module ibex_core (alert_major_o,
    alert_minor_o,
    clk_i,
    core_sleep_o,
    data_err_i,
    data_gnt_i,
    data_req_o,
    data_rvalid_i,
    data_we_o,
    debug_req_i,
    fetch_enable_i,
    instr_err_i,
    instr_gnt_i,
    instr_req_o,
    instr_rvalid_i,
    irq_external_i,
    irq_nm_i,
    irq_software_i,
    irq_timer_i,
    rst_ni,
    test_en_i,
    boot_addr_i,
    data_addr_o,
    data_be_o,
    data_rdata_i,
    data_wdata_o,
    hart_id_i,
    instr_addr_o,
    instr_rdata_i,
    irq_fast_i);
 output alert_major_o;
 output alert_minor_o;
 input clk_i;
 output core_sleep_o;
 input data_err_i;
 input data_gnt_i;
 output data_req_o;
 input data_rvalid_i;
 output data_we_o;
 input debug_req_i;
 input fetch_enable_i;
 input instr_err_i;
 input instr_gnt_i;
 output instr_req_o;
 input instr_rvalid_i;
 input irq_external_i;
 input irq_nm_i;
 input irq_software_i;
 input irq_timer_i;
 input rst_ni;
 input test_en_i;
 input [31:0] boot_addr_i;
 output [31:0] data_addr_o;
 output [3:0] data_be_o;
 input [31:0] data_rdata_i;
 output [31:0] data_wdata_o;
 input [31:0] hart_id_i;
 output [31:0] instr_addr_o;
 input [31:0] instr_rdata_i;
 input [14:0] irq_fast_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire net1083;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire net1081;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire net1077;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire net1074;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire net1067;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire net1066;
 wire net1065;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire net1064;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire net1063;
 wire net1062;
 wire net1061;
 wire net1060;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire net1059;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire net1058;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire net1057;
 wire net1056;
 wire net1055;
 wire net1054;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire net1053;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire net1052;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire net1051;
 wire _05598_;
 wire net1050;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire net1049;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire net1048;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire net1047;
 wire _05629_;
 wire _05630_;
 wire net1046;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire net1044;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire net1043;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire net1042;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire net1040;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire net1039;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire net1038;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire net1037;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire net1036;
 wire _05750_;
 wire net1035;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire net1034;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire net1033;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire net1032;
 wire net1031;
 wire _05769_;
 wire net1030;
 wire _05771_;
 wire net1029;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire net1028;
 wire _05779_;
 wire net1027;
 wire _05781_;
 wire _05782_;
 wire net1026;
 wire net1025;
 wire net1024;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire net1023;
 wire _05805_;
 wire net1022;
 wire net1021;
 wire _05808_;
 wire net1020;
 wire _05810_;
 wire net1019;
 wire net1018;
 wire _05813_;
 wire net1017;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire net1016;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire net1015;
 wire _05823_;
 wire _05824_;
 wire net1014;
 wire _05826_;
 wire _05827_;
 wire net1013;
 wire net1012;
 wire net1011;
 wire net1010;
 wire _05832_;
 wire _05833_;
 wire net1009;
 wire net1008;
 wire _05836_;
 wire _05837_;
 wire net1007;
 wire _05839_;
 wire _05840_;
 wire net1006;
 wire net1005;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire net1004;
 wire net1003;
 wire _05848_;
 wire _05849_;
 wire net1002;
 wire _05851_;
 wire _05852_;
 wire net1001;
 wire _05854_;
 wire _05855_;
 wire net1000;
 wire net999;
 wire _05858_;
 wire _05859_;
 wire net998;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire net997;
 wire net996;
 wire _05866_;
 wire _05867_;
 wire net995;
 wire _05869_;
 wire _05870_;
 wire net994;
 wire net993;
 wire _05873_;
 wire _05874_;
 wire net992;
 wire net991;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire net990;
 wire net989;
 wire _05882_;
 wire _05883_;
 wire net988;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire net987;
 wire net986;
 wire net985;
 wire net984;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire net983;
 wire net982;
 wire net981;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire net980;
 wire net979;
 wire _05903_;
 wire _05904_;
 wire net978;
 wire net977;
 wire _05907_;
 wire _05908_;
 wire net976;
 wire net975;
 wire _05911_;
 wire _05912_;
 wire net974;
 wire net973;
 wire net972;
 wire _05916_;
 wire _05917_;
 wire net971;
 wire net970;
 wire net969;
 wire _05921_;
 wire _05922_;
 wire net968;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire net967;
 wire net966;
 wire _05929_;
 wire _05930_;
 wire net965;
 wire _05932_;
 wire _05933_;
 wire net964;
 wire net963;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire net962;
 wire net961;
 wire net960;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire net959;
 wire _05946_;
 wire net957;
 wire net956;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire net955;
 wire net954;
 wire _05954_;
 wire _05955_;
 wire net953;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire net952;
 wire net951;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire net950;
 wire _05966_;
 wire _05967_;
 wire net949;
 wire net948;
 wire net947;
 wire _05971_;
 wire _05972_;
 wire net946;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire net945;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire net944;
 wire net943;
 wire net942;
 wire net941;
 wire net940;
 wire net939;
 wire net938;
 wire net937;
 wire _06103_;
 wire _06104_;
 wire net936;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire net935;
 wire _06112_;
 wire net934;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire net933;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire net932;
 wire net931;
 wire _06137_;
 wire _06138_;
 wire net930;
 wire net929;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire net928;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire net927;
 wire _06221_;
 wire net926;
 wire _06223_;
 wire net925;
 wire _06225_;
 wire net924;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire net923;
 wire net922;
 wire net921;
 wire net920;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire net919;
 wire net918;
 wire net917;
 wire _06300_;
 wire _06301_;
 wire net916;
 wire net915;
 wire _06304_;
 wire net914;
 wire net913;
 wire net912;
 wire _06308_;
 wire net911;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire net910;
 wire net909;
 wire net908;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire net907;
 wire _06332_;
 wire net906;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire net905;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire net904;
 wire _06364_;
 wire net903;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire net902;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire net901;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire net900;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire net899;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire net898;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire net897;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire net896;
 wire net895;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire net894;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire net893;
 wire _06580_;
 wire net892;
 wire net891;
 wire net890;
 wire _06584_;
 wire net889;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire net888;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire net887;
 wire net886;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire net885;
 wire net884;
 wire net883;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire net882;
 wire net881;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire net880;
 wire net879;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire net878;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire net877;
 wire net876;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire net875;
 wire net874;
 wire _06733_;
 wire _06734_;
 wire net873;
 wire net872;
 wire _06737_;
 wire net871;
 wire net870;
 wire _06740_;
 wire _06741_;
 wire net869;
 wire net868;
 wire _06744_;
 wire net867;
 wire net866;
 wire net865;
 wire net864;
 wire net863;
 wire _06750_;
 wire net862;
 wire _06752_;
 wire net861;
 wire net860;
 wire _06755_;
 wire net859;
 wire net858;
 wire _06758_;
 wire net857;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire net856;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire net855;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire net854;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire net853;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire net852;
 wire _06833_;
 wire _06834_;
 wire net851;
 wire net850;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire net849;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire net847;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire net846;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire net845;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire net844;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire net843;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire net842;
 wire _06987_;
 wire net841;
 wire net840;
 wire _06990_;
 wire net839;
 wire _06992_;
 wire net838;
 wire _06994_;
 wire net837;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire net836;
 wire _07000_;
 wire net835;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire net834;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire net833;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire net832;
 wire _07016_;
 wire net831;
 wire net830;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire net829;
 wire _07026_;
 wire net828;
 wire _07028_;
 wire net827;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire net826;
 wire _07041_;
 wire net825;
 wire net824;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire net823;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire net822;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire net821;
 wire net820;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire net819;
 wire _07064_;
 wire _07065_;
 wire net818;
 wire _07067_;
 wire _07068_;
 wire net817;
 wire net816;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire net815;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire net814;
 wire net813;
 wire _07080_;
 wire net812;
 wire _07082_;
 wire _07083_;
 wire net811;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire net810;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire net809;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire net808;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire net807;
 wire _07120_;
 wire _07121_;
 wire net806;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire net805;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire net804;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire net803;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire net802;
 wire net801;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire net800;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire net799;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire net798;
 wire net797;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire net796;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire net795;
 wire _07227_;
 wire net794;
 wire _07229_;
 wire net793;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire net792;
 wire net791;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire net790;
 wire _07250_;
 wire net789;
 wire net788;
 wire _07253_;
 wire net787;
 wire net786;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire net785;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire net784;
 wire _07264_;
 wire _07265_;
 wire net783;
 wire _07267_;
 wire net782;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire net781;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire net780;
 wire _07283_;
 wire net779;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire net778;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire net777;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire net776;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire net775;
 wire net774;
 wire net773;
 wire net772;
 wire net771;
 wire net770;
 wire net769;
 wire _07350_;
 wire net768;
 wire _07352_;
 wire _07353_;
 wire net767;
 wire _07355_;
 wire _07356_;
 wire net766;
 wire net765;
 wire _07359_;
 wire _07360_;
 wire net764;
 wire net763;
 wire _07363_;
 wire _07364_;
 wire net762;
 wire _07366_;
 wire _07367_;
 wire net761;
 wire _07369_;
 wire net760;
 wire _07371_;
 wire _07372_;
 wire net759;
 wire net758;
 wire net757;
 wire _07376_;
 wire net756;
 wire net755;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire net754;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire net753;
 wire _07421_;
 wire net752;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire net751;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire net750;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire net749;
 wire net748;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire net747;
 wire net746;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire net745;
 wire net744;
 wire net743;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire net742;
 wire net741;
 wire net740;
 wire net739;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire net738;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire net737;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire net736;
 wire _07524_;
 wire net735;
 wire _07526_;
 wire net734;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire net733;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire net732;
 wire net731;
 wire net730;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire net729;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire net728;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire net727;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire net726;
 wire _07590_;
 wire _07591_;
 wire net725;
 wire net724;
 wire net723;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire net722;
 wire net721;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire net720;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire net719;
 wire _07634_;
 wire net718;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire net717;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire net716;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire net715;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire net714;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire net713;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire net712;
 wire net711;
 wire net710;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire net709;
 wire _07762_;
 wire _07763_;
 wire net708;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire net707;
 wire net706;
 wire net705;
 wire _07784_;
 wire _07785_;
 wire net704;
 wire net703;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire net702;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire net701;
 wire net700;
 wire net699;
 wire net698;
 wire _07803_;
 wire _07804_;
 wire net697;
 wire net696;
 wire _07807_;
 wire net695;
 wire _07809_;
 wire _07810_;
 wire net694;
 wire _07812_;
 wire _07813_;
 wire net693;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire net692;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire net691;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire net690;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire net689;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire net688;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire net687;
 wire net686;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire net685;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire net684;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire net683;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire net682;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire net681;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire net680;
 wire net679;
 wire net678;
 wire _08664_;
 wire _08665_;
 wire net677;
 wire net676;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire net675;
 wire net674;
 wire _08675_;
 wire net673;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire net672;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire net671;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire net670;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire net669;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire net668;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire net667;
 wire net666;
 wire _08768_;
 wire net665;
 wire net664;
 wire _08771_;
 wire _08772_;
 wire net663;
 wire _08774_;
 wire net662;
 wire net661;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire net660;
 wire _08788_;
 wire _08789_;
 wire net659;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire net658;
 wire _08798_;
 wire net657;
 wire _08800_;
 wire net656;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire net655;
 wire net654;
 wire net653;
 wire net652;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire net651;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire net650;
 wire net649;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire net648;
 wire net647;
 wire _08845_;
 wire _08846_;
 wire net646;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire net645;
 wire net644;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire net643;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire net642;
 wire net641;
 wire _09142_;
 wire net640;
 wire net639;
 wire _09145_;
 wire _09146_;
 wire net638;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire net633;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire net632;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire net631;
 wire net630;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire net629;
 wire _09229_;
 wire net628;
 wire _09231_;
 wire net627;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire net626;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire net625;
 wire net624;
 wire net623;
 wire _09261_;
 wire _09262_;
 wire net622;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire net621;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire net620;
 wire _09276_;
 wire _09277_;
 wire net619;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire net618;
 wire net617;
 wire net616;
 wire net615;
 wire _09324_;
 wire net614;
 wire net613;
 wire _09327_;
 wire net612;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire net611;
 wire net610;
 wire _09335_;
 wire _09336_;
 wire net609;
 wire net608;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire net607;
 wire net606;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire net605;
 wire _09398_;
 wire net604;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire net603;
 wire _09445_;
 wire _09446_;
 wire net602;
 wire net601;
 wire _09449_;
 wire _09450_;
 wire net600;
 wire _09452_;
 wire net599;
 wire _09454_;
 wire net598;
 wire _09456_;
 wire net597;
 wire _09458_;
 wire net596;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire net595;
 wire net594;
 wire net593;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire net592;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire net591;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire net590;
 wire _09493_;
 wire net589;
 wire net588;
 wire net587;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire net586;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire net585;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire net584;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire net583;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire net582;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire net581;
 wire net580;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire net579;
 wire _09568_;
 wire _09569_;
 wire net578;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire net577;
 wire net576;
 wire net575;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire net574;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire net573;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire net572;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire net571;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire net570;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire net569;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire net568;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire net567;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire net566;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire net565;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire net564;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire net563;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire net562;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire net561;
 wire net560;
 wire _09760_;
 wire net559;
 wire _09762_;
 wire net558;
 wire net557;
 wire _09765_;
 wire net556;
 wire _09767_;
 wire net555;
 wire net554;
 wire _09770_;
 wire net553;
 wire _09772_;
 wire net552;
 wire _09774_;
 wire net551;
 wire _09776_;
 wire net550;
 wire _09778_;
 wire net549;
 wire _09780_;
 wire net548;
 wire _09782_;
 wire net547;
 wire _09784_;
 wire net546;
 wire net545;
 wire _09787_;
 wire net544;
 wire _09789_;
 wire net543;
 wire _09791_;
 wire net542;
 wire _09793_;
 wire net541;
 wire _09795_;
 wire net540;
 wire _09797_;
 wire net539;
 wire _09799_;
 wire net538;
 wire _09801_;
 wire net537;
 wire _09803_;
 wire net536;
 wire _09805_;
 wire net535;
 wire net534;
 wire _09808_;
 wire net533;
 wire _09810_;
 wire net532;
 wire _09812_;
 wire net531;
 wire _09814_;
 wire net530;
 wire _09816_;
 wire net529;
 wire _09818_;
 wire net528;
 wire _09820_;
 wire net527;
 wire _09822_;
 wire net526;
 wire _09824_;
 wire net525;
 wire _09826_;
 wire net524;
 wire _09828_;
 wire _09829_;
 wire net523;
 wire _09831_;
 wire net522;
 wire net521;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire net520;
 wire _09842_;
 wire _09843_;
 wire net519;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire net518;
 wire _09854_;
 wire _09855_;
 wire net517;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire net516;
 wire net515;
 wire net514;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire net513;
 wire _09885_;
 wire _09886_;
 wire net512;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire net511;
 wire _09897_;
 wire _09898_;
 wire net510;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire net509;
 wire net508;
 wire _09918_;
 wire net507;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire net506;
 wire net505;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire net504;
 wire net503;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire net502;
 wire _09957_;
 wire _09958_;
 wire net501;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire net500;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire net499;
 wire _09972_;
 wire net498;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire net497;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire net496;
 wire _09995_;
 wire _09996_;
 wire net495;
 wire net494;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire net493;
 wire _10007_;
 wire _10008_;
 wire net492;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire net491;
 wire _10019_;
 wire _10020_;
 wire net490;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire net489;
 wire net488;
 wire net487;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire net486;
 wire _10049_;
 wire _10050_;
 wire net485;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire net484;
 wire _10061_;
 wire _10062_;
 wire net483;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire net482;
 wire _10080_;
 wire net481;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire net480;
 wire net479;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire net478;
 wire net477;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire net476;
 wire _10119_;
 wire _10120_;
 wire net475;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire net474;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire net473;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire net472;
 wire _10139_;
 wire _10140_;
 wire net471;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire net470;
 wire _10147_;
 wire net469;
 wire _10149_;
 wire _10150_;
 wire net468;
 wire _10152_;
 wire _10153_;
 wire net466;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire net465;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire net464;
 wire net463;
 wire _10165_;
 wire net462;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire net461;
 wire _10172_;
 wire _10173_;
 wire net460;
 wire _10175_;
 wire net459;
 wire _10177_;
 wire net458;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire net457;
 wire _10183_;
 wire net456;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire net455;
 wire _10189_;
 wire net454;
 wire _10191_;
 wire net453;
 wire _10193_;
 wire net452;
 wire _10195_;
 wire net451;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire net450;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire net449;
 wire _10207_;
 wire net448;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire net447;
 wire net446;
 wire net445;
 wire _10218_;
 wire _10219_;
 wire net444;
 wire _10221_;
 wire net443;
 wire _10223_;
 wire net442;
 wire _10225_;
 wire _10226_;
 wire net441;
 wire _10228_;
 wire net440;
 wire net439;
 wire _10231_;
 wire _10232_;
 wire net438;
 wire net437;
 wire _10235_;
 wire net436;
 wire _10237_;
 wire net435;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire net434;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire net433;
 wire net432;
 wire _10248_;
 wire _10249_;
 wire net431;
 wire net430;
 wire _10252_;
 wire _10253_;
 wire net429;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire net428;
 wire _10260_;
 wire _10261_;
 wire net427;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire net426;
 wire _10271_;
 wire net425;
 wire net424;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire net423;
 wire _10282_;
 wire _10283_;
 wire net422;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire net421;
 wire _10294_;
 wire _10295_;
 wire net420;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire net419;
 wire net418;
 wire net417;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire net416;
 wire _10322_;
 wire _10323_;
 wire net415;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire net414;
 wire _10334_;
 wire _10335_;
 wire net413;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire net412;
 wire _10352_;
 wire _10353_;
 wire net411;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire net410;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire net409;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire net408;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire net407;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire net406;
 wire _10392_;
 wire net405;
 wire _10394_;
 wire _10395_;
 wire net404;
 wire _10397_;
 wire net403;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire net402;
 wire net401;
 wire _10410_;
 wire net400;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net399;
 wire _10434_;
 wire net398;
 wire _10436_;
 wire net397;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire net396;
 wire net395;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire net394;
 wire net393;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire net392;
 wire net391;
 wire net390;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire net389;
 wire _10486_;
 wire _10487_;
 wire net388;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire net387;
 wire _10498_;
 wire _10499_;
 wire net386;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire net385;
 wire _10516_;
 wire net384;
 wire _10518_;
 wire _10519_;
 wire net383;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire net382;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire net381;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire net380;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire net379;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire net378;
 wire _10559_;
 wire net377;
 wire net376;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire net375;
 wire _10573_;
 wire _10574_;
 wire net374;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire net373;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire net372;
 wire _10598_;
 wire net371;
 wire net370;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire net369;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire net368;
 wire _10610_;
 wire net367;
 wire net366;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire net365;
 wire _10618_;
 wire _10619_;
 wire net364;
 wire _10621_;
 wire net363;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire net362;
 wire net361;
 wire _10628_;
 wire net360;
 wire _10630_;
 wire _10631_;
 wire net359;
 wire _10633_;
 wire _10634_;
 wire net358;
 wire _10636_;
 wire _10637_;
 wire net357;
 wire _10639_;
 wire _10640_;
 wire net356;
 wire _10642_;
 wire _10643_;
 wire net355;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire net354;
 wire _10649_;
 wire _10650_;
 wire net353;
 wire _10652_;
 wire net352;
 wire _10654_;
 wire net351;
 wire _10656_;
 wire net350;
 wire _10658_;
 wire _10659_;
 wire net349;
 wire _10661_;
 wire net348;
 wire net347;
 wire _10664_;
 wire _10665_;
 wire net346;
 wire _10667_;
 wire net345;
 wire _10669_;
 wire net344;
 wire net343;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire net342;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire net341;
 wire _10680_;
 wire net340;
 wire net339;
 wire _10683_;
 wire net338;
 wire _10685_;
 wire _10686_;
 wire net337;
 wire _10688_;
 wire net336;
 wire _10690_;
 wire net335;
 wire _10692_;
 wire _10693_;
 wire net334;
 wire _10695_;
 wire _10696_;
 wire net333;
 wire _10698_;
 wire _10699_;
 wire net332;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire net331;
 wire _10706_;
 wire _10707_;
 wire net330;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire net329;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire net328;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire net327;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire net326;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire net325;
 wire _10746_;
 wire net324;
 wire _10748_;
 wire net323;
 wire net322;
 wire _10751_;
 wire net321;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire net320;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire net319;
 wire net318;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire net317;
 wire _10796_;
 wire net316;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire net315;
 wire _10808_;
 wire net314;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire net313;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire net312;
 wire net311;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire net310;
 wire net309;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire net308;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire net307;
 wire _10865_;
 wire _10866_;
 wire net306;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire net305;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire net304;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire net303;
 wire _10889_;
 wire _10890_;
 wire net302;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire net301;
 wire net300;
 wire net299;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire net298;
 wire _10916_;
 wire _10917_;
 wire net297;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire net296;
 wire _10928_;
 wire _10929_;
 wire net295;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire net294;
 wire net293;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire net292;
 wire _10958_;
 wire net291;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire net290;
 wire _10970_;
 wire net289;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire net288;
 wire net287;
 wire net286;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire net285;
 wire _10997_;
 wire _10998_;
 wire net284;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire net283;
 wire _11009_;
 wire _11010_;
 wire net282;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire net281;
 wire _11027_;
 wire _11028_;
 wire net280;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire net279;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire net278;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire net277;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire net276;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire net275;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire net274;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire net273;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire net272;
 wire net271;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire net270;
 wire _11122_;
 wire _11123_;
 wire net269;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire net268;
 wire _11143_;
 wire _11144_;
 wire net267;
 wire net266;
 wire _11147_;
 wire _11148_;
 wire net265;
 wire _11150_;
 wire net264;
 wire _11152_;
 wire net263;
 wire net262;
 wire _11155_;
 wire _11156_;
 wire net261;
 wire net260;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire net259;
 wire net258;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire net257;
 wire _11169_;
 wire net256;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire net255;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire net254;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire net253;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire net252;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire net251;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire net250;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire net249;
 wire _11292_;
 wire net248;
 wire net247;
 wire _11295_;
 wire net246;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire net245;
 wire net244;
 wire _11302_;
 wire net243;
 wire net242;
 wire _11305_;
 wire _11306_;
 wire net241;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire net240;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire net239;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire net238;
 wire net237;
 wire _11411_;
 wire _11412_;
 wire net236;
 wire _11414_;
 wire net235;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire net234;
 wire net233;
 wire net232;
 wire _11435_;
 wire net231;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire net230;
 wire net229;
 wire _11443_;
 wire _11444_;
 wire net228;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire net227;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire net226;
 wire _11477_;
 wire net225;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire net224;
 wire net223;
 wire net222;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire net221;
 wire net220;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire net219;
 wire net218;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire net217;
 wire net216;
 wire _11550_;
 wire net215;
 wire _11552_;
 wire _11553_;
 wire net214;
 wire _11555_;
 wire _11556_;
 wire net213;
 wire _11558_;
 wire net212;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire net211;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire net210;
 wire net209;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire net208;
 wire _11647_;
 wire net207;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire net206;
 wire _11659_;
 wire net205;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire net204;
 wire _11675_;
 wire net203;
 wire net202;
 wire _11678_;
 wire net201;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire net200;
 wire net199;
 wire net198;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire net197;
 wire net196;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire net195;
 wire _11707_;
 wire net194;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire net193;
 wire _11719_;
 wire net192;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire net191;
 wire _11736_;
 wire net190;
 wire _11738_;
 wire net189;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire net188;
 wire net187;
 wire net186;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire net185;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire net184;
 wire _11800_;
 wire net183;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire net182;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire net181;
 wire net180;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire net179;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire net178;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire net177;
 wire net176;
 wire net175;
 wire net174;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire net173;
 wire _11915_;
 wire _11916_;
 wire net172;
 wire _11918_;
 wire _11919_;
 wire net171;
 wire net170;
 wire net169;
 wire net168;
 wire net167;
 wire _11925_;
 wire net166;
 wire net165;
 wire net164;
 wire net163;
 wire _11930_;
 wire _11931_;
 wire net162;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire net161;
 wire _11937_;
 wire net160;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire net159;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire net158;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire net157;
 wire net156;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire net155;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire net154;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire net153;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire net152;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire net151;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire net150;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire net149;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire net148;
 wire net147;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire net146;
 wire _12176_;
 wire _12177_;
 wire net145;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire net144;
 wire _12188_;
 wire _12189_;
 wire net143;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire net142;
 wire net141;
 wire _12209_;
 wire _12210_;
 wire net140;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire net139;
 wire _12234_;
 wire net138;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire net137;
 wire _12242_;
 wire _12243_;
 wire net136;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire net135;
 wire net134;
 wire net133;
 wire net132;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire net131;
 wire net130;
 wire net129;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire net128;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire net127;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire net126;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire net125;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire net124;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire net123;
 wire net122;
 wire _12442_;
 wire net121;
 wire net120;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire net119;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire net118;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire net117;
 wire _12480_;
 wire _12481_;
 wire net116;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire net115;
 wire _12501_;
 wire _12502_;
 wire net114;
 wire _12504_;
 wire net113;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire net112;
 wire _12524_;
 wire _12525_;
 wire net111;
 wire _12527_;
 wire net110;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire net109;
 wire net108;
 wire _12559_;
 wire net107;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire net106;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire net105;
 wire _12597_;
 wire net104;
 wire _12599_;
 wire net103;
 wire _12601_;
 wire _12602_;
 wire net102;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire net101;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire net100;
 wire _12632_;
 wire net99;
 wire _12634_;
 wire net98;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire net97;
 wire net96;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire net95;
 wire net94;
 wire net93;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire net92;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire net91;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire net90;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire net89;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire net88;
 wire net87;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire net86;
 wire net85;
 wire net84;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire net83;
 wire net82;
 wire _12736_;
 wire net81;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire net80;
 wire _12744_;
 wire net79;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire net78;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire net77;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire net76;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire net75;
 wire _12773_;
 wire net74;
 wire net73;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire net72;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire net71;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire net70;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire net69;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire net68;
 wire net67;
 wire net66;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire net65;
 wire net64;
 wire net63;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire net62;
 wire net61;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire net60;
 wire net59;
 wire _12843_;
 wire net58;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire net57;
 wire net56;
 wire net55;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire net54;
 wire net53;
 wire net52;
 wire _12869_;
 wire net51;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire net50;
 wire net49;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire net48;
 wire net47;
 wire _12918_;
 wire _12919_;
 wire net46;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire net45;
 wire _12932_;
 wire net44;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire net43;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire net42;
 wire _12943_;
 wire net41;
 wire _12945_;
 wire net40;
 wire _12947_;
 wire _12948_;
 wire net39;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire net38;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire net37;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire net36;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire net35;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire net34;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire net33;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire net32;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire net31;
 wire _13141_;
 wire _13142_;
 wire net30;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire net1654;
 wire net1653;
 wire net1652;
 wire net1651;
 wire net1650;
 wire _13340_;
 wire net1649;
 wire _13342_;
 wire net1648;
 wire net1647;
 wire _13345_;
 wire net1646;
 wire net1645;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire net1644;
 wire net1643;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire net1642;
 wire _13359_;
 wire net1641;
 wire net1640;
 wire net1639;
 wire net1638;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire net1637;
 wire net1636;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire net1635;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire net1634;
 wire net1633;
 wire _13380_;
 wire net1632;
 wire _13382_;
 wire _13383_;
 wire net1631;
 wire _13385_;
 wire net1630;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire net1629;
 wire net1628;
 wire _13394_;
 wire _13395_;
 wire net1627;
 wire net1626;
 wire net1625;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire net1624;
 wire net1623;
 wire _13405_;
 wire _13406_;
 wire net1622;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire net1621;
 wire _13414_;
 wire _13415_;
 wire net1620;
 wire net1619;
 wire _13418_;
 wire _13419_;
 wire net1618;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire net1617;
 wire net1616;
 wire _13426_;
 wire net1615;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire net1614;
 wire net1613;
 wire _13433_;
 wire _13434_;
 wire net1612;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire net1611;
 wire _13441_;
 wire _13442_;
 wire net1610;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire net1609;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire net1608;
 wire net1607;
 wire net1606;
 wire net1605;
 wire net1604;
 wire _13456_;
 wire _13457_;
 wire net1603;
 wire _13459_;
 wire _13460_;
 wire net1602;
 wire net1601;
 wire _13463_;
 wire net1600;
 wire _13465_;
 wire net1599;
 wire _13467_;
 wire net1598;
 wire net1597;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire net1596;
 wire _13476_;
 wire net1595;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire net1594;
 wire _13492_;
 wire net1593;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire net1592;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire net1591;
 wire net1590;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire net1589;
 wire _13525_;
 wire net1586;
 wire net1585;
 wire _13528_;
 wire net1584;
 wire net1583;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire net1582;
 wire net1581;
 wire _13537_;
 wire _13538_;
 wire net1580;
 wire net1579;
 wire net1578;
 wire net1577;
 wire net1576;
 wire net1575;
 wire net1574;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire net1573;
 wire net1572;
 wire _13558_;
 wire _13559_;
 wire net1571;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire net1570;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire net1569;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire net1568;
 wire _13620_;
 wire net1567;
 wire net1566;
 wire _13623_;
 wire net1565;
 wire net1564;
 wire _13626_;
 wire net1563;
 wire net1562;
 wire net1561;
 wire _13630_;
 wire net1560;
 wire net1559;
 wire net1558;
 wire net1557;
 wire net1556;
 wire _13636_;
 wire net1555;
 wire _13638_;
 wire net1554;
 wire net1553;
 wire net1552;
 wire net1551;
 wire net1550;
 wire net1549;
 wire net1548;
 wire net1547;
 wire _13647_;
 wire net1546;
 wire _13649_;
 wire net1545;
 wire net1544;
 wire net1543;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire net1542;
 wire net1541;
 wire net1540;
 wire net1539;
 wire _13660_;
 wire _13661_;
 wire net1538;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire net1537;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire net1536;
 wire net1535;
 wire net1534;
 wire _13675_;
 wire net1533;
 wire net1532;
 wire net1531;
 wire _13679_;
 wire net1530;
 wire net1529;
 wire net1528;
 wire net1527;
 wire net1526;
 wire _13685_;
 wire net1525;
 wire _13687_;
 wire _13688_;
 wire net1524;
 wire net1523;
 wire net1522;
 wire net1521;
 wire net1520;
 wire net1519;
 wire net1518;
 wire net1517;
 wire net1516;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire net1515;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire net1514;
 wire net1513;
 wire net1512;
 wire net1511;
 wire net1510;
 wire _13710_;
 wire _13711_;
 wire net1509;
 wire net1508;
 wire net1507;
 wire net1506;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire net1505;
 wire net1504;
 wire net1503;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire net1502;
 wire net1501;
 wire net1500;
 wire net1499;
 wire net1498;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire net1497;
 wire net1496;
 wire net1495;
 wire _13740_;
 wire net1494;
 wire net1493;
 wire net1492;
 wire _13744_;
 wire _13745_;
 wire net1491;
 wire net1490;
 wire net1489;
 wire net1488;
 wire net1487;
 wire _13751_;
 wire net1486;
 wire net1485;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire net1484;
 wire net1483;
 wire net1482;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire net1481;
 wire net1480;
 wire net1479;
 wire _13771_;
 wire _13772_;
 wire net1478;
 wire net1477;
 wire _13775_;
 wire net1476;
 wire net1475;
 wire _13778_;
 wire net1474;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire net1473;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire net1472;
 wire net1471;
 wire _13797_;
 wire net1470;
 wire net1469;
 wire net1468;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire net1467;
 wire net1466;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire net1465;
 wire _13817_;
 wire net1464;
 wire net1463;
 wire net1462;
 wire net1461;
 wire _13822_;
 wire _13823_;
 wire net1460;
 wire _13825_;
 wire net1459;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire net1458;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire net1457;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire net1456;
 wire _13853_;
 wire net1455;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire net1454;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire net1453;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire net1452;
 wire net1451;
 wire net1449;
 wire net1448;
 wire net1447;
 wire net1445;
 wire net1444;
 wire net1443;
 wire _13903_;
 wire net1442;
 wire net1441;
 wire _13906_;
 wire net1440;
 wire net1439;
 wire _13909_;
 wire _13910_;
 wire net1438;
 wire net1437;
 wire net1436;
 wire _13914_;
 wire _13915_;
 wire net1435;
 wire net1434;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire net1433;
 wire net1432;
 wire net1431;
 wire net1430;
 wire net1429;
 wire _13927_;
 wire net1428;
 wire _13929_;
 wire net1427;
 wire _13931_;
 wire net1426;
 wire net1425;
 wire _13934_;
 wire net1424;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire net1423;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire net1422;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire net1421;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire net1420;
 wire net1419;
 wire net1418;
 wire net1417;
 wire _13964_;
 wire _13965_;
 wire net1416;
 wire net1415;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire net1414;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire net1413;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire net1412;
 wire net1411;
 wire net1410;
 wire _13985_;
 wire _13986_;
 wire net1409;
 wire _13988_;
 wire _13989_;
 wire net1408;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire net1407;
 wire net1406;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire net1404;
 wire _14001_;
 wire _14002_;
 wire net1403;
 wire net1401;
 wire _14005_;
 wire net1400;
 wire net1399;
 wire _14008_;
 wire net1398;
 wire net1397;
 wire _14011_;
 wire _14012_;
 wire net1396;
 wire _14014_;
 wire _14015_;
 wire net1395;
 wire net1394;
 wire net1393;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire net1392;
 wire _14029_;
 wire _14030_;
 wire net1391;
 wire net1390;
 wire _14033_;
 wire net1389;
 wire net1388;
 wire _14036_;
 wire net1387;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire net1386;
 wire net1385;
 wire _14049_;
 wire _14050_;
 wire net1384;
 wire _14052_;
 wire net1383;
 wire net1382;
 wire _14055_;
 wire net1381;
 wire _14057_;
 wire net1380;
 wire _14059_;
 wire _14060_;
 wire net1379;
 wire _14062_;
 wire _14063_;
 wire net1378;
 wire net1377;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire net1376;
 wire net1375;
 wire _14072_;
 wire net1374;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire net1373;
 wire _14078_;
 wire _14079_;
 wire net1372;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire net1371;
 wire _14085_;
 wire _14086_;
 wire net1370;
 wire net1369;
 wire net1368;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire net1367;
 wire net1366;
 wire net1365;
 wire _14103_;
 wire _14104_;
 wire net1364;
 wire net1363;
 wire _14107_;
 wire net1362;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire net1361;
 wire _14114_;
 wire net1360;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire net1359;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire net1358;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire net1357;
 wire _14158_;
 wire _14159_;
 wire net1356;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire net1355;
 wire _14171_;
 wire net1354;
 wire _14173_;
 wire _14174_;
 wire net1353;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire net1351;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire net1350;
 wire net1349;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire net1348;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire net1345;
 wire net1344;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire net1343;
 wire net1341;
 wire net1339;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire net1338;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire net1337;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire net1336;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire net1335;
 wire net1333;
 wire _14362_;
 wire _14363_;
 wire net1332;
 wire net1331;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire net1330;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire net1329;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire net1328;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire net1326;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire net1325;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire net1324;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire net1323;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire net1322;
 wire _14546_;
 wire net1321;
 wire net1320;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire net1319;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire net1317;
 wire net1316;
 wire _14614_;
 wire _14615_;
 wire net1315;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire net1311;
 wire _14716_;
 wire net1310;
 wire _14718_;
 wire _14719_;
 wire net1309;
 wire net1308;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire net1307;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire net1306;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire net1305;
 wire net1304;
 wire _14745_;
 wire net1303;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire net1302;
 wire net1301;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire net1300;
 wire net1299;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire net1298;
 wire net1297;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire net1296;
 wire _14782_;
 wire _14783_;
 wire net1295;
 wire net1294;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire net1293;
 wire net1292;
 wire _14791_;
 wire net1291;
 wire _14793_;
 wire _14794_;
 wire net1290;
 wire _14796_;
 wire _14797_;
 wire net1289;
 wire _14799_;
 wire net1288;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire net1287;
 wire _14845_;
 wire net1286;
 wire net1285;
 wire net1284;
 wire net1283;
 wire net1282;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire net1281;
 wire net1280;
 wire _14857_;
 wire net1279;
 wire net1278;
 wire _14860_;
 wire net1277;
 wire net1276;
 wire net1275;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire net1274;
 wire net1273;
 wire _14870_;
 wire net1272;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire net1271;
 wire _14882_;
 wire _14883_;
 wire net1270;
 wire _14885_;
 wire _14886_;
 wire net1269;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire net1268;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire net1267;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire net1266;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire net1265;
 wire _14945_;
 wire _14946_;
 wire net1264;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire net1263;
 wire _14952_;
 wire net1262;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire net1261;
 wire _14982_;
 wire _14983_;
 wire net1260;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire net1259;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire net1258;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire net1257;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire net1256;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire net1255;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire net1254;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire _15051_;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire _15056_;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire net1253;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire net1252;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire net1251;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire net1250;
 wire _15105_;
 wire _15106_;
 wire net1249;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire _15123_;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire _15128_;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire net1247;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire net1245;
 wire _15174_;
 wire _15175_;
 wire net1244;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire net1243;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire _15200_;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire _15227_;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire net1241;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire _15332_;
 wire _15333_;
 wire _15334_;
 wire _15335_;
 wire _15336_;
 wire _15337_;
 wire net1238;
 wire _15339_;
 wire _15340_;
 wire _15341_;
 wire _15342_;
 wire _15343_;
 wire _15344_;
 wire _15345_;
 wire _15346_;
 wire _15347_;
 wire _15348_;
 wire _15349_;
 wire _15350_;
 wire _15351_;
 wire _15352_;
 wire _15353_;
 wire _15354_;
 wire _15355_;
 wire _15356_;
 wire _15357_;
 wire _15358_;
 wire _15359_;
 wire _15360_;
 wire _15361_;
 wire _15362_;
 wire _15363_;
 wire _15364_;
 wire _15365_;
 wire _15366_;
 wire _15367_;
 wire _15368_;
 wire _15369_;
 wire _15370_;
 wire _15371_;
 wire _15372_;
 wire _15373_;
 wire _15374_;
 wire _15375_;
 wire _15376_;
 wire _15377_;
 wire _15378_;
 wire _15379_;
 wire _15380_;
 wire _15381_;
 wire _15382_;
 wire _15383_;
 wire _15384_;
 wire _15385_;
 wire _15386_;
 wire _15387_;
 wire _15388_;
 wire _15389_;
 wire _15390_;
 wire _15391_;
 wire _15392_;
 wire _15393_;
 wire _15394_;
 wire _15395_;
 wire _15396_;
 wire net1237;
 wire _15398_;
 wire _15399_;
 wire _15400_;
 wire _15401_;
 wire _15402_;
 wire net1235;
 wire _15404_;
 wire _15405_;
 wire _15406_;
 wire _15407_;
 wire _15408_;
 wire _15409_;
 wire _15410_;
 wire net1234;
 wire net1233;
 wire net1232;
 wire net1231;
 wire net1230;
 wire net1229;
 wire net1228;
 wire net1227;
 wire net1226;
 wire net1225;
 wire _15421_;
 wire _15422_;
 wire net1224;
 wire net1223;
 wire net1222;
 wire _15426_;
 wire net1221;
 wire net1220;
 wire net1219;
 wire net1218;
 wire _15431_;
 wire net1217;
 wire net1216;
 wire _15434_;
 wire net1215;
 wire _15436_;
 wire net1214;
 wire _15438_;
 wire _15439_;
 wire _15440_;
 wire net1213;
 wire net1212;
 wire net1211;
 wire _15444_;
 wire _15445_;
 wire net1210;
 wire _15447_;
 wire net1209;
 wire _15449_;
 wire _15450_;
 wire _15451_;
 wire net1208;
 wire _15453_;
 wire _15454_;
 wire _15455_;
 wire _15456_;
 wire _15457_;
 wire _15458_;
 wire net1207;
 wire net1206;
 wire _15461_;
 wire _15462_;
 wire _15463_;
 wire _15464_;
 wire _15465_;
 wire _15466_;
 wire _15467_;
 wire net1205;
 wire net1204;
 wire _15470_;
 wire _15471_;
 wire _15472_;
 wire _15473_;
 wire net1203;
 wire _15475_;
 wire _15476_;
 wire _15477_;
 wire _15478_;
 wire _15479_;
 wire _15480_;
 wire _15481_;
 wire _15482_;
 wire _15483_;
 wire _15484_;
 wire _15485_;
 wire _15486_;
 wire _15487_;
 wire _15488_;
 wire _15489_;
 wire _15490_;
 wire net1202;
 wire _15492_;
 wire net1201;
 wire _15494_;
 wire net1200;
 wire net1199;
 wire net1198;
 wire net1197;
 wire net1196;
 wire net1195;
 wire net1194;
 wire net1193;
 wire net1192;
 wire net1191;
 wire _15505_;
 wire net1190;
 wire _15507_;
 wire _15508_;
 wire net1189;
 wire _15510_;
 wire net1188;
 wire _15512_;
 wire net1187;
 wire _15514_;
 wire _15515_;
 wire net1186;
 wire net1185;
 wire _15518_;
 wire net1184;
 wire _15520_;
 wire net1183;
 wire _15522_;
 wire _15523_;
 wire _15524_;
 wire net1182;
 wire _15526_;
 wire _15527_;
 wire _15528_;
 wire net1181;
 wire net1180;
 wire net1179;
 wire net1178;
 wire _15533_;
 wire _15534_;
 wire _15535_;
 wire net1177;
 wire _15537_;
 wire _15538_;
 wire net1176;
 wire _15540_;
 wire _15541_;
 wire _15542_;
 wire net1175;
 wire _15544_;
 wire _15545_;
 wire _15546_;
 wire _15547_;
 wire net1174;
 wire net1173;
 wire net1172;
 wire _15551_;
 wire net1171;
 wire _15553_;
 wire net1170;
 wire _15555_;
 wire net1169;
 wire _15557_;
 wire net1168;
 wire _15559_;
 wire net1167;
 wire _15561_;
 wire _15562_;
 wire net1166;
 wire _15564_;
 wire _15565_;
 wire _15566_;
 wire _15567_;
 wire net1165;
 wire _15569_;
 wire _15570_;
 wire _15571_;
 wire _15572_;
 wire _15573_;
 wire _15574_;
 wire _15575_;
 wire net1164;
 wire _15577_;
 wire _15578_;
 wire _15579_;
 wire _15580_;
 wire _15581_;
 wire _15582_;
 wire _15583_;
 wire _15584_;
 wire _15585_;
 wire _15586_;
 wire _15587_;
 wire _15588_;
 wire _15589_;
 wire _15590_;
 wire _15591_;
 wire _15592_;
 wire _15593_;
 wire _15594_;
 wire _15595_;
 wire _15596_;
 wire _15597_;
 wire _15598_;
 wire _15599_;
 wire _15600_;
 wire _15601_;
 wire _15602_;
 wire _15603_;
 wire _15604_;
 wire _15605_;
 wire net1163;
 wire _15607_;
 wire _15608_;
 wire _15609_;
 wire _15610_;
 wire _15611_;
 wire _15612_;
 wire _15613_;
 wire _15614_;
 wire _15615_;
 wire _15616_;
 wire _15617_;
 wire _15618_;
 wire _15619_;
 wire _15620_;
 wire _15621_;
 wire net1162;
 wire net1161;
 wire _15624_;
 wire _15625_;
 wire _15626_;
 wire _15627_;
 wire _15628_;
 wire _15629_;
 wire _15630_;
 wire net1160;
 wire _15632_;
 wire _15633_;
 wire _15634_;
 wire _15635_;
 wire _15636_;
 wire _15637_;
 wire _15638_;
 wire _15639_;
 wire _15640_;
 wire _15641_;
 wire _15642_;
 wire _15643_;
 wire net1159;
 wire _15645_;
 wire _15646_;
 wire _15647_;
 wire _15648_;
 wire _15649_;
 wire _15650_;
 wire _15651_;
 wire _15652_;
 wire _15653_;
 wire _15654_;
 wire _15655_;
 wire _15656_;
 wire net1158;
 wire net1157;
 wire _15659_;
 wire _15660_;
 wire _15661_;
 wire net1156;
 wire _15663_;
 wire _15664_;
 wire _15665_;
 wire _15666_;
 wire net1155;
 wire _15668_;
 wire _15669_;
 wire _15670_;
 wire _15671_;
 wire net1154;
 wire net1153;
 wire _15674_;
 wire net1152;
 wire _15676_;
 wire _15677_;
 wire net1151;
 wire _15679_;
 wire _15680_;
 wire _15681_;
 wire _15682_;
 wire _15683_;
 wire _15684_;
 wire _15685_;
 wire _15686_;
 wire _15687_;
 wire _15688_;
 wire _15689_;
 wire _15690_;
 wire _15691_;
 wire _15692_;
 wire _15693_;
 wire _15694_;
 wire _15695_;
 wire _15696_;
 wire _15697_;
 wire _15698_;
 wire _15699_;
 wire _15700_;
 wire _15701_;
 wire _15702_;
 wire _15703_;
 wire _15704_;
 wire _15705_;
 wire _15706_;
 wire _15707_;
 wire _15708_;
 wire _15709_;
 wire _15710_;
 wire _15711_;
 wire _15712_;
 wire _15713_;
 wire _15714_;
 wire _15715_;
 wire _15716_;
 wire _15717_;
 wire _15718_;
 wire _15719_;
 wire _15720_;
 wire _15721_;
 wire _15722_;
 wire _15723_;
 wire _15724_;
 wire _15725_;
 wire _15726_;
 wire _15727_;
 wire _15728_;
 wire _15729_;
 wire _15730_;
 wire _15731_;
 wire _15732_;
 wire _15733_;
 wire _15734_;
 wire _15735_;
 wire _15736_;
 wire _15737_;
 wire _15738_;
 wire _15739_;
 wire _15740_;
 wire _15741_;
 wire _15742_;
 wire _15743_;
 wire _15744_;
 wire _15745_;
 wire _15746_;
 wire _15747_;
 wire _15748_;
 wire _15749_;
 wire _15750_;
 wire _15751_;
 wire _15752_;
 wire _15753_;
 wire _15754_;
 wire _15755_;
 wire _15756_;
 wire _15757_;
 wire _15758_;
 wire net1150;
 wire _15760_;
 wire _15761_;
 wire _15762_;
 wire _15763_;
 wire _15764_;
 wire _15765_;
 wire _15766_;
 wire _15767_;
 wire _15768_;
 wire _15769_;
 wire _15770_;
 wire _15771_;
 wire _15772_;
 wire _15773_;
 wire net1149;
 wire _15775_;
 wire _15776_;
 wire _15777_;
 wire _15778_;
 wire net1148;
 wire _15780_;
 wire _15781_;
 wire _15782_;
 wire net1147;
 wire _15784_;
 wire _15785_;
 wire _15786_;
 wire _15787_;
 wire _15788_;
 wire _15789_;
 wire _15790_;
 wire _15791_;
 wire _15792_;
 wire _15793_;
 wire _15794_;
 wire _15795_;
 wire _15796_;
 wire _15797_;
 wire _15798_;
 wire _15799_;
 wire _15800_;
 wire _15801_;
 wire _15802_;
 wire _15803_;
 wire _15804_;
 wire _15805_;
 wire _15806_;
 wire _15807_;
 wire _15808_;
 wire _15809_;
 wire _15810_;
 wire _15811_;
 wire _15812_;
 wire _15813_;
 wire _15814_;
 wire _15815_;
 wire _15816_;
 wire _15817_;
 wire _15818_;
 wire _15819_;
 wire _15820_;
 wire _15821_;
 wire _15822_;
 wire _15823_;
 wire _15824_;
 wire _15825_;
 wire _15826_;
 wire _15827_;
 wire _15828_;
 wire _15829_;
 wire _15830_;
 wire _15831_;
 wire _15832_;
 wire _15833_;
 wire _15834_;
 wire _15835_;
 wire _15836_;
 wire _15837_;
 wire _15838_;
 wire _15839_;
 wire _15840_;
 wire _15841_;
 wire _15842_;
 wire _15843_;
 wire _15844_;
 wire _15845_;
 wire _15846_;
 wire _15847_;
 wire _15848_;
 wire _15849_;
 wire _15850_;
 wire _15851_;
 wire _15852_;
 wire _15853_;
 wire _15854_;
 wire _15855_;
 wire _15856_;
 wire _15857_;
 wire _15858_;
 wire _15859_;
 wire _15860_;
 wire _15861_;
 wire _15862_;
 wire _15863_;
 wire _15864_;
 wire _15865_;
 wire _15866_;
 wire _15867_;
 wire _15868_;
 wire _15869_;
 wire _15870_;
 wire _15871_;
 wire _15872_;
 wire _15873_;
 wire _15874_;
 wire _15875_;
 wire _15876_;
 wire _15877_;
 wire _15878_;
 wire _15879_;
 wire _15880_;
 wire _15881_;
 wire _15882_;
 wire _15883_;
 wire _15884_;
 wire _15885_;
 wire _15886_;
 wire _15887_;
 wire _15888_;
 wire _15889_;
 wire _15890_;
 wire net1144;
 wire _15892_;
 wire _15893_;
 wire net1143;
 wire net1142;
 wire net1141;
 wire _15897_;
 wire net1140;
 wire _15899_;
 wire _15900_;
 wire net1139;
 wire _15902_;
 wire net1138;
 wire _15904_;
 wire _15905_;
 wire _15906_;
 wire _15907_;
 wire net1137;
 wire _15909_;
 wire net1136;
 wire _15911_;
 wire _15912_;
 wire net1135;
 wire net1134;
 wire _15915_;
 wire net1133;
 wire _15917_;
 wire net1132;
 wire _15919_;
 wire net1131;
 wire _15921_;
 wire _15922_;
 wire net1130;
 wire _15924_;
 wire net1129;
 wire _15926_;
 wire _15927_;
 wire _15928_;
 wire _15929_;
 wire _15930_;
 wire _15931_;
 wire _15932_;
 wire _15933_;
 wire net1128;
 wire net1127;
 wire _15936_;
 wire _15937_;
 wire _15938_;
 wire _15939_;
 wire _15940_;
 wire _15941_;
 wire _15942_;
 wire _15943_;
 wire _15944_;
 wire net1126;
 wire _15946_;
 wire net1125;
 wire net1124;
 wire _15949_;
 wire _15950_;
 wire net1123;
 wire _15952_;
 wire _15953_;
 wire _15954_;
 wire _15955_;
 wire _15956_;
 wire _15957_;
 wire net1122;
 wire _15959_;
 wire _15960_;
 wire _15961_;
 wire _15962_;
 wire _15963_;
 wire _15964_;
 wire _15965_;
 wire _15966_;
 wire _15967_;
 wire _15968_;
 wire _15969_;
 wire _15970_;
 wire _15971_;
 wire _15972_;
 wire _15973_;
 wire _15974_;
 wire _15975_;
 wire _15976_;
 wire _15977_;
 wire _15978_;
 wire _15979_;
 wire _15980_;
 wire _15981_;
 wire _15982_;
 wire _15983_;
 wire _15984_;
 wire _15985_;
 wire _15986_;
 wire _15987_;
 wire _15988_;
 wire _15989_;
 wire _15990_;
 wire _15991_;
 wire _15992_;
 wire _15993_;
 wire _15994_;
 wire _15995_;
 wire _15996_;
 wire _15997_;
 wire _15998_;
 wire _15999_;
 wire _16000_;
 wire _16001_;
 wire _16002_;
 wire _16003_;
 wire _16004_;
 wire _16005_;
 wire _16006_;
 wire _16007_;
 wire _16008_;
 wire _16009_;
 wire _16010_;
 wire _16011_;
 wire _16012_;
 wire _16013_;
 wire _16014_;
 wire _16015_;
 wire _16016_;
 wire _16017_;
 wire _16018_;
 wire _16019_;
 wire _16020_;
 wire _16021_;
 wire _16022_;
 wire _16023_;
 wire _16024_;
 wire _16025_;
 wire net1120;
 wire _16027_;
 wire _16028_;
 wire _16029_;
 wire _16030_;
 wire _16031_;
 wire net1119;
 wire _16033_;
 wire _16034_;
 wire net1118;
 wire _16036_;
 wire _16037_;
 wire _16038_;
 wire _16039_;
 wire net1117;
 wire _16041_;
 wire _16042_;
 wire _16043_;
 wire _16044_;
 wire _16045_;
 wire _16046_;
 wire _16047_;
 wire _16048_;
 wire _16049_;
 wire _16050_;
 wire _16051_;
 wire net1116;
 wire _16053_;
 wire net1115;
 wire _16055_;
 wire _16056_;
 wire _16057_;
 wire _16058_;
 wire _16059_;
 wire _16060_;
 wire _16061_;
 wire _16062_;
 wire _16063_;
 wire net1114;
 wire _16065_;
 wire _16066_;
 wire _16067_;
 wire _16068_;
 wire _16069_;
 wire _16070_;
 wire _16071_;
 wire _16072_;
 wire _16073_;
 wire _16074_;
 wire _16075_;
 wire _16076_;
 wire _16077_;
 wire _16078_;
 wire _16079_;
 wire net1113;
 wire _16081_;
 wire _16082_;
 wire _16083_;
 wire _16084_;
 wire _16085_;
 wire _16086_;
 wire _16087_;
 wire _16088_;
 wire _16089_;
 wire _16090_;
 wire _16091_;
 wire _16092_;
 wire _16093_;
 wire _16094_;
 wire _16095_;
 wire _16096_;
 wire _16097_;
 wire _16098_;
 wire _16099_;
 wire _16100_;
 wire _16101_;
 wire _16102_;
 wire _16103_;
 wire _16104_;
 wire _16105_;
 wire _16106_;
 wire _16107_;
 wire _16108_;
 wire _16109_;
 wire _16110_;
 wire _16111_;
 wire _16112_;
 wire _16113_;
 wire _16114_;
 wire _16115_;
 wire _16116_;
 wire _16117_;
 wire _16118_;
 wire _16119_;
 wire _16120_;
 wire _16121_;
 wire _16122_;
 wire _16123_;
 wire _16124_;
 wire _16125_;
 wire _16126_;
 wire _16127_;
 wire _16128_;
 wire _16129_;
 wire _16130_;
 wire _16131_;
 wire _16132_;
 wire _16133_;
 wire _16134_;
 wire _16135_;
 wire _16136_;
 wire _16137_;
 wire _16138_;
 wire net1112;
 wire _16140_;
 wire _16141_;
 wire _16142_;
 wire _16143_;
 wire _16144_;
 wire _16145_;
 wire _16146_;
 wire _16147_;
 wire _16148_;
 wire _16149_;
 wire _16150_;
 wire _16151_;
 wire net1110;
 wire _16153_;
 wire net1109;
 wire _16155_;
 wire _16156_;
 wire _16157_;
 wire _16158_;
 wire _16159_;
 wire _16160_;
 wire _16161_;
 wire _16162_;
 wire _16163_;
 wire net1108;
 wire _16165_;
 wire _16166_;
 wire _16167_;
 wire _16168_;
 wire _16169_;
 wire _16170_;
 wire _16171_;
 wire _16172_;
 wire _16173_;
 wire _16174_;
 wire _16175_;
 wire _16176_;
 wire _16177_;
 wire _16178_;
 wire _16179_;
 wire _16180_;
 wire _16181_;
 wire _16182_;
 wire _16183_;
 wire _16184_;
 wire _16185_;
 wire _16186_;
 wire _16187_;
 wire _16188_;
 wire _16189_;
 wire _16190_;
 wire _16191_;
 wire _16192_;
 wire net1107;
 wire net1106;
 wire _16195_;
 wire net1105;
 wire _16197_;
 wire _16198_;
 wire net1104;
 wire _16200_;
 wire _16201_;
 wire _16202_;
 wire _16203_;
 wire _16204_;
 wire _16205_;
 wire _16206_;
 wire _16207_;
 wire _16208_;
 wire _16209_;
 wire _16210_;
 wire _16211_;
 wire _16212_;
 wire _16213_;
 wire _16214_;
 wire _16215_;
 wire _16216_;
 wire _16217_;
 wire net1103;
 wire _16219_;
 wire _16220_;
 wire _16221_;
 wire _16222_;
 wire _16223_;
 wire _16224_;
 wire net1102;
 wire _16226_;
 wire _16227_;
 wire _16228_;
 wire _16229_;
 wire _16230_;
 wire _16231_;
 wire _16232_;
 wire _16233_;
 wire _16234_;
 wire _16235_;
 wire _16236_;
 wire _16237_;
 wire _16238_;
 wire _16239_;
 wire _16240_;
 wire _16241_;
 wire _16242_;
 wire _16243_;
 wire _16244_;
 wire _16245_;
 wire _16246_;
 wire _16247_;
 wire _16248_;
 wire _16249_;
 wire _16250_;
 wire _16251_;
 wire _16252_;
 wire _16253_;
 wire _16254_;
 wire _16255_;
 wire _16256_;
 wire _16257_;
 wire _16258_;
 wire _16259_;
 wire _16260_;
 wire _16261_;
 wire _16262_;
 wire _16263_;
 wire net1100;
 wire _16265_;
 wire _16266_;
 wire _16267_;
 wire _16268_;
 wire _16269_;
 wire _16270_;
 wire _16271_;
 wire _16272_;
 wire _16273_;
 wire _16274_;
 wire _16275_;
 wire _16276_;
 wire _16277_;
 wire _16278_;
 wire _16279_;
 wire _16280_;
 wire _16281_;
 wire _16282_;
 wire _16283_;
 wire _16284_;
 wire _16285_;
 wire _16286_;
 wire _16287_;
 wire _16288_;
 wire _16289_;
 wire _16290_;
 wire _16291_;
 wire _16292_;
 wire _16293_;
 wire _16294_;
 wire _16295_;
 wire _16296_;
 wire _16297_;
 wire _16298_;
 wire _16299_;
 wire _16300_;
 wire _16301_;
 wire _16302_;
 wire _16303_;
 wire _16304_;
 wire _16305_;
 wire _16306_;
 wire _16307_;
 wire _16308_;
 wire _16309_;
 wire net1099;
 wire _16311_;
 wire _16312_;
 wire _16313_;
 wire _16314_;
 wire _16315_;
 wire _16316_;
 wire _16317_;
 wire _16318_;
 wire _16319_;
 wire _16320_;
 wire _16321_;
 wire _16322_;
 wire _16323_;
 wire _16324_;
 wire net1098;
 wire _16326_;
 wire net1097;
 wire _16328_;
 wire _16329_;
 wire _16330_;
 wire _16331_;
 wire net1096;
 wire _16333_;
 wire _16334_;
 wire _16335_;
 wire _16336_;
 wire _16337_;
 wire _16338_;
 wire _16339_;
 wire _16340_;
 wire _16341_;
 wire _16342_;
 wire _16343_;
 wire _16344_;
 wire _16345_;
 wire _16346_;
 wire _16347_;
 wire _16348_;
 wire _16349_;
 wire _16350_;
 wire _16351_;
 wire _16352_;
 wire _16353_;
 wire _16354_;
 wire _16355_;
 wire _16356_;
 wire _16357_;
 wire _16358_;
 wire _16359_;
 wire _16360_;
 wire _16361_;
 wire _16362_;
 wire _16363_;
 wire _16364_;
 wire net1095;
 wire _16366_;
 wire _16367_;
 wire _16368_;
 wire _16369_;
 wire _16370_;
 wire _16371_;
 wire _16372_;
 wire _16373_;
 wire _16374_;
 wire _16375_;
 wire _16376_;
 wire _16377_;
 wire _16378_;
 wire _16379_;
 wire net1094;
 wire _16381_;
 wire _16382_;
 wire _16383_;
 wire _16384_;
 wire _16385_;
 wire _16386_;
 wire _16387_;
 wire _16388_;
 wire _16389_;
 wire _16390_;
 wire _16391_;
 wire _16392_;
 wire _16393_;
 wire _16394_;
 wire _16395_;
 wire _16396_;
 wire _16397_;
 wire _16398_;
 wire _16399_;
 wire _16400_;
 wire _16401_;
 wire _16402_;
 wire _16403_;
 wire _16404_;
 wire _16405_;
 wire net1092;
 wire _16407_;
 wire _16408_;
 wire _16409_;
 wire _16410_;
 wire _16411_;
 wire net1091;
 wire _16413_;
 wire _16414_;
 wire _16415_;
 wire _16416_;
 wire _16417_;
 wire _16418_;
 wire _16419_;
 wire _16420_;
 wire _16421_;
 wire _16422_;
 wire _16423_;
 wire _16424_;
 wire _16425_;
 wire _16426_;
 wire _16427_;
 wire _16428_;
 wire _16429_;
 wire _16430_;
 wire _16431_;
 wire _16432_;
 wire _16433_;
 wire _16434_;
 wire _16435_;
 wire _16436_;
 wire _16437_;
 wire _16438_;
 wire _16439_;
 wire _16440_;
 wire _16441_;
 wire _16442_;
 wire net1090;
 wire _16444_;
 wire _16445_;
 wire _16446_;
 wire _16447_;
 wire _16448_;
 wire _16449_;
 wire _16450_;
 wire _16451_;
 wire _16452_;
 wire _16453_;
 wire _16454_;
 wire _16455_;
 wire _16456_;
 wire _16457_;
 wire net1089;
 wire _16459_;
 wire net1088;
 wire _16461_;
 wire _16462_;
 wire _16463_;
 wire _16464_;
 wire _16465_;
 wire _16466_;
 wire _16467_;
 wire _16468_;
 wire _16469_;
 wire _16470_;
 wire _16471_;
 wire _16472_;
 wire _16473_;
 wire _16474_;
 wire _16475_;
 wire _16476_;
 wire _16477_;
 wire _16478_;
 wire _16479_;
 wire _16480_;
 wire _16481_;
 wire _16482_;
 wire _16483_;
 wire _16484_;
 wire _16485_;
 wire _16486_;
 wire _16487_;
 wire _16488_;
 wire _16489_;
 wire _16490_;
 wire _16491_;
 wire _16492_;
 wire _16493_;
 wire _16494_;
 wire _16495_;
 wire _16496_;
 wire _16497_;
 wire _16498_;
 wire _16499_;
 wire _16500_;
 wire _16501_;
 wire _16502_;
 wire _16503_;
 wire _16504_;
 wire _16505_;
 wire _16506_;
 wire _16507_;
 wire _16508_;
 wire _16509_;
 wire _16510_;
 wire _16511_;
 wire _16512_;
 wire _16513_;
 wire _16514_;
 wire _16515_;
 wire _16516_;
 wire _16517_;
 wire _16518_;
 wire _16519_;
 wire _16520_;
 wire _16521_;
 wire _16522_;
 wire _16523_;
 wire _16524_;
 wire _16525_;
 wire _16526_;
 wire _16527_;
 wire _16528_;
 wire _16529_;
 wire _16530_;
 wire _16531_;
 wire _16532_;
 wire _16533_;
 wire _16534_;
 wire _16535_;
 wire _16536_;
 wire _16537_;
 wire _16538_;
 wire _16539_;
 wire _16540_;
 wire _16541_;
 wire _16542_;
 wire _16543_;
 wire _16544_;
 wire _16545_;
 wire _16546_;
 wire _16547_;
 wire _16548_;
 wire _16549_;
 wire _16550_;
 wire _16551_;
 wire _16552_;
 wire _16553_;
 wire _16554_;
 wire _16555_;
 wire _16556_;
 wire _16557_;
 wire _16558_;
 wire _16559_;
 wire _16560_;
 wire _16561_;
 wire _16562_;
 wire _16563_;
 wire _16564_;
 wire _16565_;
 wire _16566_;
 wire _16567_;
 wire _16568_;
 wire net1087;
 wire _16570_;
 wire _16571_;
 wire _16572_;
 wire _16573_;
 wire _16574_;
 wire _16575_;
 wire _16576_;
 wire _16577_;
 wire _16578_;
 wire _16579_;
 wire _16580_;
 wire _16581_;
 wire _16582_;
 wire _16583_;
 wire _16584_;
 wire _16585_;
 wire _16586_;
 wire _16587_;
 wire _16588_;
 wire _16589_;
 wire _16590_;
 wire _16591_;
 wire _16592_;
 wire _16593_;
 wire _16594_;
 wire _16595_;
 wire _16596_;
 wire _16597_;
 wire _16598_;
 wire _16599_;
 wire _16600_;
 wire _16601_;
 wire _16602_;
 wire _16603_;
 wire _16604_;
 wire _16605_;
 wire _16606_;
 wire _16607_;
 wire _16608_;
 wire _16609_;
 wire _16610_;
 wire _16611_;
 wire _16612_;
 wire _16613_;
 wire _16614_;
 wire _16615_;
 wire _16616_;
 wire _16617_;
 wire _16618_;
 wire _16619_;
 wire _16620_;
 wire _16621_;
 wire _16622_;
 wire _16623_;
 wire _16624_;
 wire _16625_;
 wire _16626_;
 wire _16627_;
 wire _16628_;
 wire _16629_;
 wire _16630_;
 wire _16631_;
 wire _16632_;
 wire _16633_;
 wire _16634_;
 wire _16635_;
 wire _16636_;
 wire _16637_;
 wire _16638_;
 wire _16639_;
 wire _16640_;
 wire _16641_;
 wire _16642_;
 wire _16643_;
 wire _16644_;
 wire _16645_;
 wire _16646_;
 wire _16647_;
 wire _16648_;
 wire _16649_;
 wire _16650_;
 wire _16651_;
 wire _16652_;
 wire _16653_;
 wire _16654_;
 wire _16655_;
 wire _16656_;
 wire _16657_;
 wire _16658_;
 wire _16659_;
 wire _16660_;
 wire _16661_;
 wire _16662_;
 wire _16663_;
 wire _16664_;
 wire _16665_;
 wire _16666_;
 wire _16667_;
 wire _16668_;
 wire _16669_;
 wire _16670_;
 wire _16671_;
 wire _16672_;
 wire _16673_;
 wire _16674_;
 wire _16675_;
 wire _16676_;
 wire _16677_;
 wire _16678_;
 wire _16679_;
 wire _16680_;
 wire _16681_;
 wire _16682_;
 wire _16683_;
 wire _16684_;
 wire _16685_;
 wire _16686_;
 wire _16687_;
 wire _16688_;
 wire _16689_;
 wire _16690_;
 wire _16691_;
 wire _16692_;
 wire _16693_;
 wire _16694_;
 wire _16695_;
 wire _16696_;
 wire _16697_;
 wire _16698_;
 wire _16699_;
 wire _16700_;
 wire _16701_;
 wire _16702_;
 wire _16703_;
 wire _16704_;
 wire _16705_;
 wire _16706_;
 wire _16707_;
 wire _16708_;
 wire _16709_;
 wire _16710_;
 wire _16711_;
 wire _16712_;
 wire _16713_;
 wire _16714_;
 wire _16715_;
 wire _16716_;
 wire _16717_;
 wire _16718_;
 wire _16719_;
 wire net1402;
 wire _16721_;
 wire _16722_;
 wire _16723_;
 wire _16724_;
 wire _16725_;
 wire _16726_;
 wire _16727_;
 wire _16728_;
 wire _16729_;
 wire _16730_;
 wire _16731_;
 wire _16732_;
 wire _16733_;
 wire _16734_;
 wire _16735_;
 wire _16736_;
 wire _16737_;
 wire _16738_;
 wire _16739_;
 wire _16740_;
 wire _16741_;
 wire _16742_;
 wire _16743_;
 wire _16744_;
 wire _16745_;
 wire _16746_;
 wire _16747_;
 wire _16748_;
 wire _16749_;
 wire _16750_;
 wire _16751_;
 wire _16752_;
 wire _16753_;
 wire _16754_;
 wire _16755_;
 wire _16756_;
 wire _16757_;
 wire _16758_;
 wire _16759_;
 wire _16760_;
 wire _16761_;
 wire _16762_;
 wire _16763_;
 wire _16764_;
 wire _16765_;
 wire _16766_;
 wire _16767_;
 wire _16768_;
 wire _16769_;
 wire _16770_;
 wire _16771_;
 wire _16772_;
 wire _16773_;
 wire _16774_;
 wire _16775_;
 wire _16776_;
 wire _16777_;
 wire _16778_;
 wire _16779_;
 wire _16780_;
 wire _16781_;
 wire _16782_;
 wire _16783_;
 wire _16784_;
 wire _16785_;
 wire _16786_;
 wire _16787_;
 wire _16788_;
 wire _16789_;
 wire _16790_;
 wire _16791_;
 wire _16792_;
 wire _16793_;
 wire _16794_;
 wire _16795_;
 wire _16796_;
 wire _16797_;
 wire _16798_;
 wire _16799_;
 wire _16800_;
 wire _16801_;
 wire _16802_;
 wire _16803_;
 wire _16804_;
 wire _16805_;
 wire _16806_;
 wire _16807_;
 wire _16808_;
 wire _16809_;
 wire _16810_;
 wire _16811_;
 wire _16812_;
 wire _16813_;
 wire _16814_;
 wire _16815_;
 wire _16816_;
 wire _16817_;
 wire _16818_;
 wire _16819_;
 wire _16820_;
 wire _16821_;
 wire _16822_;
 wire _16823_;
 wire _16824_;
 wire _16825_;
 wire _16826_;
 wire _16827_;
 wire _16828_;
 wire _16829_;
 wire _16830_;
 wire _16831_;
 wire _16832_;
 wire _16833_;
 wire _16834_;
 wire _16835_;
 wire _16836_;
 wire _16837_;
 wire _16838_;
 wire _16839_;
 wire _16840_;
 wire _16841_;
 wire _16842_;
 wire _16843_;
 wire _16844_;
 wire _16845_;
 wire _16846_;
 wire _16847_;
 wire _16848_;
 wire _16849_;
 wire _16850_;
 wire _16851_;
 wire _16852_;
 wire _16853_;
 wire _16854_;
 wire _16855_;
 wire _16856_;
 wire _16857_;
 wire _16858_;
 wire _16859_;
 wire _16860_;
 wire _16861_;
 wire _16862_;
 wire _16863_;
 wire _16864_;
 wire _16865_;
 wire _16866_;
 wire _16867_;
 wire _16868_;
 wire _16869_;
 wire _16870_;
 wire _16871_;
 wire _16872_;
 wire _16873_;
 wire _16874_;
 wire _16875_;
 wire _16876_;
 wire _16877_;
 wire _16878_;
 wire _16879_;
 wire _16880_;
 wire _16881_;
 wire _16882_;
 wire _16883_;
 wire _16884_;
 wire _16885_;
 wire _16886_;
 wire _16887_;
 wire _16888_;
 wire _16889_;
 wire _16890_;
 wire _16891_;
 wire _16892_;
 wire _16893_;
 wire _16894_;
 wire _16895_;
 wire _16896_;
 wire _16897_;
 wire _16898_;
 wire _16899_;
 wire _16900_;
 wire _16901_;
 wire _16902_;
 wire _16903_;
 wire _16904_;
 wire _16905_;
 wire _16906_;
 wire _16907_;
 wire _16908_;
 wire _16909_;
 wire _16910_;
 wire _16911_;
 wire _16912_;
 wire _16913_;
 wire _16914_;
 wire _16915_;
 wire _16916_;
 wire _16917_;
 wire _16918_;
 wire _16919_;
 wire _16920_;
 wire _16921_;
 wire _16922_;
 wire _16923_;
 wire _16924_;
 wire _16925_;
 wire _16926_;
 wire _16927_;
 wire _16928_;
 wire _16929_;
 wire _16930_;
 wire _16931_;
 wire _16932_;
 wire _16933_;
 wire _16934_;
 wire _16935_;
 wire _16936_;
 wire _16937_;
 wire _16938_;
 wire _16939_;
 wire _16940_;
 wire _16941_;
 wire _16942_;
 wire _16943_;
 wire _16944_;
 wire _16945_;
 wire _16946_;
 wire _16947_;
 wire _16948_;
 wire _16949_;
 wire _16950_;
 wire _16951_;
 wire _16952_;
 wire _16953_;
 wire _16954_;
 wire _16955_;
 wire _16956_;
 wire _16957_;
 wire _16958_;
 wire _16959_;
 wire _16960_;
 wire _16961_;
 wire _16962_;
 wire _16963_;
 wire _16964_;
 wire _16965_;
 wire _16966_;
 wire _16967_;
 wire _16968_;
 wire _16969_;
 wire _16970_;
 wire _16971_;
 wire _16972_;
 wire _16973_;
 wire _16974_;
 wire _16975_;
 wire _16976_;
 wire _16977_;
 wire _16978_;
 wire _16979_;
 wire _16980_;
 wire _16981_;
 wire _16982_;
 wire _16983_;
 wire _16984_;
 wire _16985_;
 wire _16986_;
 wire _16987_;
 wire _16988_;
 wire _16989_;
 wire _16990_;
 wire _16991_;
 wire _16992_;
 wire _16993_;
 wire _16994_;
 wire _16995_;
 wire _16996_;
 wire _16997_;
 wire _16998_;
 wire _16999_;
 wire _17000_;
 wire _17001_;
 wire _17002_;
 wire _17003_;
 wire _17004_;
 wire _17005_;
 wire _17006_;
 wire _17007_;
 wire _17008_;
 wire _17009_;
 wire _17010_;
 wire _17011_;
 wire _17012_;
 wire _17013_;
 wire _17014_;
 wire _17015_;
 wire _17016_;
 wire _17017_;
 wire _17018_;
 wire _17019_;
 wire _17020_;
 wire _17021_;
 wire _17022_;
 wire _17023_;
 wire _17024_;
 wire _17025_;
 wire _17026_;
 wire _17027_;
 wire _17028_;
 wire _17029_;
 wire _17030_;
 wire _17031_;
 wire _17032_;
 wire _17033_;
 wire _17034_;
 wire _17035_;
 wire _17036_;
 wire _17037_;
 wire _17038_;
 wire _17039_;
 wire _17040_;
 wire _17041_;
 wire _17042_;
 wire _17043_;
 wire _17044_;
 wire _17045_;
 wire _17046_;
 wire _17047_;
 wire _17048_;
 wire _17049_;
 wire _17050_;
 wire _17051_;
 wire _17052_;
 wire _17053_;
 wire _17054_;
 wire _17055_;
 wire _17056_;
 wire _17057_;
 wire _17058_;
 wire _17059_;
 wire _17060_;
 wire _17061_;
 wire _17062_;
 wire _17063_;
 wire _17064_;
 wire _17065_;
 wire _17066_;
 wire _17067_;
 wire _17068_;
 wire _17069_;
 wire _17070_;
 wire _17071_;
 wire _17072_;
 wire _17073_;
 wire _17074_;
 wire _17075_;
 wire _17076_;
 wire _17077_;
 wire _17078_;
 wire _17079_;
 wire _17080_;
 wire _17081_;
 wire _17082_;
 wire _17083_;
 wire _17084_;
 wire _17085_;
 wire _17086_;
 wire _17087_;
 wire _17088_;
 wire _17089_;
 wire _17090_;
 wire _17091_;
 wire _17092_;
 wire _17093_;
 wire _17094_;
 wire _17095_;
 wire _17096_;
 wire _17097_;
 wire _17098_;
 wire _17099_;
 wire _17100_;
 wire _17101_;
 wire _17102_;
 wire _17103_;
 wire _17104_;
 wire _17105_;
 wire _17106_;
 wire _17107_;
 wire _17108_;
 wire _17109_;
 wire _17110_;
 wire _17111_;
 wire _17112_;
 wire _17113_;
 wire _17114_;
 wire _17115_;
 wire _17116_;
 wire _17117_;
 wire _17118_;
 wire _17119_;
 wire _17120_;
 wire net958;
 wire _17122_;
 wire _17123_;
 wire _17124_;
 wire _17125_;
 wire _17126_;
 wire _17127_;
 wire _17128_;
 wire _17129_;
 wire _17130_;
 wire _17131_;
 wire _17132_;
 wire _17133_;
 wire _17134_;
 wire _17135_;
 wire _17136_;
 wire _17137_;
 wire _17138_;
 wire _17139_;
 wire _17140_;
 wire _17141_;
 wire _17142_;
 wire _17143_;
 wire _17144_;
 wire _17145_;
 wire _17146_;
 wire _17147_;
 wire _17148_;
 wire _17149_;
 wire _17150_;
 wire _17151_;
 wire _17152_;
 wire _17153_;
 wire _17154_;
 wire _17155_;
 wire _17156_;
 wire _17157_;
 wire _17158_;
 wire _17159_;
 wire _17160_;
 wire _17161_;
 wire _17162_;
 wire _17163_;
 wire _17164_;
 wire _17165_;
 wire _17166_;
 wire _17167_;
 wire _17168_;
 wire _17169_;
 wire _17170_;
 wire _17171_;
 wire _17172_;
 wire _17173_;
 wire _17174_;
 wire _17175_;
 wire _17176_;
 wire _17177_;
 wire _17178_;
 wire _17179_;
 wire _17180_;
 wire _17181_;
 wire _17182_;
 wire _17183_;
 wire _17184_;
 wire _17185_;
 wire _17186_;
 wire _17187_;
 wire _17188_;
 wire _17189_;
 wire _17190_;
 wire _17191_;
 wire _17192_;
 wire _17193_;
 wire _17194_;
 wire _17195_;
 wire _17196_;
 wire _17197_;
 wire _17198_;
 wire _17199_;
 wire _17200_;
 wire _17201_;
 wire _17202_;
 wire _17203_;
 wire _17204_;
 wire _17205_;
 wire _17206_;
 wire _17207_;
 wire _17208_;
 wire _17209_;
 wire _17210_;
 wire _17211_;
 wire _17212_;
 wire _17213_;
 wire _17214_;
 wire _17215_;
 wire _17216_;
 wire _17217_;
 wire _17218_;
 wire _17219_;
 wire _17220_;
 wire _17221_;
 wire _17222_;
 wire _17223_;
 wire _17224_;
 wire _17225_;
 wire _17226_;
 wire _17227_;
 wire _17228_;
 wire _17229_;
 wire _17230_;
 wire _17231_;
 wire _17232_;
 wire _17233_;
 wire _17234_;
 wire _17235_;
 wire _17236_;
 wire _17237_;
 wire _17238_;
 wire _17239_;
 wire _17240_;
 wire _17241_;
 wire _17242_;
 wire _17243_;
 wire _17244_;
 wire _17245_;
 wire _17246_;
 wire _17247_;
 wire _17248_;
 wire _17249_;
 wire _17250_;
 wire _17251_;
 wire _17252_;
 wire _17253_;
 wire _17254_;
 wire _17255_;
 wire _17256_;
 wire _17257_;
 wire _17258_;
 wire _17259_;
 wire _17260_;
 wire _17261_;
 wire _17262_;
 wire _17263_;
 wire _17264_;
 wire _17265_;
 wire _17266_;
 wire _17267_;
 wire _17268_;
 wire _17269_;
 wire _17270_;
 wire _17271_;
 wire _17272_;
 wire _17273_;
 wire _17274_;
 wire _17275_;
 wire _17276_;
 wire _17277_;
 wire _17278_;
 wire _17279_;
 wire _17280_;
 wire _17281_;
 wire _17282_;
 wire _17283_;
 wire _17284_;
 wire _17285_;
 wire _17286_;
 wire _17287_;
 wire _17288_;
 wire _17289_;
 wire _17290_;
 wire _17291_;
 wire _17292_;
 wire _17293_;
 wire _17294_;
 wire _17295_;
 wire _17296_;
 wire _17297_;
 wire _17298_;
 wire _17299_;
 wire _17300_;
 wire _17301_;
 wire _17302_;
 wire _17303_;
 wire _17304_;
 wire _17305_;
 wire _17306_;
 wire _17307_;
 wire _17308_;
 wire _17309_;
 wire _17310_;
 wire _17311_;
 wire _17312_;
 wire _17313_;
 wire _17314_;
 wire _17315_;
 wire _17316_;
 wire _17317_;
 wire _17318_;
 wire _17319_;
 wire _17320_;
 wire _17321_;
 wire _17322_;
 wire _17323_;
 wire _17324_;
 wire _17325_;
 wire _17326_;
 wire _17327_;
 wire _17328_;
 wire _17329_;
 wire _17330_;
 wire _17331_;
 wire _17332_;
 wire _17333_;
 wire _17334_;
 wire _17335_;
 wire _17336_;
 wire _17337_;
 wire _17338_;
 wire _17339_;
 wire _17340_;
 wire _17341_;
 wire _17342_;
 wire _17343_;
 wire _17344_;
 wire _17345_;
 wire _17346_;
 wire _17347_;
 wire _17348_;
 wire _17349_;
 wire _17350_;
 wire _17351_;
 wire _17352_;
 wire _17353_;
 wire _17354_;
 wire _17355_;
 wire _17356_;
 wire _17357_;
 wire _17358_;
 wire _17359_;
 wire _17360_;
 wire _17361_;
 wire _17362_;
 wire _17363_;
 wire _17364_;
 wire _17365_;
 wire _17366_;
 wire _17367_;
 wire _17368_;
 wire _17369_;
 wire _17370_;
 wire _17371_;
 wire _17372_;
 wire _17373_;
 wire _17374_;
 wire _17375_;
 wire _17376_;
 wire _17377_;
 wire _17378_;
 wire _17379_;
 wire _17380_;
 wire _17381_;
 wire _17382_;
 wire _17383_;
 wire _17384_;
 wire _17385_;
 wire _17386_;
 wire _17387_;
 wire _17388_;
 wire _17389_;
 wire _17390_;
 wire _17391_;
 wire _17392_;
 wire _17393_;
 wire _17394_;
 wire _17395_;
 wire _17396_;
 wire _17397_;
 wire _17398_;
 wire _17399_;
 wire _17400_;
 wire _17401_;
 wire _17402_;
 wire _17403_;
 wire _17404_;
 wire _17405_;
 wire _17406_;
 wire _17407_;
 wire _17408_;
 wire _17409_;
 wire _17410_;
 wire _17411_;
 wire _17412_;
 wire _17413_;
 wire _17414_;
 wire _17415_;
 wire _17416_;
 wire _17417_;
 wire _17418_;
 wire _17419_;
 wire _17420_;
 wire _17421_;
 wire _17422_;
 wire _17423_;
 wire _17424_;
 wire _17425_;
 wire _17426_;
 wire _17427_;
 wire _17428_;
 wire _17429_;
 wire _17430_;
 wire _17431_;
 wire _17432_;
 wire _17433_;
 wire _17434_;
 wire _17435_;
 wire _17436_;
 wire _17437_;
 wire _17438_;
 wire _17439_;
 wire _17440_;
 wire _17441_;
 wire _17442_;
 wire _17443_;
 wire _17444_;
 wire _17445_;
 wire _17446_;
 wire _17447_;
 wire _17448_;
 wire _17449_;
 wire _17450_;
 wire _17451_;
 wire _17452_;
 wire _17453_;
 wire _17454_;
 wire _17455_;
 wire _17456_;
 wire _17457_;
 wire _17458_;
 wire _17459_;
 wire _17460_;
 wire _17461_;
 wire _17462_;
 wire _17463_;
 wire _17464_;
 wire _17465_;
 wire _17466_;
 wire _17467_;
 wire _17468_;
 wire _17469_;
 wire _17470_;
 wire _17471_;
 wire _17472_;
 wire _17473_;
 wire _17474_;
 wire _17475_;
 wire _17476_;
 wire _17477_;
 wire _17478_;
 wire _17479_;
 wire _17480_;
 wire _17481_;
 wire _17482_;
 wire _17483_;
 wire _17484_;
 wire _17485_;
 wire _17486_;
 wire _17487_;
 wire _17488_;
 wire _17489_;
 wire _17490_;
 wire _17491_;
 wire _17492_;
 wire _17493_;
 wire _17494_;
 wire _17495_;
 wire _17496_;
 wire _17497_;
 wire _17498_;
 wire _17499_;
 wire _17500_;
 wire _17501_;
 wire _17502_;
 wire _17503_;
 wire _17504_;
 wire _17505_;
 wire _17506_;
 wire _17507_;
 wire _17508_;
 wire _17509_;
 wire _17510_;
 wire _17511_;
 wire _17512_;
 wire _17513_;
 wire _17514_;
 wire _17515_;
 wire _17516_;
 wire _17517_;
 wire _17518_;
 wire _17519_;
 wire _17520_;
 wire _17521_;
 wire _17522_;
 wire _17523_;
 wire _17524_;
 wire _17525_;
 wire _17526_;
 wire _17527_;
 wire _17528_;
 wire _17529_;
 wire _17530_;
 wire _17531_;
 wire _17532_;
 wire _17533_;
 wire _17534_;
 wire _17535_;
 wire _17536_;
 wire _17537_;
 wire _17538_;
 wire _17539_;
 wire _17540_;
 wire _17541_;
 wire _17542_;
 wire _17543_;
 wire _17544_;
 wire _17545_;
 wire _17546_;
 wire _17547_;
 wire _17548_;
 wire _17549_;
 wire _17550_;
 wire _17551_;
 wire _17552_;
 wire _17553_;
 wire _17554_;
 wire _17555_;
 wire _17556_;
 wire _17557_;
 wire _17558_;
 wire _17559_;
 wire _17560_;
 wire _17561_;
 wire _17562_;
 wire _17563_;
 wire _17564_;
 wire _17565_;
 wire _17566_;
 wire _17567_;
 wire _17568_;
 wire _17569_;
 wire _17570_;
 wire _17571_;
 wire _17572_;
 wire _17573_;
 wire _17574_;
 wire _17575_;
 wire _17576_;
 wire _17577_;
 wire _17578_;
 wire _17579_;
 wire _17580_;
 wire _17581_;
 wire _17582_;
 wire _17583_;
 wire _17584_;
 wire _17585_;
 wire _17586_;
 wire _17587_;
 wire _17588_;
 wire _17589_;
 wire _17590_;
 wire _17591_;
 wire _17592_;
 wire _17593_;
 wire _17594_;
 wire _17595_;
 wire _17596_;
 wire _17597_;
 wire _17598_;
 wire _17599_;
 wire _17600_;
 wire _17601_;
 wire _17602_;
 wire _17603_;
 wire _17604_;
 wire _17605_;
 wire _17606_;
 wire _17607_;
 wire _17608_;
 wire _17609_;
 wire _17610_;
 wire _17611_;
 wire _17612_;
 wire _17613_;
 wire _17614_;
 wire _17615_;
 wire _17616_;
 wire _17617_;
 wire _17618_;
 wire _17619_;
 wire _17620_;
 wire _17621_;
 wire _17622_;
 wire _17623_;
 wire _17624_;
 wire _17625_;
 wire _17626_;
 wire _17627_;
 wire _17628_;
 wire _17629_;
 wire _17630_;
 wire _17631_;
 wire _17632_;
 wire _17633_;
 wire _17634_;
 wire _17635_;
 wire _17636_;
 wire _17637_;
 wire _17638_;
 wire _17639_;
 wire _17640_;
 wire _17641_;
 wire _17642_;
 wire _17643_;
 wire _17644_;
 wire _17645_;
 wire _17646_;
 wire _17647_;
 wire _17648_;
 wire _17649_;
 wire _17650_;
 wire _17651_;
 wire _17652_;
 wire _17653_;
 wire _17654_;
 wire _17655_;
 wire _17656_;
 wire _17657_;
 wire _17658_;
 wire _17659_;
 wire _17660_;
 wire _17661_;
 wire _17662_;
 wire _17663_;
 wire _17664_;
 wire _17665_;
 wire _17666_;
 wire _17667_;
 wire _17668_;
 wire _17669_;
 wire _17670_;
 wire _17671_;
 wire _17672_;
 wire _17673_;
 wire _17674_;
 wire _17675_;
 wire _17676_;
 wire _17677_;
 wire _17678_;
 wire _17679_;
 wire _17680_;
 wire _17681_;
 wire _17682_;
 wire _17683_;
 wire _17684_;
 wire _17685_;
 wire _17686_;
 wire _17687_;
 wire _17688_;
 wire _17689_;
 wire _17690_;
 wire _17691_;
 wire _17692_;
 wire _17693_;
 wire _17694_;
 wire _17695_;
 wire _17696_;
 wire _17697_;
 wire _17698_;
 wire _17699_;
 wire _17700_;
 wire _17701_;
 wire _17702_;
 wire _17703_;
 wire _17704_;
 wire _17705_;
 wire _17706_;
 wire _17707_;
 wire _17708_;
 wire _17709_;
 wire _17710_;
 wire _17711_;
 wire _17712_;
 wire _17713_;
 wire _17714_;
 wire _17715_;
 wire _17716_;
 wire _17717_;
 wire _17718_;
 wire _17719_;
 wire _17720_;
 wire _17721_;
 wire _17722_;
 wire _17723_;
 wire _17724_;
 wire _17725_;
 wire _17726_;
 wire _17727_;
 wire _17728_;
 wire _17729_;
 wire _17730_;
 wire _17731_;
 wire _17732_;
 wire _17733_;
 wire _17734_;
 wire _17735_;
 wire _17736_;
 wire _17737_;
 wire _17738_;
 wire _17739_;
 wire _17740_;
 wire _17741_;
 wire _17742_;
 wire _17743_;
 wire _17744_;
 wire _17745_;
 wire _17746_;
 wire _17747_;
 wire _17748_;
 wire _17749_;
 wire _17750_;
 wire _17751_;
 wire _17752_;
 wire _17753_;
 wire _17754_;
 wire _17755_;
 wire _17756_;
 wire _17757_;
 wire _17758_;
 wire _17759_;
 wire _17760_;
 wire _17761_;
 wire _17762_;
 wire _17763_;
 wire _17764_;
 wire _17765_;
 wire _17766_;
 wire _17767_;
 wire _17768_;
 wire _17769_;
 wire _17770_;
 wire _17771_;
 wire _17772_;
 wire _17773_;
 wire _17774_;
 wire _17775_;
 wire _17776_;
 wire _17777_;
 wire _17778_;
 wire _17779_;
 wire _17780_;
 wire _17781_;
 wire _17782_;
 wire _17783_;
 wire _17784_;
 wire _17785_;
 wire _17786_;
 wire _17787_;
 wire _17788_;
 wire _17789_;
 wire _17790_;
 wire _17791_;
 wire _17792_;
 wire _17793_;
 wire _17794_;
 wire _17795_;
 wire _17796_;
 wire _17797_;
 wire _17798_;
 wire _17799_;
 wire _17800_;
 wire _17801_;
 wire _17802_;
 wire _17803_;
 wire _17804_;
 wire _17805_;
 wire _17806_;
 wire _17807_;
 wire _17808_;
 wire _17809_;
 wire _17810_;
 wire _17811_;
 wire _17812_;
 wire net848;
 wire net1312;
 wire _17815_;
 wire _17816_;
 wire _17817_;
 wire _17818_;
 wire _17819_;
 wire _17820_;
 wire _17821_;
 wire _17822_;
 wire _17823_;
 wire _17824_;
 wire _17825_;
 wire _17826_;
 wire _17827_;
 wire _17828_;
 wire _17829_;
 wire _17830_;
 wire _17831_;
 wire _17832_;
 wire _17833_;
 wire _17834_;
 wire _17835_;
 wire _17836_;
 wire _17837_;
 wire _17838_;
 wire _17839_;
 wire _17840_;
 wire _17841_;
 wire _17842_;
 wire _17843_;
 wire _17844_;
 wire _17845_;
 wire _17846_;
 wire _17847_;
 wire _17848_;
 wire _17849_;
 wire _17850_;
 wire _17851_;
 wire _17852_;
 wire _17853_;
 wire _17854_;
 wire _17855_;
 wire _17856_;
 wire _17857_;
 wire _17858_;
 wire _17859_;
 wire _17860_;
 wire _17861_;
 wire _17862_;
 wire _17863_;
 wire _17864_;
 wire _17865_;
 wire _17866_;
 wire _17867_;
 wire _17868_;
 wire _17869_;
 wire _17870_;
 wire _17871_;
 wire _17872_;
 wire _17873_;
 wire _17874_;
 wire _17875_;
 wire _17876_;
 wire _17877_;
 wire _17878_;
 wire _17879_;
 wire _17880_;
 wire _17881_;
 wire _17882_;
 wire _17883_;
 wire _17884_;
 wire _17885_;
 wire _17886_;
 wire _17887_;
 wire _17888_;
 wire _17889_;
 wire _17890_;
 wire _17891_;
 wire _17892_;
 wire _17893_;
 wire _17894_;
 wire _17895_;
 wire _17896_;
 wire _17897_;
 wire _17898_;
 wire _17899_;
 wire _17900_;
 wire _17901_;
 wire _17902_;
 wire _17903_;
 wire _17904_;
 wire _17905_;
 wire _17906_;
 wire _17907_;
 wire _17908_;
 wire _17909_;
 wire _17910_;
 wire _17911_;
 wire _17912_;
 wire _17913_;
 wire _17914_;
 wire _17915_;
 wire _17916_;
 wire _17917_;
 wire _17918_;
 wire _17919_;
 wire _17920_;
 wire _17921_;
 wire _17922_;
 wire _17923_;
 wire _17924_;
 wire _17925_;
 wire _17926_;
 wire _17927_;
 wire _17928_;
 wire _17929_;
 wire _17930_;
 wire _17931_;
 wire _17932_;
 wire _17933_;
 wire _17934_;
 wire _17935_;
 wire _17936_;
 wire _17937_;
 wire _17938_;
 wire _17939_;
 wire _17940_;
 wire _17941_;
 wire _17942_;
 wire _17943_;
 wire _17944_;
 wire _17945_;
 wire _17946_;
 wire _17947_;
 wire _17948_;
 wire _17949_;
 wire _17950_;
 wire _17951_;
 wire _17952_;
 wire _17953_;
 wire _17954_;
 wire _17955_;
 wire _17956_;
 wire _17957_;
 wire _17958_;
 wire _17959_;
 wire _17960_;
 wire _17961_;
 wire _17962_;
 wire _17963_;
 wire _17964_;
 wire _17965_;
 wire _17966_;
 wire _17967_;
 wire _17968_;
 wire _17969_;
 wire _17970_;
 wire _17971_;
 wire _17972_;
 wire _17973_;
 wire _17974_;
 wire _17975_;
 wire _17976_;
 wire _17977_;
 wire _17978_;
 wire _17979_;
 wire _17980_;
 wire _17981_;
 wire _17982_;
 wire _17983_;
 wire _17984_;
 wire _17985_;
 wire _17986_;
 wire _17987_;
 wire _17988_;
 wire _17989_;
 wire _17990_;
 wire _17991_;
 wire _17992_;
 wire _17993_;
 wire _17994_;
 wire _17995_;
 wire _17996_;
 wire _17997_;
 wire _17998_;
 wire _17999_;
 wire _18000_;
 wire _18001_;
 wire _18002_;
 wire _18003_;
 wire _18004_;
 wire _18005_;
 wire _18006_;
 wire _18007_;
 wire _18008_;
 wire _18009_;
 wire _18010_;
 wire _18011_;
 wire _18012_;
 wire _18013_;
 wire _18014_;
 wire _18015_;
 wire _18016_;
 wire _18017_;
 wire _18018_;
 wire _18019_;
 wire _18020_;
 wire _18021_;
 wire _18022_;
 wire _18023_;
 wire _18024_;
 wire _18025_;
 wire _18026_;
 wire _18027_;
 wire _18028_;
 wire _18029_;
 wire _18030_;
 wire _18031_;
 wire _18032_;
 wire _18033_;
 wire _18034_;
 wire _18035_;
 wire _18036_;
 wire _18037_;
 wire _18038_;
 wire _18039_;
 wire _18040_;
 wire _18041_;
 wire _18042_;
 wire _18043_;
 wire _18044_;
 wire _18045_;
 wire _18046_;
 wire _18047_;
 wire _18048_;
 wire _18049_;
 wire _18050_;
 wire _18051_;
 wire _18052_;
 wire _18053_;
 wire _18054_;
 wire _18055_;
 wire _18056_;
 wire _18057_;
 wire _18058_;
 wire _18059_;
 wire _18060_;
 wire _18061_;
 wire _18062_;
 wire _18063_;
 wire _18064_;
 wire _18065_;
 wire _18066_;
 wire _18067_;
 wire _18068_;
 wire _18069_;
 wire _18070_;
 wire _18071_;
 wire _18072_;
 wire _18073_;
 wire _18074_;
 wire _18075_;
 wire _18076_;
 wire _18077_;
 wire _18078_;
 wire _18079_;
 wire _18080_;
 wire _18081_;
 wire _18082_;
 wire _18083_;
 wire _18084_;
 wire _18085_;
 wire _18086_;
 wire _18087_;
 wire _18088_;
 wire _18089_;
 wire _18090_;
 wire _18091_;
 wire _18092_;
 wire _18093_;
 wire _18094_;
 wire _18095_;
 wire _18096_;
 wire _18097_;
 wire _18098_;
 wire _18099_;
 wire _18100_;
 wire _18101_;
 wire _18102_;
 wire _18103_;
 wire _18104_;
 wire _18105_;
 wire _18106_;
 wire _18107_;
 wire _18108_;
 wire _18109_;
 wire _18110_;
 wire _18111_;
 wire _18112_;
 wire _18113_;
 wire _18114_;
 wire _18115_;
 wire _18116_;
 wire _18117_;
 wire _18118_;
 wire _18119_;
 wire _18120_;
 wire _18121_;
 wire _18122_;
 wire _18123_;
 wire _18124_;
 wire _18125_;
 wire _18126_;
 wire _18127_;
 wire _18128_;
 wire _18129_;
 wire _18130_;
 wire _18131_;
 wire _18132_;
 wire _18133_;
 wire _18134_;
 wire _18135_;
 wire _18136_;
 wire _18137_;
 wire _18138_;
 wire _18139_;
 wire _18140_;
 wire _18141_;
 wire _18142_;
 wire _18143_;
 wire _18144_;
 wire _18145_;
 wire _18146_;
 wire _18147_;
 wire _18148_;
 wire _18149_;
 wire _18150_;
 wire _18151_;
 wire _18152_;
 wire _18153_;
 wire _18154_;
 wire _18155_;
 wire _18156_;
 wire _18157_;
 wire _18158_;
 wire _18159_;
 wire _18160_;
 wire _18161_;
 wire _18162_;
 wire _18163_;
 wire _18164_;
 wire _18165_;
 wire _18166_;
 wire _18167_;
 wire _18168_;
 wire _18169_;
 wire _18170_;
 wire _18171_;
 wire _18172_;
 wire _18173_;
 wire _18174_;
 wire _18175_;
 wire _18176_;
 wire _18177_;
 wire _18178_;
 wire _18179_;
 wire _18180_;
 wire _18181_;
 wire _18182_;
 wire _18183_;
 wire _18184_;
 wire _18185_;
 wire _18186_;
 wire _18187_;
 wire _18188_;
 wire _18189_;
 wire _18190_;
 wire _18191_;
 wire _18192_;
 wire _18193_;
 wire _18194_;
 wire _18195_;
 wire _18196_;
 wire _18197_;
 wire _18198_;
 wire _18199_;
 wire _18200_;
 wire _18201_;
 wire _18202_;
 wire _18203_;
 wire _18204_;
 wire _18205_;
 wire _18206_;
 wire _18207_;
 wire _18208_;
 wire _18209_;
 wire _18210_;
 wire _18211_;
 wire _18212_;
 wire _18213_;
 wire _18214_;
 wire _18215_;
 wire _18216_;
 wire _18217_;
 wire _18218_;
 wire _18219_;
 wire _18220_;
 wire _18221_;
 wire _18222_;
 wire _18223_;
 wire _18224_;
 wire _18225_;
 wire _18226_;
 wire _18227_;
 wire _18228_;
 wire _18229_;
 wire _18230_;
 wire _18231_;
 wire _18232_;
 wire _18233_;
 wire _18234_;
 wire _18235_;
 wire _18236_;
 wire _18237_;
 wire _18238_;
 wire _18239_;
 wire _18240_;
 wire _18241_;
 wire _18242_;
 wire _18243_;
 wire _18244_;
 wire _18245_;
 wire _18246_;
 wire _18247_;
 wire _18248_;
 wire _18249_;
 wire _18250_;
 wire _18251_;
 wire _18252_;
 wire _18253_;
 wire _18254_;
 wire _18255_;
 wire _18256_;
 wire _18257_;
 wire _18258_;
 wire _18259_;
 wire _18260_;
 wire _18261_;
 wire _18262_;
 wire _18263_;
 wire _18264_;
 wire _18265_;
 wire _18266_;
 wire _18267_;
 wire _18268_;
 wire _18269_;
 wire _18270_;
 wire _18271_;
 wire _18272_;
 wire _18273_;
 wire _18274_;
 wire _18275_;
 wire _18276_;
 wire _18277_;
 wire _18278_;
 wire _18279_;
 wire _18280_;
 wire _18281_;
 wire _18282_;
 wire _18283_;
 wire _18284_;
 wire _18285_;
 wire _18286_;
 wire _18287_;
 wire _18288_;
 wire _18289_;
 wire _18290_;
 wire _18291_;
 wire _18292_;
 wire _18293_;
 wire _18294_;
 wire _18295_;
 wire _18296_;
 wire _18297_;
 wire _18298_;
 wire _18299_;
 wire _18300_;
 wire _18301_;
 wire _18302_;
 wire _18303_;
 wire _18304_;
 wire _18305_;
 wire _18306_;
 wire _18307_;
 wire _18308_;
 wire _18309_;
 wire _18310_;
 wire _18311_;
 wire _18312_;
 wire _18313_;
 wire _18314_;
 wire _18315_;
 wire _18316_;
 wire _18317_;
 wire _18318_;
 wire _18319_;
 wire _18320_;
 wire _18321_;
 wire net1446;
 wire net1587;
 wire _18324_;
 wire net1352;
 wire _18326_;
 wire net1450;
 wire net1405;
 wire _18329_;
 wire _18330_;
 wire net1588;
 wire _18332_;
 wire _18333_;
 wire net1045;
 wire _18335_;
 wire _18336_;
 wire _18337_;
 wire net1346;
 wire _18339_;
 wire net1347;
 wire _18341_;
 wire _18342_;
 wire net1340;
 wire _18344_;
 wire net1342;
 wire _18346_;
 wire _18347_;
 wire net1041;
 wire net1248;
 wire net1334;
 wire _18351_;
 wire _18352_;
 wire _18353_;
 wire net1246;
 wire _18355_;
 wire _18356_;
 wire _18357_;
 wire net1327;
 wire net1242;
 wire _18360_;
 wire _18361_;
 wire _18362_;
 wire _18363_;
 wire net1240;
 wire _18365_;
 wire _18366_;
 wire _18367_;
 wire net1318;
 wire net1239;
 wire _18370_;
 wire _18371_;
 wire _18372_;
 wire net1314;
 wire net1236;
 wire _18375_;
 wire _18376_;
 wire _18377_;
 wire net1313;
 wire _18379_;
 wire _18380_;
 wire _18381_;
 wire _18382_;
 wire _18383_;
 wire _18384_;
 wire _18385_;
 wire _18386_;
 wire _18387_;
 wire _18388_;
 wire _18389_;
 wire _18390_;
 wire _18391_;
 wire _18392_;
 wire _18393_;
 wire _18394_;
 wire _18395_;
 wire _18396_;
 wire _18397_;
 wire net1145;
 wire _18399_;
 wire _18400_;
 wire net1146;
 wire _18402_;
 wire _18403_;
 wire _18404_;
 wire _18405_;
 wire net1121;
 wire _18407_;
 wire _18408_;
 wire _18409_;
 wire _18410_;
 wire net1111;
 wire _18412_;
 wire _18413_;
 wire net1101;
 wire _18415_;
 wire _18416_;
 wire _18417_;
 wire _18418_;
 wire _18419_;
 wire net1093;
 wire _18421_;
 wire _18422_;
 wire _18423_;
 wire _18424_;
 wire _18425_;
 wire _18426_;
 wire _18427_;
 wire net1086;
 wire _18429_;
 wire _18430_;
 wire net1085;
 wire _18432_;
 wire net1084;
 wire _18434_;
 wire _18435_;
 wire _18436_;
 wire _18437_;
 wire net1082;
 wire _18439_;
 wire _18440_;
 wire _18441_;
 wire _18442_;
 wire net1080;
 wire _18444_;
 wire _18445_;
 wire _18446_;
 wire _18447_;
 wire net1079;
 wire _18449_;
 wire _18450_;
 wire net1078;
 wire _18452_;
 wire net1075;
 wire net1076;
 wire _18455_;
 wire _18456_;
 wire _18457_;
 wire net1072;
 wire _18459_;
 wire _18460_;
 wire net1073;
 wire _18462_;
 wire net1071;
 wire net1070;
 wire _18465_;
 wire _18466_;
 wire _18467_;
 wire net1069;
 wire _18469_;
 wire _18470_;
 wire _18471_;
 wire _18472_;
 wire net1068;
 wire _18474_;
 wire _18475_;
 wire _18476_;
 wire _18477_;
 wire _18478_;
 wire _18479_;
 wire _18480_;
 wire _18481_;
 wire _18482_;
 wire _18483_;
 wire _18484_;
 wire _18485_;
 wire _18486_;
 wire _18487_;
 wire _18488_;
 wire _18489_;
 wire _18490_;
 wire _18491_;
 wire _18492_;
 wire _18493_;
 wire _18494_;
 wire _18495_;
 wire _18496_;
 wire _18497_;
 wire _18498_;
 wire _18499_;
 wire _18500_;
 wire _18501_;
 wire _18502_;
 wire _18503_;
 wire _18504_;
 wire _18505_;
 wire _18506_;
 wire _18507_;
 wire _18508_;
 wire _18509_;
 wire _18510_;
 wire _18511_;
 wire _18512_;
 wire _18513_;
 wire _18514_;
 wire _18515_;
 wire _18516_;
 wire _18517_;
 wire _18518_;
 wire _18519_;
 wire _18520_;
 wire _18521_;
 wire _18522_;
 wire _18523_;
 wire _18524_;
 wire _18525_;
 wire _18526_;
 wire _18527_;
 wire _18528_;
 wire _18529_;
 wire _18530_;
 wire _18531_;
 wire _18532_;
 wire _18533_;
 wire _18534_;
 wire _18535_;
 wire _18536_;
 wire _18537_;
 wire _18538_;
 wire _18539_;
 wire _18540_;
 wire _18541_;
 wire _18542_;
 wire _18543_;
 wire _18544_;
 wire _18545_;
 wire _18546_;
 wire _18547_;
 wire _18548_;
 wire _18549_;
 wire _18550_;
 wire _18551_;
 wire _18552_;
 wire _18553_;
 wire _18554_;
 wire _18555_;
 wire _18556_;
 wire _18557_;
 wire _18558_;
 wire _18559_;
 wire _18560_;
 wire _18561_;
 wire _18562_;
 wire _18563_;
 wire _18564_;
 wire _18565_;
 wire _18566_;
 wire _18567_;
 wire _18568_;
 wire _18569_;
 wire _18570_;
 wire _18571_;
 wire _18572_;
 wire _18573_;
 wire _18574_;
 wire _18575_;
 wire _18576_;
 wire _18577_;
 wire _18578_;
 wire _18579_;
 wire _18580_;
 wire _18581_;
 wire _18582_;
 wire _18583_;
 wire _18584_;
 wire _18585_;
 wire _18586_;
 wire _18587_;
 wire _18588_;
 wire _18589_;
 wire _18590_;
 wire _18591_;
 wire _18592_;
 wire _18593_;
 wire _18594_;
 wire _18595_;
 wire _18596_;
 wire _18597_;
 wire _18598_;
 wire _18599_;
 wire _18600_;
 wire _18601_;
 wire _18602_;
 wire _18603_;
 wire _18604_;
 wire _18605_;
 wire clknet_leaf_0_clk_i;
 wire net29;
 wire net467;
 wire core_busy_d;
 wire \core_clock_gate_i.clk_o ;
 wire \core_clock_gate_i.en_latch ;
 wire \cs_registers_i.mcycle_counter_i.counter[0] ;
 wire \cs_registers_i.mcycle_counter_i.counter[10] ;
 wire \cs_registers_i.mcycle_counter_i.counter[12] ;
 wire \cs_registers_i.mcycle_counter_i.counter[14] ;
 wire \cs_registers_i.mcycle_counter_i.counter[16] ;
 wire \cs_registers_i.mcycle_counter_i.counter[18] ;
 wire \cs_registers_i.mcycle_counter_i.counter[1] ;
 wire \cs_registers_i.mcycle_counter_i.counter[20] ;
 wire \cs_registers_i.mcycle_counter_i.counter[22] ;
 wire \cs_registers_i.mcycle_counter_i.counter[24] ;
 wire \cs_registers_i.mcycle_counter_i.counter[26] ;
 wire \cs_registers_i.mcycle_counter_i.counter[28] ;
 wire \cs_registers_i.mcycle_counter_i.counter[2] ;
 wire \cs_registers_i.mcycle_counter_i.counter[30] ;
 wire \cs_registers_i.mcycle_counter_i.counter[32] ;
 wire \cs_registers_i.mcycle_counter_i.counter[34] ;
 wire \cs_registers_i.mcycle_counter_i.counter[36] ;
 wire \cs_registers_i.mcycle_counter_i.counter[38] ;
 wire \cs_registers_i.mcycle_counter_i.counter[40] ;
 wire \cs_registers_i.mcycle_counter_i.counter[42] ;
 wire \cs_registers_i.mcycle_counter_i.counter[44] ;
 wire \cs_registers_i.mcycle_counter_i.counter[46] ;
 wire \cs_registers_i.mcycle_counter_i.counter[48] ;
 wire \cs_registers_i.mcycle_counter_i.counter[4] ;
 wire \cs_registers_i.mcycle_counter_i.counter[50] ;
 wire \cs_registers_i.mcycle_counter_i.counter[52] ;
 wire \cs_registers_i.mcycle_counter_i.counter[54] ;
 wire \cs_registers_i.mcycle_counter_i.counter[56] ;
 wire \cs_registers_i.mcycle_counter_i.counter[58] ;
 wire \cs_registers_i.mcycle_counter_i.counter[60] ;
 wire \cs_registers_i.mcycle_counter_i.counter[62] ;
 wire \cs_registers_i.mcycle_counter_i.counter[6] ;
 wire \cs_registers_i.mcycle_counter_i.counter[8] ;
 wire \cs_registers_i.mhpmcounter[2][0] ;
 wire \cs_registers_i.mhpmcounter[2][10] ;
 wire \cs_registers_i.mhpmcounter[2][12] ;
 wire \cs_registers_i.mhpmcounter[2][14] ;
 wire \cs_registers_i.mhpmcounter[2][16] ;
 wire \cs_registers_i.mhpmcounter[2][18] ;
 wire \cs_registers_i.mhpmcounter[2][1] ;
 wire \cs_registers_i.mhpmcounter[2][20] ;
 wire \cs_registers_i.mhpmcounter[2][22] ;
 wire \cs_registers_i.mhpmcounter[2][24] ;
 wire \cs_registers_i.mhpmcounter[2][26] ;
 wire \cs_registers_i.mhpmcounter[2][28] ;
 wire \cs_registers_i.mhpmcounter[2][2] ;
 wire \cs_registers_i.mhpmcounter[2][30] ;
 wire \cs_registers_i.mhpmcounter[2][32] ;
 wire \cs_registers_i.mhpmcounter[2][34] ;
 wire \cs_registers_i.mhpmcounter[2][36] ;
 wire \cs_registers_i.mhpmcounter[2][38] ;
 wire \cs_registers_i.mhpmcounter[2][40] ;
 wire \cs_registers_i.mhpmcounter[2][42] ;
 wire \cs_registers_i.mhpmcounter[2][44] ;
 wire \cs_registers_i.mhpmcounter[2][46] ;
 wire \cs_registers_i.mhpmcounter[2][48] ;
 wire \cs_registers_i.mhpmcounter[2][4] ;
 wire \cs_registers_i.mhpmcounter[2][50] ;
 wire \cs_registers_i.mhpmcounter[2][52] ;
 wire \cs_registers_i.mhpmcounter[2][54] ;
 wire \cs_registers_i.mhpmcounter[2][56] ;
 wire \cs_registers_i.mhpmcounter[2][58] ;
 wire \cs_registers_i.mhpmcounter[2][60] ;
 wire \cs_registers_i.mhpmcounter[2][62] ;
 wire \cs_registers_i.mhpmcounter[2][6] ;
 wire \cs_registers_i.mhpmcounter[2][8] ;
 wire \cs_registers_i.pc_id_i[11] ;
 wire \cs_registers_i.pc_id_i[13] ;
 wire \cs_registers_i.pc_id_i[15] ;
 wire \cs_registers_i.pc_id_i[17] ;
 wire \cs_registers_i.pc_id_i[19] ;
 wire \cs_registers_i.pc_id_i[1] ;
 wire \cs_registers_i.pc_id_i[21] ;
 wire \cs_registers_i.pc_id_i[23] ;
 wire \cs_registers_i.pc_id_i[25] ;
 wire \cs_registers_i.pc_id_i[27] ;
 wire \cs_registers_i.pc_id_i[29] ;
 wire \cs_registers_i.pc_id_i[2] ;
 wire \cs_registers_i.pc_id_i[3] ;
 wire \cs_registers_i.pc_id_i[5] ;
 wire \cs_registers_i.pc_id_i[7] ;
 wire \cs_registers_i.pc_id_i[9] ;
 wire \cs_registers_i.pc_if_i[11] ;
 wire \cs_registers_i.pc_if_i[13] ;
 wire \cs_registers_i.pc_if_i[15] ;
 wire \cs_registers_i.pc_if_i[17] ;
 wire \cs_registers_i.pc_if_i[19] ;
 wire \cs_registers_i.pc_if_i[21] ;
 wire \cs_registers_i.pc_if_i[23] ;
 wire \cs_registers_i.pc_if_i[25] ;
 wire \cs_registers_i.pc_if_i[27] ;
 wire \cs_registers_i.pc_if_i[29] ;
 wire \cs_registers_i.pc_if_i[2] ;
 wire \cs_registers_i.pc_if_i[3] ;
 wire \cs_registers_i.pc_if_i[5] ;
 wire \cs_registers_i.pc_if_i[7] ;
 wire \cs_registers_i.pc_if_i[9] ;
 wire \cs_registers_i.priv_lvl_q[0] ;
 wire \ex_block_i.alu_adder_result_ex_o[0] ;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire \ex_block_i.alu_adder_result_ex_o[1] ;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \id_stage_i.branch_set_d ;
 wire \id_stage_i.controller_i.exc_req_d ;
 wire \id_stage_i.controller_i.illegal_insn_d ;
 wire \id_stage_i.controller_i.load_err_d ;
 wire \id_stage_i.controller_i.store_err_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \if_stage_i.instr_valid_id_d ;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_0_clk_i;
 wire clknet_2_0__leaf_clk_i;
 wire clknet_2_1__leaf_clk_i;
 wire clknet_2_2__leaf_clk_i;
 wire clknet_2_3__leaf_clk_i;
 wire clknet_level_0_1_10_clk_i;
 wire clknet_level_1_1_11_clk_i;
 wire clknet_level_2_1_12_clk_i;
 wire clknet_level_3_1_13_clk_i;
 wire clknet_level_0_1_24_clk_i;
 wire clknet_level_1_1_25_clk_i;
 wire clknet_level_2_1_26_clk_i;
 wire clknet_level_3_1_27_clk_i;
 wire clknet_level_0_1_38_clk_i;
 wire clknet_level_1_1_39_clk_i;
 wire clknet_level_2_1_310_clk_i;
 wire clknet_level_3_1_311_clk_i;
 wire clknet_level_0_1_412_clk_i;
 wire clknet_level_1_1_413_clk_i;
 wire clknet_level_2_1_414_clk_i;
 wire clknet_level_3_1_415_clk_i;
 wire clknet_level_0_1_516_clk_i;
 wire clknet_level_1_1_517_clk_i;
 wire clknet_level_2_1_518_clk_i;
 wire clknet_level_3_1_519_clk_i;
 wire clknet_level_0_1_620_clk_i;
 wire clknet_level_1_1_621_clk_i;
 wire clknet_level_2_1_622_clk_i;
 wire clknet_level_3_1_623_clk_i;
 wire clknet_level_0_1_724_clk_i;
 wire clknet_level_1_1_725_clk_i;
 wire clknet_level_2_1_726_clk_i;
 wire clknet_level_3_1_727_clk_i;
 wire clknet_level_0_1_828_clk_i;
 wire clknet_level_1_1_829_clk_i;
 wire clknet_level_2_1_830_clk_i;
 wire clknet_level_3_1_831_clk_i;
 wire clknet_level_0_1_932_clk_i;
 wire clknet_level_1_1_933_clk_i;
 wire clknet_level_2_1_934_clk_i;
 wire clknet_level_3_1_935_clk_i;
 wire clknet_level_0_1_1036_clk_i;
 wire clknet_level_1_1_1037_clk_i;
 wire clknet_level_2_1_1038_clk_i;
 wire clknet_level_3_1_1039_clk_i;
 wire clknet_level_0_1_1140_clk_i;
 wire clknet_level_1_1_1141_clk_i;
 wire clknet_level_2_1_1142_clk_i;
 wire clknet_level_3_1_1143_clk_i;
 wire clknet_level_0_1_1244_clk_i;
 wire clknet_level_1_1_1245_clk_i;
 wire clknet_level_2_1_1246_clk_i;
 wire clknet_level_3_1_1247_clk_i;
 wire clknet_level_0_1_1348_clk_i;
 wire clknet_level_1_1_1349_clk_i;
 wire clknet_level_2_1_1350_clk_i;
 wire clknet_level_3_1_1351_clk_i;
 wire clknet_level_0_1_1452_clk_i;
 wire clknet_level_1_1_1453_clk_i;
 wire clknet_level_2_1_1454_clk_i;
 wire clknet_level_3_1_1455_clk_i;
 wire clknet_level_0_1_1556_clk_i;
 wire clknet_level_1_1_1557_clk_i;
 wire clknet_level_2_1_1558_clk_i;
 wire clknet_level_3_1_1559_clk_i;
 wire clknet_level_0_1_1660_clk_i;
 wire clknet_level_1_1_1661_clk_i;
 wire clknet_level_2_1_1662_clk_i;
 wire clknet_level_3_1_1663_clk_i;
 wire clknet_level_0_1_1764_clk_i;
 wire clknet_level_1_1_1765_clk_i;
 wire clknet_level_2_1_1766_clk_i;
 wire clknet_level_3_1_1767_clk_i;
 wire clknet_level_0_1_1868_clk_i;
 wire clknet_level_1_1_1869_clk_i;
 wire clknet_level_2_1_1870_clk_i;
 wire clknet_level_3_1_1871_clk_i;
 wire clknet_level_0_1_1972_clk_i;
 wire clknet_level_1_1_1973_clk_i;
 wire clknet_level_2_1_1974_clk_i;
 wire clknet_level_3_1_1975_clk_i;
 wire clknet_level_0_1_2076_clk_i;
 wire clknet_level_1_1_2077_clk_i;
 wire clknet_level_2_1_2078_clk_i;
 wire clknet_level_3_1_2079_clk_i;
 wire clknet_level_0_1_2180_clk_i;
 wire clknet_level_1_1_2181_clk_i;
 wire clknet_level_2_1_2182_clk_i;
 wire clknet_level_3_1_2183_clk_i;
 wire clknet_level_0_1_2284_clk_i;
 wire clknet_level_1_1_2285_clk_i;
 wire clknet_level_2_1_2286_clk_i;
 wire clknet_level_3_1_2287_clk_i;
 wire clknet_level_0_1_2388_clk_i;
 wire clknet_level_1_1_2389_clk_i;
 wire clknet_level_2_1_2390_clk_i;
 wire clknet_level_3_1_2391_clk_i;
 wire clknet_level_0_1_2492_clk_i;
 wire clknet_level_1_1_2493_clk_i;
 wire clknet_level_2_1_2494_clk_i;
 wire clknet_level_3_1_2495_clk_i;
 wire clknet_level_0_1_2596_clk_i;
 wire clknet_level_1_1_2597_clk_i;
 wire clknet_level_2_1_2598_clk_i;
 wire clknet_level_3_1_2599_clk_i;
 wire clknet_level_0_1_26100_clk_i;
 wire clknet_level_1_1_26101_clk_i;
 wire clknet_level_2_1_26102_clk_i;
 wire clknet_level_3_1_26103_clk_i;
 wire clknet_level_0_1_27104_clk_i;
 wire clknet_level_1_1_27105_clk_i;
 wire clknet_level_2_1_27106_clk_i;
 wire clknet_level_3_1_27107_clk_i;
 wire clknet_level_0_1_28108_clk_i;
 wire clknet_level_1_1_28109_clk_i;
 wire clknet_level_2_1_28110_clk_i;
 wire clknet_level_3_1_28111_clk_i;
 wire clknet_level_0_1_29112_clk_i;
 wire clknet_level_1_1_29113_clk_i;
 wire clknet_level_2_1_29114_clk_i;
 wire clknet_level_3_1_29115_clk_i;
 wire clknet_level_0_1_30116_clk_i;
 wire clknet_level_1_1_30117_clk_i;
 wire clknet_level_2_1_30118_clk_i;
 wire clknet_level_3_1_30119_clk_i;
 wire clknet_level_0_1_31120_clk_i;
 wire clknet_level_1_1_31121_clk_i;
 wire clknet_level_2_1_31122_clk_i;
 wire clknet_level_3_1_31123_clk_i;
 wire clknet_level_0_1_32124_clk_i;
 wire clknet_level_1_1_32125_clk_i;
 wire clknet_level_2_1_32126_clk_i;
 wire clknet_level_3_1_32127_clk_i;
 wire clknet_level_0_1_33128_clk_i;
 wire clknet_level_1_1_33129_clk_i;
 wire clknet_level_2_1_33130_clk_i;
 wire clknet_level_3_1_33131_clk_i;
 wire clknet_level_0_1_34132_clk_i;
 wire clknet_level_1_1_34133_clk_i;
 wire clknet_level_2_1_34134_clk_i;
 wire clknet_level_3_1_34135_clk_i;
 wire \clknet_leaf_0_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_1_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_2_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_3_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_4_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_5_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_6_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_7_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_8_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_9_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_10_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_11_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_12_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_13_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_14_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_15_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_16_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_17_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_18_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_19_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_20_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_21_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_22_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_23_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_24_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_25_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_26_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_27_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_28_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_29_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_30_core_clock_gate_i.clk_o ;
 wire \clknet_leaf_31_core_clock_gate_i.clk_o ;
 wire \clknet_0_core_clock_gate_i.clk_o ;
 wire \clknet_2_0__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_1__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_2__leaf_core_clock_gate_i.clk_o ;
 wire \clknet_2_3__leaf_core_clock_gate_i.clk_o ;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;

 TIEHIx1_ASAP7_75t_R _34951__538 (.H(net538));
 TIEHIx1_ASAP7_75t_R _34950__537 (.H(net537));
 TIEHIx1_ASAP7_75t_R _34949__536 (.H(net536));
 TIEHIx1_ASAP7_75t_R _34948__535 (.H(net535));
 TIEHIx1_ASAP7_75t_R _34947__534 (.H(net534));
 INVx1_ASAP7_75t_R _18613_ (.A(_00264_),
    .Y(_13340_));
 TIEHIx1_ASAP7_75t_R _34946__533 (.H(net533));
 NAND2x1_ASAP7_75t_R _18615_ (.A(net346),
    .B(_00262_),
    .Y(_13342_));
 TIEHIx1_ASAP7_75t_R _34945__532 (.H(net532));
 TIEHIx1_ASAP7_75t_R _34944__531 (.H(net531));
 OA211x2_ASAP7_75t_R _18618_ (.A1(net346),
    .A2(_13340_),
    .B(_13342_),
    .C(net336),
    .Y(_13345_));
 TIEHIx1_ASAP7_75t_R _34943__530 (.H(net530));
 TIEHIx1_ASAP7_75t_R _34942__529 (.H(net529));
 INVx1_ASAP7_75t_R _18621_ (.A(_00268_),
    .Y(_13348_));
 NAND2x1_ASAP7_75t_R _18622_ (.A(net2248),
    .B(_00266_),
    .Y(_13349_));
 CKINVDCx20_ASAP7_75t_R _18623_ (.A(net337),
    .Y(_13350_));
 OA211x2_ASAP7_75t_R _18624_ (.A1(net367),
    .A2(_13348_),
    .B(_13349_),
    .C(_13350_),
    .Y(_13351_));
 OR3x1_ASAP7_75t_R _18625_ (.A(net375),
    .B(_13345_),
    .C(_13351_),
    .Y(_13352_));
 TIEHIx1_ASAP7_75t_R _34941__528 (.H(net528));
 TIEHIx1_ASAP7_75t_R _34940__527 (.H(net527));
 CKINVDCx20_ASAP7_75t_R _18628_ (.A(_00244_),
    .Y(_13355_));
 AND2x6_ASAP7_75t_R _18629_ (.A(net332),
    .B(_13355_),
    .Y(_13356_));
 AND2x6_ASAP7_75t_R _18630_ (.A(net376),
    .B(net338),
    .Y(_13357_));
 TIEHIx1_ASAP7_75t_R _34939__526 (.H(net526));
 CKINVDCx20_ASAP7_75t_R _18632_ (.A(net359),
    .Y(_13359_));
 TIEHIx1_ASAP7_75t_R _34938__525 (.H(net525));
 TIEHIx1_ASAP7_75t_R _34937__524 (.H(net524));
 TIEHIx1_ASAP7_75t_R _34936__523 (.H(net523));
 TIEHIx1_ASAP7_75t_R _34935__522 (.H(net522));
 AND2x2_ASAP7_75t_R _18637_ (.A(net346),
    .B(_00261_),
    .Y(_13364_));
 AO21x1_ASAP7_75t_R _18638_ (.A1(net2278),
    .A2(_00263_),
    .B(_13364_),
    .Y(_13365_));
 AND2x6_ASAP7_75t_R _18639_ (.A(net374),
    .B(_13350_),
    .Y(_13366_));
 TIEHIx1_ASAP7_75t_R _34934__521 (.H(net521));
 TIEHIx1_ASAP7_75t_R _34933__520 (.H(net520));
 AND2x2_ASAP7_75t_R _18642_ (.A(net346),
    .B(_00265_),
    .Y(_13369_));
 AO21x1_ASAP7_75t_R _18643_ (.A1(net2278),
    .A2(_00267_),
    .B(_13369_),
    .Y(_13370_));
 AOI22x1_ASAP7_75t_R _18644_ (.A1(_13357_),
    .A2(_13365_),
    .B1(_13366_),
    .B2(_13370_),
    .Y(_13371_));
 AND3x2_ASAP7_75t_R _18645_ (.A(_13352_),
    .B(_13356_),
    .C(_13371_),
    .Y(_13372_));
 CKINVDCx20_ASAP7_75t_R _18646_ (.A(net332),
    .Y(_13373_));
 TIEHIx1_ASAP7_75t_R _34932__519 (.H(net519));
 AND2x2_ASAP7_75t_R _18648_ (.A(_13373_),
    .B(net328),
    .Y(_13375_));
 CKINVDCx20_ASAP7_75t_R _18649_ (.A(net370),
    .Y(_13376_));
 AND2x6_ASAP7_75t_R _18650_ (.A(net323),
    .B(net336),
    .Y(_13377_));
 TIEHIx1_ASAP7_75t_R _34931__518 (.H(net518));
 TIEHIx1_ASAP7_75t_R _34930__517 (.H(net517));
 INVx1_ASAP7_75t_R _18653_ (.A(_00254_),
    .Y(_13380_));
 TIEHIx1_ASAP7_75t_R _34929__516 (.H(net516));
 NOR2x1_ASAP7_75t_R _18655_ (.A(net342),
    .B(_00256_),
    .Y(_13382_));
 AO21x1_ASAP7_75t_R _18656_ (.A1(net342),
    .A2(_13380_),
    .B(_13382_),
    .Y(_13383_));
 TIEHIx1_ASAP7_75t_R _34928__515 (.H(net515));
 INVx1_ASAP7_75t_R _18658_ (.A(_00255_),
    .Y(_13385_));
 TIEHIx1_ASAP7_75t_R _34927__514 (.H(net514));
 NAND2x1_ASAP7_75t_R _18660_ (.A(net342),
    .B(_00253_),
    .Y(_13387_));
 OA211x2_ASAP7_75t_R _18661_ (.A1(net341),
    .A2(_13385_),
    .B(_13357_),
    .C(_13387_),
    .Y(_13388_));
 AO21x1_ASAP7_75t_R _18662_ (.A1(_13377_),
    .A2(_13383_),
    .B(_13388_),
    .Y(_13389_));
 AND2x6_ASAP7_75t_R _18663_ (.A(net370),
    .B(net341),
    .Y(_13390_));
 AND2x6_ASAP7_75t_R _18664_ (.A(net374),
    .B(net326),
    .Y(_13391_));
 TIEHIx1_ASAP7_75t_R _34926__513 (.H(net513));
 TIEHIx1_ASAP7_75t_R _34925__512 (.H(net512));
 OR3x1_ASAP7_75t_R _18667_ (.A(net337),
    .B(_00245_),
    .C(_13355_),
    .Y(_13394_));
 AOI221x1_ASAP7_75t_R _18668_ (.A1(_00257_),
    .A2(_13390_),
    .B1(net2242),
    .B2(_00259_),
    .C(_13394_),
    .Y(_13395_));
 TIEHIx1_ASAP7_75t_R _34924__511 (.H(net511));
 TIEHIx1_ASAP7_75t_R _34923__510 (.H(net510));
 TIEHIx1_ASAP7_75t_R _34922__509 (.H(net509));
 AND2x2_ASAP7_75t_R _18672_ (.A(net341),
    .B(_00258_),
    .Y(_13399_));
 AO21x1_ASAP7_75t_R _18673_ (.A1(net2278),
    .A2(_00260_),
    .B(_13399_),
    .Y(_13400_));
 NAND2x1_ASAP7_75t_R _18674_ (.A(net323),
    .B(_13400_),
    .Y(_13401_));
 NOR2x2_ASAP7_75t_R _18675_ (.A(net374),
    .B(net336),
    .Y(_13402_));
 TIEHIx1_ASAP7_75t_R _34921__508 (.H(net508));
 TIEHIx1_ASAP7_75t_R _34920__507 (.H(net507));
 AND2x2_ASAP7_75t_R _18678_ (.A(net342),
    .B(_00250_),
    .Y(_13405_));
 AO21x1_ASAP7_75t_R _18679_ (.A1(net326),
    .A2(_00252_),
    .B(_13405_),
    .Y(_13406_));
 TIEHIx1_ASAP7_75t_R _34919__506 (.H(net506));
 AND2x2_ASAP7_75t_R _18681_ (.A(net342),
    .B(_00249_),
    .Y(_13408_));
 AO21x1_ASAP7_75t_R _18682_ (.A1(net326),
    .A2(_00251_),
    .B(_13408_),
    .Y(_13409_));
 NAND2x1_ASAP7_75t_R _18683_ (.A(_00245_),
    .B(net328),
    .Y(_13410_));
 AOI221x1_ASAP7_75t_R _18684_ (.A1(_13402_),
    .A2(_13406_),
    .B1(_13409_),
    .B2(_13366_),
    .C(_13410_),
    .Y(_13411_));
 INVx1_ASAP7_75t_R _18685_ (.A(_00247_),
    .Y(_13412_));
 TIEHIx1_ASAP7_75t_R _34918__505 (.H(net505));
 OR2x2_ASAP7_75t_R _18687_ (.A(_00248_),
    .B(net341),
    .Y(_13414_));
 OAI21x1_ASAP7_75t_R _18688_ (.A1(net2278),
    .A2(_01708_),
    .B(_13414_),
    .Y(_13415_));
 TIEHIx1_ASAP7_75t_R _34917__504 (.H(net504));
 TIEHIx1_ASAP7_75t_R _34916__503 (.H(net503));
 AO221x1_ASAP7_75t_R _18691_ (.A1(_13412_),
    .A2(net2244),
    .B1(_13415_),
    .B2(net323),
    .C(_13350_),
    .Y(_13418_));
 AO222x2_ASAP7_75t_R _18692_ (.A1(_13375_),
    .A2(_13389_),
    .B1(_13395_),
    .B2(_13401_),
    .C1(_13411_),
    .C2(_13418_),
    .Y(_13419_));
 TIEHIx1_ASAP7_75t_R _34915__502 (.H(net502));
 INVx1_ASAP7_75t_R _18694_ (.A(_00270_),
    .Y(_13421_));
 NOR2x1_ASAP7_75t_R _18695_ (.A(net352),
    .B(_00272_),
    .Y(_13422_));
 AO21x1_ASAP7_75t_R _18696_ (.A1(net352),
    .A2(_13421_),
    .B(_13422_),
    .Y(_13423_));
 TIEHIx1_ASAP7_75t_R _34914__501 (.H(net501));
 TIEHIx1_ASAP7_75t_R _34913__500 (.H(net500));
 INVx1_ASAP7_75t_R _18699_ (.A(_00276_),
    .Y(_13426_));
 TIEHIx1_ASAP7_75t_R _34912__499 (.H(net499));
 NAND2x1_ASAP7_75t_R _18701_ (.A(net2276),
    .B(_00274_),
    .Y(_13428_));
 OA211x2_ASAP7_75t_R _18702_ (.A1(net352),
    .A2(_13426_),
    .B(_13402_),
    .C(_13428_),
    .Y(_13429_));
 AO21x1_ASAP7_75t_R _18703_ (.A1(_13377_),
    .A2(_13423_),
    .B(_13429_),
    .Y(_13430_));
 TIEHIx1_ASAP7_75t_R _34911__498 (.H(net498));
 TIEHIx1_ASAP7_75t_R _34910__497 (.H(net497));
 NAND2x1_ASAP7_75t_R _18706_ (.A(net352),
    .B(_00269_),
    .Y(_13433_));
 NAND2x1_ASAP7_75t_R _18707_ (.A(net2278),
    .B(_00271_),
    .Y(_13434_));
 TIEHIx1_ASAP7_75t_R _34909__496 (.H(net496));
 NAND2x1_ASAP7_75t_R _18709_ (.A(net2269),
    .B(_00273_),
    .Y(_13436_));
 NAND2x1_ASAP7_75t_R _18710_ (.A(net2278),
    .B(_00275_),
    .Y(_13437_));
 AO33x2_ASAP7_75t_R _18711_ (.A1(_13357_),
    .A2(_13433_),
    .A3(_13434_),
    .B1(_13436_),
    .B2(_13437_),
    .B3(_13366_),
    .Y(_13438_));
 NOR2x2_ASAP7_75t_R _18712_ (.A(net331),
    .B(net328),
    .Y(_13439_));
 TIEHIx1_ASAP7_75t_R _34908__495 (.H(net495));
 OA21x2_ASAP7_75t_R _18714_ (.A1(_13430_),
    .A2(_13438_),
    .B(_13439_),
    .Y(_13441_));
 NOR3x2_ASAP7_75t_R _18715_ (.B(_13419_),
    .C(_13441_),
    .Y(_13442_),
    .A(_13372_));
 TIEHIx1_ASAP7_75t_R _34907__494 (.H(net494));
 NAND2x2_ASAP7_75t_R _18717_ (.A(_01608_),
    .B(_01609_),
    .Y(_13444_));
 OR2x4_ASAP7_75t_R _18718_ (.A(_00277_),
    .B(_13444_),
    .Y(_13445_));
 INVx2_ASAP7_75t_R _18719_ (.A(_01609_),
    .Y(_13446_));
 TIEHIx1_ASAP7_75t_R _34906__493 (.H(net493));
 INVx1_ASAP7_75t_R _18721_ (.A(_00277_),
    .Y(_13448_));
 AO211x2_ASAP7_75t_R _18722_ (.A1(_18554_),
    .A2(_13446_),
    .B(_01608_),
    .C(_13448_),
    .Y(_13449_));
 NAND2x2_ASAP7_75t_R _18723_ (.A(_13445_),
    .B(_13449_),
    .Y(_13450_));
 TIEHIx1_ASAP7_75t_R _34905__492 (.H(net492));
 TIEHIx1_ASAP7_75t_R _34904__491 (.H(net491));
 TIEHIx1_ASAP7_75t_R _34903__490 (.H(net490));
 TIEHIx1_ASAP7_75t_R _34902__489 (.H(net489));
 TIEHIx1_ASAP7_75t_R _34901__488 (.H(net488));
 INVx6_ASAP7_75t_R _18729_ (.A(_00175_),
    .Y(_13456_));
 AND4x2_ASAP7_75t_R _18730_ (.A(_00278_),
    .B(_00279_),
    .C(_00172_),
    .D(_13456_),
    .Y(_13457_));
 TIEHIx1_ASAP7_75t_R _34900__487 (.H(net487));
 CKINVDCx9p33_ASAP7_75t_R _18732_ (.A(_01317_),
    .Y(_13459_));
 CKINVDCx6p67_ASAP7_75t_R _18733_ (.A(_00172_),
    .Y(_13460_));
 TIEHIx1_ASAP7_75t_R _34899__486 (.H(net486));
 TIEHIx1_ASAP7_75t_R _34898__485 (.H(net485));
 OR4x2_ASAP7_75t_R _18736_ (.A(_00278_),
    .B(_00163_),
    .C(_00175_),
    .D(_01746_),
    .Y(_13463_));
 TIEHIx1_ASAP7_75t_R _34897__484 (.H(net484));
 AOI211x1_ASAP7_75t_R _18738_ (.A1(_01713_),
    .A2(_13459_),
    .B(_13460_),
    .C(_13463_),
    .Y(_13465_));
 TIEHIx1_ASAP7_75t_R _34896__483 (.H(net483));
 OR2x2_ASAP7_75t_R _18740_ (.A(_00163_),
    .B(_01746_),
    .Y(_13467_));
 TIEHIx1_ASAP7_75t_R _34895__482 (.H(net482));
 TIEHIx1_ASAP7_75t_R _34894__481 (.H(net481));
 NAND2x2_ASAP7_75t_R _18743_ (.A(_00165_),
    .B(_00168_),
    .Y(_13470_));
 NOR2x1_ASAP7_75t_R _18744_ (.A(_00278_),
    .B(_00172_),
    .Y(_13471_));
 OR4x1_ASAP7_75t_R _18745_ (.A(_00175_),
    .B(_13467_),
    .C(_13470_),
    .D(_13471_),
    .Y(_13472_));
 OR3x4_ASAP7_75t_R _18746_ (.A(_13457_),
    .B(_13465_),
    .C(_13472_),
    .Y(_13473_));
 NOR2x2_ASAP7_75t_R _18747_ (.A(_13450_),
    .B(_13473_),
    .Y(_13474_));
 TIEHIx1_ASAP7_75t_R _34893__480 (.H(net480));
 AND2x6_ASAP7_75t_R _18749_ (.A(_00165_),
    .B(_00168_),
    .Y(_13476_));
 TIEHIx1_ASAP7_75t_R _34892__479 (.H(net479));
 NAND2x1_ASAP7_75t_R _18751_ (.A(_13476_),
    .B(_13465_),
    .Y(_13478_));
 INVx2_ASAP7_75t_R _18752_ (.A(_00278_),
    .Y(_13479_));
 INVx3_ASAP7_75t_R _18753_ (.A(_00168_),
    .Y(_13480_));
 OR5x2_ASAP7_75t_R _18754_ (.A(_13479_),
    .B(_00165_),
    .C(_13480_),
    .D(_00172_),
    .E(_13467_),
    .Y(_13481_));
 AND3x1_ASAP7_75t_R _18755_ (.A(_13445_),
    .B(_13449_),
    .C(_13481_),
    .Y(_13482_));
 CKINVDCx12_ASAP7_75t_R _18756_ (.A(_00281_),
    .Y(_13483_));
 AND2x2_ASAP7_75t_R _18757_ (.A(_00279_),
    .B(_00282_),
    .Y(_13484_));
 NAND2x2_ASAP7_75t_R _18758_ (.A(_13483_),
    .B(_13484_),
    .Y(_13485_));
 NAND2x1_ASAP7_75t_R _18759_ (.A(_00278_),
    .B(_00175_),
    .Y(_13486_));
 OR5x2_ASAP7_75t_R _18760_ (.A(_00165_),
    .B(_00168_),
    .C(_13460_),
    .D(_13467_),
    .E(_13486_),
    .Y(_13487_));
 OR2x2_ASAP7_75t_R _18761_ (.A(_13485_),
    .B(_13487_),
    .Y(_13488_));
 NOR2x2_ASAP7_75t_R _18762_ (.A(_00163_),
    .B(_01746_),
    .Y(_13489_));
 AND2x2_ASAP7_75t_R _18763_ (.A(_13489_),
    .B(_13476_),
    .Y(_13490_));
 TIEHIx1_ASAP7_75t_R _34891__478 (.H(net478));
 AOI211x1_ASAP7_75t_R _18765_ (.A1(_01713_),
    .A2(_13459_),
    .B(_00165_),
    .C(_13463_),
    .Y(_13492_));
 TIEHIx1_ASAP7_75t_R _34890__477 (.H(net477));
 AOI22x1_ASAP7_75t_R _18767_ (.A1(_13457_),
    .A2(_13490_),
    .B1(_13492_),
    .B2(_00172_),
    .Y(_13494_));
 AND4x2_ASAP7_75t_R _18768_ (.A(_13478_),
    .B(_13482_),
    .C(_13488_),
    .D(_13494_),
    .Y(_13495_));
 INVx5_ASAP7_75t_R _18769_ (.A(_00165_),
    .Y(_13496_));
 AND5x2_ASAP7_75t_R _18770_ (.A(_00278_),
    .B(_13496_),
    .C(_00168_),
    .D(_13460_),
    .E(_13489_),
    .Y(_13497_));
 AND2x2_ASAP7_75t_R _18771_ (.A(_00278_),
    .B(_00175_),
    .Y(_13498_));
 NOR2x1_ASAP7_75t_R _18772_ (.A(_00278_),
    .B(_00175_),
    .Y(_13499_));
 AO31x2_ASAP7_75t_R _18773_ (.A1(_13483_),
    .A2(_13484_),
    .A3(_13498_),
    .B(_13499_),
    .Y(_13500_));
 TIEHIx1_ASAP7_75t_R _34889__476 (.H(net476));
 AND4x1_ASAP7_75t_R _18775_ (.A(_13496_),
    .B(_13480_),
    .C(_00172_),
    .D(_13489_),
    .Y(_13502_));
 NAND2x1_ASAP7_75t_R _18776_ (.A(_00168_),
    .B(_00172_),
    .Y(_13503_));
 AOI211x1_ASAP7_75t_R _18777_ (.A1(_01713_),
    .A2(_13459_),
    .B(_13463_),
    .C(_13503_),
    .Y(_13504_));
 AO22x2_ASAP7_75t_R _18778_ (.A1(_13500_),
    .A2(_13502_),
    .B1(_13504_),
    .B2(_13496_),
    .Y(_13505_));
 OR3x1_ASAP7_75t_R _18779_ (.A(_13450_),
    .B(_13497_),
    .C(_13505_),
    .Y(_13506_));
 NOR2x2_ASAP7_75t_R _18780_ (.A(_00277_),
    .B(_13444_),
    .Y(_13507_));
 INVx2_ASAP7_75t_R _18781_ (.A(_18554_),
    .Y(_13508_));
 INVx1_ASAP7_75t_R _18782_ (.A(_01608_),
    .Y(_13509_));
 OA211x2_ASAP7_75t_R _18783_ (.A1(_13508_),
    .A2(_01609_),
    .B(_13509_),
    .C(_00277_),
    .Y(_13510_));
 OR3x1_ASAP7_75t_R _18784_ (.A(_13507_),
    .B(_13510_),
    .C(_13497_),
    .Y(_13511_));
 AO221x1_ASAP7_75t_R _18785_ (.A1(_13476_),
    .A2(_13465_),
    .B1(_13488_),
    .B2(_13494_),
    .C(_13511_),
    .Y(_13512_));
 AOI22x1_ASAP7_75t_R _18786_ (.A1(_13500_),
    .A2(_13502_),
    .B1(_13504_),
    .B2(_13496_),
    .Y(_13513_));
 OA33x2_ASAP7_75t_R _18787_ (.A1(_00184_),
    .A2(_13495_),
    .A3(_13506_),
    .B1(_13512_),
    .B2(_13513_),
    .B3(_00385_),
    .Y(_13514_));
 TIEHIx1_ASAP7_75t_R _34888__475 (.H(net475));
 TIEHIx1_ASAP7_75t_R _34887__474 (.H(net474));
 AND2x2_ASAP7_75t_R _18790_ (.A(_13476_),
    .B(_13465_),
    .Y(_13517_));
 NOR2x1_ASAP7_75t_R _18791_ (.A(_13485_),
    .B(_13487_),
    .Y(_13518_));
 AO32x1_ASAP7_75t_R _18792_ (.A1(_13457_),
    .A2(_13489_),
    .A3(_13476_),
    .B1(_13492_),
    .B2(_00172_),
    .Y(_13519_));
 OR4x2_ASAP7_75t_R _18793_ (.A(_13517_),
    .B(_13511_),
    .C(_13518_),
    .D(_13519_),
    .Y(_13520_));
 OR2x6_ASAP7_75t_R _18794_ (.A(_13450_),
    .B(_13473_),
    .Y(_13521_));
 OA21x2_ASAP7_75t_R _18795_ (.A1(net2269),
    .A2(_13520_),
    .B(_13521_),
    .Y(_13522_));
 AO22x2_ASAP7_75t_R _18796_ (.A1(_13442_),
    .A2(_13474_),
    .B1(_13514_),
    .B2(_13522_),
    .Y(_13523_));
 TIEHIx1_ASAP7_75t_R _34886__473 (.H(net473));
 INVx8_ASAP7_75t_R _18798_ (.A(_13523_),
    .Y(_13525_));
 TIEHIx1_ASAP7_75t_R _34885__472 (.H(net472));
 TIEHIx1_ASAP7_75t_R _34884__471 (.H(net471));
 TIEHIx1_ASAP7_75t_R _34883__470 (.H(net470));
 TIEHIx1_ASAP7_75t_R _34882__469 (.H(net469));
 INVx5_ASAP7_75t_R _18803_ (.A(_01743_),
    .Y(_13528_));
 TIEHIx1_ASAP7_75t_R _34881__468 (.H(net468));
 TIELOx1_ASAP7_75t_R _36799__466 (.L(net466));
 AND2x6_ASAP7_75t_R _18806_ (.A(_00283_),
    .B(_01742_),
    .Y(_13531_));
 AND3x2_ASAP7_75t_R _18807_ (.A(_00280_),
    .B(_01740_),
    .C(_01741_),
    .Y(_13532_));
 AND2x2_ASAP7_75t_R _18808_ (.A(_13531_),
    .B(_13532_),
    .Y(_13533_));
 AND3x4_ASAP7_75t_R _18809_ (.A(_01739_),
    .B(_13528_),
    .C(_13533_),
    .Y(_13534_));
 TIELOx1_ASAP7_75t_R _36798__465 (.L(net465));
 TIELOx1_ASAP7_75t_R _36767__464 (.L(net464));
 AND5x2_ASAP7_75t_R _18812_ (.A(_00278_),
    .B(_13460_),
    .C(_13456_),
    .D(_13489_),
    .E(_13476_),
    .Y(_13537_));
 NAND2x2_ASAP7_75t_R _18813_ (.A(_13534_),
    .B(_13537_),
    .Y(_13538_));
 TIELOx1_ASAP7_75t_R _36766__463 (.L(net463));
 TIELOx1_ASAP7_75t_R _36765__462 (.L(net462));
 TIELOx1_ASAP7_75t_R ibex_core_461 (.L(net461));
 BUFx16f_ASAP7_75t_R load_slew460 (.A(net2385),
    .Y(net460));
 BUFx16f_ASAP7_75t_R load_slew459 (.A(net2385),
    .Y(net459));
 BUFx16f_ASAP7_75t_R max_length458 (.A(net459),
    .Y(net458));
 BUFx16f_ASAP7_75t_R load_slew457 (.A(net459),
    .Y(net457));
 NAND2x1_ASAP7_75t_R _18821_ (.A(_00279_),
    .B(_00282_),
    .Y(_13546_));
 AND5x2_ASAP7_75t_R _18822_ (.A(_13496_),
    .B(_13480_),
    .C(_00172_),
    .D(_13489_),
    .E(_13498_),
    .Y(_13547_));
 NAND2x1_ASAP7_75t_R _18823_ (.A(_13546_),
    .B(_13547_),
    .Y(_13548_));
 AND3x1_ASAP7_75t_R _18824_ (.A(_13496_),
    .B(_00172_),
    .C(_13489_),
    .Y(_13549_));
 AO21x1_ASAP7_75t_R _18825_ (.A1(_13480_),
    .A2(_13498_),
    .B(_13499_),
    .Y(_13550_));
 OA21x2_ASAP7_75t_R _18826_ (.A1(_00278_),
    .A2(_13456_),
    .B(_00172_),
    .Y(_13551_));
 AND4x1_ASAP7_75t_R _18827_ (.A(_00278_),
    .B(_00168_),
    .C(_13460_),
    .D(_13489_),
    .Y(_13552_));
 AO221x2_ASAP7_75t_R _18828_ (.A1(_13549_),
    .A2(_13550_),
    .B1(_13551_),
    .B2(_13490_),
    .C(_13552_),
    .Y(_13553_));
 AND2x2_ASAP7_75t_R _18829_ (.A(_13548_),
    .B(_13553_),
    .Y(_13554_));
 AND4x2_ASAP7_75t_R _18830_ (.A(_00278_),
    .B(_13460_),
    .C(_13489_),
    .D(_13476_),
    .Y(_13555_));
 BUFx16f_ASAP7_75t_R load_slew456 (.A(net457),
    .Y(net456));
 BUFx16f_ASAP7_75t_R load_slew455 (.A(net456),
    .Y(net455));
 NAND2x1_ASAP7_75t_R _18833_ (.A(_00279_),
    .B(_00281_),
    .Y(_13558_));
 INVx5_ASAP7_75t_R _18834_ (.A(_00282_),
    .Y(_13559_));
 BUFx16f_ASAP7_75t_R load_slew454 (.A(net456),
    .Y(net454));
 AND4x2_ASAP7_75t_R _18836_ (.A(_00280_),
    .B(_01740_),
    .C(_01741_),
    .D(_01742_),
    .Y(_13561_));
 NOR2x2_ASAP7_75t_R _18837_ (.A(_00279_),
    .B(_00281_),
    .Y(_13562_));
 OAI21x1_ASAP7_75t_R _18838_ (.A1(_13559_),
    .A2(_13561_),
    .B(_13562_),
    .Y(_13563_));
 AND4x2_ASAP7_75t_R _18839_ (.A(_00175_),
    .B(_13555_),
    .C(_13558_),
    .D(_13563_),
    .Y(_13564_));
 NAND2x1_ASAP7_75t_R _18840_ (.A(_13531_),
    .B(_13532_),
    .Y(_13565_));
 XOR2x1_ASAP7_75t_R _18841_ (.A(_00279_),
    .Y(_13566_),
    .B(_00281_));
 AOI21x1_ASAP7_75t_R _18842_ (.A1(_00282_),
    .A2(_01743_),
    .B(_01739_),
    .Y(_13567_));
 AO21x1_ASAP7_75t_R _18843_ (.A1(_01743_),
    .A2(_13566_),
    .B(_13567_),
    .Y(_13568_));
 OA21x2_ASAP7_75t_R _18844_ (.A1(_13565_),
    .A2(_13568_),
    .B(_13537_),
    .Y(_13569_));
 CKINVDCx11_ASAP7_75t_R _18845_ (.A(_00279_),
    .Y(_13570_));
 AND2x2_ASAP7_75t_R _18846_ (.A(_13570_),
    .B(_00281_),
    .Y(_13571_));
 INVx1_ASAP7_75t_R _18847_ (.A(_01713_),
    .Y(_13572_));
 OR5x2_ASAP7_75t_R _18848_ (.A(_13572_),
    .B(_01317_),
    .C(_13460_),
    .D(_13470_),
    .E(_13463_),
    .Y(_13573_));
 AND2x4_ASAP7_75t_R _18849_ (.A(_13483_),
    .B(_00282_),
    .Y(_13574_));
 AOI211x1_ASAP7_75t_R _18850_ (.A1(_13559_),
    .A2(_13571_),
    .B(_13573_),
    .C(_13574_),
    .Y(_13575_));
 NOR3x2_ASAP7_75t_R _18851_ (.B(_13569_),
    .C(_13575_),
    .Y(_13576_),
    .A(_13564_));
 NAND2x2_ASAP7_75t_R _18852_ (.A(_13554_),
    .B(_13576_),
    .Y(_13577_));
 AND2x2_ASAP7_75t_R _18853_ (.A(_13574_),
    .B(_13555_),
    .Y(_13578_));
 AND3x1_ASAP7_75t_R _18854_ (.A(_00283_),
    .B(_01742_),
    .C(_01743_),
    .Y(_13579_));
 OA211x2_ASAP7_75t_R _18855_ (.A1(_13570_),
    .A2(_01739_),
    .B(_13532_),
    .C(_13579_),
    .Y(_13580_));
 OA21x2_ASAP7_75t_R _18856_ (.A1(_00279_),
    .A2(_13561_),
    .B(_00175_),
    .Y(_13581_));
 AO21x1_ASAP7_75t_R _18857_ (.A1(_13456_),
    .A2(_13580_),
    .B(_13581_),
    .Y(_13582_));
 NOR2x1_ASAP7_75t_R _18858_ (.A(_13485_),
    .B(_13573_),
    .Y(_13583_));
 AOI21x1_ASAP7_75t_R _18859_ (.A1(_13578_),
    .A2(_13582_),
    .B(_13583_),
    .Y(_13584_));
 BUFx16f_ASAP7_75t_R load_slew453 (.A(net458),
    .Y(net453));
 AND2x2_ASAP7_75t_R _18861_ (.A(_01713_),
    .B(_13459_),
    .Y(_13586_));
 NOR2x2_ASAP7_75t_R _18862_ (.A(_13460_),
    .B(_13463_),
    .Y(_13587_));
 AND3x1_ASAP7_75t_R _18863_ (.A(_13476_),
    .B(_13586_),
    .C(_13587_),
    .Y(_13588_));
 BUFx16f_ASAP7_75t_R wire452 (.A(net2385),
    .Y(net452));
 NAND2x1_ASAP7_75t_R _18865_ (.A(_00282_),
    .B(_13566_),
    .Y(_13590_));
 AND4x1_ASAP7_75t_R _18866_ (.A(_13570_),
    .B(_01739_),
    .C(_13532_),
    .D(_13579_),
    .Y(_13591_));
 NOR2x2_ASAP7_75t_R _18867_ (.A(_00281_),
    .B(_00282_),
    .Y(_13592_));
 OA211x2_ASAP7_75t_R _18868_ (.A1(_00175_),
    .A2(_13591_),
    .B(_13592_),
    .C(_13555_),
    .Y(_13593_));
 AOI21x1_ASAP7_75t_R _18869_ (.A1(_13588_),
    .A2(_13590_),
    .B(_13593_),
    .Y(_13594_));
 INVx4_ASAP7_75t_R _18870_ (.A(_01739_),
    .Y(_13595_));
 AND2x2_ASAP7_75t_R _18871_ (.A(_00282_),
    .B(_01739_),
    .Y(_13596_));
 AO32x1_ASAP7_75t_R _18872_ (.A1(_00281_),
    .A2(_13595_),
    .A3(_13484_),
    .B1(_13562_),
    .B2(_13596_),
    .Y(_13597_));
 AND3x1_ASAP7_75t_R _18873_ (.A(_00281_),
    .B(_13559_),
    .C(_01739_),
    .Y(_13598_));
 OR2x2_ASAP7_75t_R _18874_ (.A(_13597_),
    .B(_13598_),
    .Y(_13599_));
 AND2x2_ASAP7_75t_R _18875_ (.A(_13532_),
    .B(_13579_),
    .Y(_13600_));
 AND2x2_ASAP7_75t_R _18876_ (.A(_13537_),
    .B(_13600_),
    .Y(_13601_));
 AO32x1_ASAP7_75t_R _18877_ (.A1(_13562_),
    .A2(_13561_),
    .A3(_13596_),
    .B1(_13559_),
    .B2(_00281_),
    .Y(_13602_));
 AND3x1_ASAP7_75t_R _18878_ (.A(_00175_),
    .B(_13555_),
    .C(_13602_),
    .Y(_13603_));
 OA21x2_ASAP7_75t_R _18879_ (.A1(_13570_),
    .A2(_00281_),
    .B(_00282_),
    .Y(_13604_));
 AND4x2_ASAP7_75t_R _18880_ (.A(_13476_),
    .B(_13586_),
    .C(_13587_),
    .D(_13604_),
    .Y(_13605_));
 AO211x2_ASAP7_75t_R _18881_ (.A1(_13599_),
    .A2(_13601_),
    .B(_13603_),
    .C(_13605_),
    .Y(_13606_));
 NAND3x1_ASAP7_75t_R _18882_ (.A(_13584_),
    .B(_13594_),
    .C(_13606_),
    .Y(_13607_));
 AO22x1_ASAP7_75t_R _18883_ (.A1(_13483_),
    .A2(_13595_),
    .B1(_01743_),
    .B2(_13559_),
    .Y(_13608_));
 NAND2x1_ASAP7_75t_R _18884_ (.A(_00279_),
    .B(_13608_),
    .Y(_13609_));
 OA211x2_ASAP7_75t_R _18885_ (.A1(_00279_),
    .A2(_13483_),
    .B(_00282_),
    .C(_01743_),
    .Y(_13610_));
 OA21x2_ASAP7_75t_R _18886_ (.A1(_01739_),
    .A2(_13610_),
    .B(_13533_),
    .Y(_13611_));
 NAND2x2_ASAP7_75t_R _18887_ (.A(_13456_),
    .B(_13555_),
    .Y(_13612_));
 AO21x2_ASAP7_75t_R _18888_ (.A1(_13609_),
    .A2(_13611_),
    .B(_13612_),
    .Y(_13613_));
 NAND2x1_ASAP7_75t_R _18889_ (.A(_00279_),
    .B(_13559_),
    .Y(_13614_));
 OR4x1_ASAP7_75t_R _18890_ (.A(_00279_),
    .B(_00281_),
    .C(_13559_),
    .D(_13561_),
    .Y(_13615_));
 OR5x2_ASAP7_75t_R _18891_ (.A(_13479_),
    .B(_00172_),
    .C(_13456_),
    .D(_13467_),
    .E(_13470_),
    .Y(_13616_));
 AO21x1_ASAP7_75t_R _18892_ (.A1(_13614_),
    .A2(_13615_),
    .B(_13616_),
    .Y(_13617_));
 AND4x2_ASAP7_75t_R _18893_ (.A(_13573_),
    .B(_13613_),
    .C(_13617_),
    .D(_13554_),
    .Y(_13618_));
 BUFx16f_ASAP7_75t_R load_slew451 (.A(net452),
    .Y(net451));
 OA21x2_ASAP7_75t_R _18895_ (.A1(_13577_),
    .A2(_13607_),
    .B(_13618_),
    .Y(_13620_));
 BUFx16f_ASAP7_75t_R load_slew450 (.A(net451),
    .Y(net450));
 BUFx16f_ASAP7_75t_R wire449 (.A(net450),
    .Y(net449));
 XNOR2x1_ASAP7_75t_R _18898_ (.B(_13620_),
    .Y(_13623_),
    .A(_13523_));
 BUFx16f_ASAP7_75t_R load_slew448 (.A(net451),
    .Y(net448));
 BUFx16f_ASAP7_75t_R load_slew447 (.A(net451),
    .Y(net447));
 CKINVDCx20_ASAP7_75t_R _18901_ (.A(_00286_),
    .Y(_13626_));
 BUFx16f_ASAP7_75t_R load_slew446 (.A(net447),
    .Y(net446));
 BUFx16f_ASAP7_75t_R load_slew445 (.A(net447),
    .Y(net445));
 BUFx16f_ASAP7_75t_R wire444 (.A(net445),
    .Y(net444));
 INVx13_ASAP7_75t_R _18905_ (.A(net388),
    .Y(_13630_));
 BUFx16f_ASAP7_75t_R load_slew443 (.A(net446),
    .Y(net443));
 BUFx16f_ASAP7_75t_R load_slew442 (.A(net443),
    .Y(net442));
 BUFx16f_ASAP7_75t_R load_slew441 (.A(net460),
    .Y(net441));
 BUFx16f_ASAP7_75t_R load_slew440 (.A(net460),
    .Y(net440));
 BUFx16f_ASAP7_75t_R load_slew439 (.A(net460),
    .Y(net439));
 CKINVDCx20_ASAP7_75t_R _18911_ (.A(net381),
    .Y(_13636_));
 BUFx16f_ASAP7_75t_R load_slew438 (.A(net439),
    .Y(net438));
 INVx1_ASAP7_75t_R _18913_ (.A(_00252_),
    .Y(_13638_));
 BUFx16f_ASAP7_75t_R load_slew437 (.A(net460),
    .Y(net437));
 BUFx16f_ASAP7_75t_R load_slew436 (.A(net437),
    .Y(net436));
 BUFx16f_ASAP7_75t_R load_slew435 (.A(net437),
    .Y(net435));
 BUFx16f_ASAP7_75t_R load_slew434 (.A(_01643_),
    .Y(net434));
 BUFx16f_ASAP7_75t_R load_slew433 (.A(net434),
    .Y(net433));
 BUFx16f_ASAP7_75t_R load_slew432 (.A(_01642_),
    .Y(net432));
 BUFx16f_ASAP7_75t_R load_slew431 (.A(_00662_),
    .Y(net431));
 BUFx16f_ASAP7_75t_R wire430 (.A(net431),
    .Y(net430));
 NAND2x1_ASAP7_75t_R _18922_ (.A(_00250_),
    .B(net393),
    .Y(_13647_));
 BUFx16f_ASAP7_75t_R max_cap429 (.A(_00237_),
    .Y(net429));
 CKINVDCx20_ASAP7_75t_R _18924_ (.A(net419),
    .Y(_13649_));
 BUFx16f_ASAP7_75t_R load_slew428 (.A(_00240_),
    .Y(net428));
 BUFx16f_ASAP7_75t_R load_slew427 (.A(_00290_),
    .Y(net427));
 BUFx16f_ASAP7_75t_R load_slew426 (.A(net2261),
    .Y(net426));
 OA211x2_ASAP7_75t_R _18928_ (.A1(_13638_),
    .A2(net393),
    .B(_13647_),
    .C(net319),
    .Y(_13653_));
 INVx1_ASAP7_75t_R _18929_ (.A(_00251_),
    .Y(_13654_));
 NAND2x1_ASAP7_75t_R _18930_ (.A(_00249_),
    .B(net393),
    .Y(_13655_));
 BUFx16f_ASAP7_75t_R wire425 (.A(net426),
    .Y(net425));
 BUFx16f_ASAP7_75t_R load_slew424 (.A(net425),
    .Y(net424));
 BUFx16f_ASAP7_75t_R load_slew423 (.A(net424),
    .Y(net423));
 BUFx16f_ASAP7_75t_R load_slew422 (.A(net425),
    .Y(net422));
 OA211x2_ASAP7_75t_R _18935_ (.A1(_13654_),
    .A2(net393),
    .B(_13655_),
    .C(net2261),
    .Y(_13660_));
 OR3x1_ASAP7_75t_R _18936_ (.A(_13636_),
    .B(_13653_),
    .C(_13660_),
    .Y(_13661_));
 BUFx16f_ASAP7_75t_R load_slew421 (.A(net422),
    .Y(net421));
 INVx1_ASAP7_75t_R _18938_ (.A(_00260_),
    .Y(_13663_));
 NAND2x1_ASAP7_75t_R _18939_ (.A(_00258_),
    .B(net416),
    .Y(_13664_));
 OA211x2_ASAP7_75t_R _18940_ (.A1(_13663_),
    .A2(net416),
    .B(_13664_),
    .C(net319),
    .Y(_13665_));
 INVx1_ASAP7_75t_R _18941_ (.A(_00259_),
    .Y(_13666_));
 BUFx16f_ASAP7_75t_R max_cap420 (.A(net421),
    .Y(net420));
 NAND2x1_ASAP7_75t_R _18943_ (.A(_00257_),
    .B(net416),
    .Y(_13668_));
 OA211x2_ASAP7_75t_R _18944_ (.A1(_13666_),
    .A2(net416),
    .B(_13668_),
    .C(net426),
    .Y(_13669_));
 OR3x1_ASAP7_75t_R _18945_ (.A(net382),
    .B(_13665_),
    .C(_13669_),
    .Y(_13670_));
 AND3x1_ASAP7_75t_R _18946_ (.A(_13630_),
    .B(_13661_),
    .C(_13670_),
    .Y(_13671_));
 BUFx16f_ASAP7_75t_R load_slew419 (.A(net427),
    .Y(net419));
 BUFx16f_ASAP7_75t_R load_slew418 (.A(net2209),
    .Y(net418));
 BUFx16f_ASAP7_75t_R max_cap417 (.A(net2211),
    .Y(net417));
 CKINVDCx12_ASAP7_75t_R _18950_ (.A(net389),
    .Y(_13675_));
 BUFx12f_ASAP7_75t_R load_slew416 (.A(net417),
    .Y(net416));
 BUFx16f_ASAP7_75t_R load_slew415 (.A(net417),
    .Y(net415));
 BUFx16f_ASAP7_75t_R load_slew414 (.A(net2210),
    .Y(net414));
 NAND2x1_ASAP7_75t_R _18954_ (.A(_00248_),
    .B(_13675_),
    .Y(_13679_));
 BUFx16f_ASAP7_75t_R load_slew413 (.A(net414),
    .Y(net413));
 BUFx16f_ASAP7_75t_R max_cap412 (.A(net413),
    .Y(net412));
 BUFx16f_ASAP7_75t_R max_cap411 (.A(net414),
    .Y(net411));
 BUFx16f_ASAP7_75t_R max_cap410 (.A(net414),
    .Y(net410));
 BUFx12f_ASAP7_75t_R load_slew409 (.A(net411),
    .Y(net409));
 NAND2x1_ASAP7_75t_R _18960_ (.A(net416),
    .B(_01708_),
    .Y(_13685_));
 BUFx16f_ASAP7_75t_R load_slew408 (.A(net411),
    .Y(net408));
 AND2x2_ASAP7_75t_R _18962_ (.A(net2262),
    .B(_13675_),
    .Y(_13687_));
 AO32x1_ASAP7_75t_R _18963_ (.A1(net319),
    .A2(_13679_),
    .A3(_13685_),
    .B1(_13687_),
    .B2(_13412_),
    .Y(_13688_));
 BUFx16f_ASAP7_75t_R max_cap407 (.A(net408),
    .Y(net407));
 BUFx16f_ASAP7_75t_R load_slew406 (.A(net408),
    .Y(net406));
 BUFx16f_ASAP7_75t_R load_slew405 (.A(net406),
    .Y(net405));
 BUFx16f_ASAP7_75t_R load_slew404 (.A(net405),
    .Y(net404));
 BUFx16f_ASAP7_75t_R load_slew403 (.A(net404),
    .Y(net403));
 BUFx16f_ASAP7_75t_R max_cap402 (.A(net403),
    .Y(net402));
 BUFx12f_ASAP7_75t_R load_slew401 (.A(net407),
    .Y(net401));
 BUFx16f_ASAP7_75t_R wire400 (.A(net401),
    .Y(net400));
 BUFx16f_ASAP7_75t_R load_slew399 (.A(net400),
    .Y(net399));
 NAND2x1_ASAP7_75t_R _18973_ (.A(_00253_),
    .B(net2261),
    .Y(_13698_));
 OA211x2_ASAP7_75t_R _18974_ (.A1(_13380_),
    .A2(net2261),
    .B(net417),
    .C(_13698_),
    .Y(_13699_));
 INVx1_ASAP7_75t_R _18975_ (.A(_00256_),
    .Y(_13700_));
 BUFx16f_ASAP7_75t_R max_cap398 (.A(net410),
    .Y(net398));
 NAND2x1_ASAP7_75t_R _18977_ (.A(_00255_),
    .B(net2261),
    .Y(_13702_));
 OA211x2_ASAP7_75t_R _18978_ (.A1(_13700_),
    .A2(net2261),
    .B(_13675_),
    .C(_13702_),
    .Y(_13703_));
 OR3x1_ASAP7_75t_R _18979_ (.A(net382),
    .B(_13699_),
    .C(_13703_),
    .Y(_13704_));
 BUFx16f_ASAP7_75t_R load_slew397 (.A(net398),
    .Y(net397));
 BUFx16f_ASAP7_75t_R load_slew396 (.A(net398),
    .Y(net396));
 BUFx16f_ASAP7_75t_R load_slew395 (.A(net396),
    .Y(net395));
 BUFx16f_ASAP7_75t_R wire394 (.A(net395),
    .Y(net394));
 BUFx16f_ASAP7_75t_R load_slew393 (.A(net418),
    .Y(net393));
 OA211x2_ASAP7_75t_R _18985_ (.A1(_13636_),
    .A2(_13688_),
    .B(_13704_),
    .C(net387),
    .Y(_13710_));
 OR3x4_ASAP7_75t_R _18986_ (.A(_13626_),
    .B(_13671_),
    .C(_13710_),
    .Y(_13711_));
 BUFx16f_ASAP7_75t_R load_slew392 (.A(net418),
    .Y(net392));
 BUFx16f_ASAP7_75t_R wire391 (.A(net393),
    .Y(net391));
 BUFx16f_ASAP7_75t_R max_cap390 (.A(net391),
    .Y(net390));
 BUFx12f_ASAP7_75t_R load_slew389 (.A(net391),
    .Y(net389));
 NAND2x1_ASAP7_75t_R _18991_ (.A(_00266_),
    .B(net413),
    .Y(_13716_));
 OA211x2_ASAP7_75t_R _18992_ (.A1(_13348_),
    .A2(net413),
    .B(_13716_),
    .C(net318),
    .Y(_13717_));
 INVx1_ASAP7_75t_R _18993_ (.A(_00267_),
    .Y(_13718_));
 BUFx12f_ASAP7_75t_R load_slew388 (.A(_00288_),
    .Y(net388));
 BUFx16f_ASAP7_75t_R load_slew387 (.A(net2301),
    .Y(net387));
 BUFx16f_ASAP7_75t_R load_slew386 (.A(net2301),
    .Y(net386));
 NAND2x1_ASAP7_75t_R _18997_ (.A(_00265_),
    .B(net413),
    .Y(_13722_));
 OA211x2_ASAP7_75t_R _18998_ (.A1(_13718_),
    .A2(net413),
    .B(_13722_),
    .C(net425),
    .Y(_13723_));
 OR3x1_ASAP7_75t_R _18999_ (.A(_13636_),
    .B(_13717_),
    .C(_13723_),
    .Y(_13724_));
 INVx1_ASAP7_75t_R _19000_ (.A(_00274_),
    .Y(_13725_));
 BUFx16f_ASAP7_75t_R max_cap385 (.A(net386),
    .Y(net385));
 BUFx16f_ASAP7_75t_R load_slew384 (.A(net385),
    .Y(net384));
 BUFx12f_ASAP7_75t_R load_slew383 (.A(net385),
    .Y(net383));
 BUFx16f_ASAP7_75t_R load_slew382 (.A(_00287_),
    .Y(net382));
 BUFx16f_ASAP7_75t_R max_cap381 (.A(net382),
    .Y(net381));
 NAND2x1_ASAP7_75t_R _19006_ (.A(_00273_),
    .B(net425),
    .Y(_13731_));
 OA211x2_ASAP7_75t_R _19007_ (.A1(_13725_),
    .A2(net425),
    .B(net398),
    .C(_13731_),
    .Y(_13732_));
 NAND2x1_ASAP7_75t_R _19008_ (.A(_00275_),
    .B(net425),
    .Y(_13733_));
 OA211x2_ASAP7_75t_R _19009_ (.A1(_13426_),
    .A2(net424),
    .B(net316),
    .C(_13733_),
    .Y(_13734_));
 OR3x1_ASAP7_75t_R _19010_ (.A(net380),
    .B(_13732_),
    .C(_13734_),
    .Y(_13735_));
 AND3x1_ASAP7_75t_R _19011_ (.A(net321),
    .B(_13724_),
    .C(_13735_),
    .Y(_13736_));
 BUFx16f_ASAP7_75t_R wire380 (.A(net382),
    .Y(net380));
 BUFx12_ASAP7_75t_R load_slew379 (.A(net380),
    .Y(net379));
 BUFx16f_ASAP7_75t_R load_slew378 (.A(_00286_),
    .Y(net378));
 INVx1_ASAP7_75t_R _19015_ (.A(_00261_),
    .Y(_13740_));
 BUFx16f_ASAP7_75t_R load_slew377 (.A(net378),
    .Y(net377));
 BUFx16f_ASAP7_75t_R load_slew376 (.A(_00246_),
    .Y(net376));
 BUFx16f_ASAP7_75t_R wire375 (.A(net376),
    .Y(net375));
 NOR2x1_ASAP7_75t_R _19019_ (.A(_00263_),
    .B(net416),
    .Y(_13744_));
 AO21x1_ASAP7_75t_R _19020_ (.A1(_13740_),
    .A2(net416),
    .B(_13744_),
    .Y(_13745_));
 BUFx16f_ASAP7_75t_R load_slew374 (.A(net375),
    .Y(net374));
 BUFx16f_ASAP7_75t_R load_slew373 (.A(net374),
    .Y(net373));
 BUFx16f_ASAP7_75t_R load_slew372 (.A(net373),
    .Y(net372));
 BUFx12f_ASAP7_75t_R load_slew371 (.A(net372),
    .Y(net371));
 BUFx16f_ASAP7_75t_R load_slew370 (.A(net376),
    .Y(net370));
 NAND2x1_ASAP7_75t_R _19026_ (.A(_00262_),
    .B(net416),
    .Y(_13751_));
 BUFx16f_ASAP7_75t_R load_slew369 (.A(net370),
    .Y(net369));
 BUFx16f_ASAP7_75t_R load_slew368 (.A(net2297),
    .Y(net368));
 OA211x2_ASAP7_75t_R _19029_ (.A1(_13340_),
    .A2(net416),
    .B(_13751_),
    .C(net319),
    .Y(_13754_));
 AO21x1_ASAP7_75t_R _19030_ (.A1(net425),
    .A2(_13745_),
    .B(_13754_),
    .Y(_13755_));
 NAND2x1_ASAP7_75t_R _19031_ (.A(_00269_),
    .B(net424),
    .Y(_13756_));
 OA211x2_ASAP7_75t_R _19032_ (.A1(_13421_),
    .A2(net424),
    .B(net410),
    .C(_13756_),
    .Y(_13757_));
 INVx1_ASAP7_75t_R _19033_ (.A(_00272_),
    .Y(_13758_));
 BUFx16f_ASAP7_75t_R load_slew367 (.A(net2297),
    .Y(net367));
 BUFx16f_ASAP7_75t_R load_slew366 (.A(net367),
    .Y(net366));
 BUFx16f_ASAP7_75t_R load_slew365 (.A(net366),
    .Y(net365));
 NAND2x1_ASAP7_75t_R _19037_ (.A(_00271_),
    .B(net424),
    .Y(_13762_));
 OA211x2_ASAP7_75t_R _19038_ (.A1(_13758_),
    .A2(net424),
    .B(net316),
    .C(_13762_),
    .Y(_13763_));
 OR3x1_ASAP7_75t_R _19039_ (.A(net380),
    .B(_13757_),
    .C(_13763_),
    .Y(_13764_));
 OA211x2_ASAP7_75t_R _19040_ (.A1(_13636_),
    .A2(_13755_),
    .B(_13764_),
    .C(net386),
    .Y(_13765_));
 OR3x4_ASAP7_75t_R _19041_ (.A(net378),
    .B(_13736_),
    .C(_13765_),
    .Y(_13766_));
 AND2x4_ASAP7_75t_R _19042_ (.A(_13711_),
    .B(_13766_),
    .Y(_13767_));
 BUFx16f_ASAP7_75t_R load_slew364 (.A(net365),
    .Y(net364));
 BUFx16f_ASAP7_75t_R max_cap363 (.A(net364),
    .Y(net363));
 BUFx16f_ASAP7_75t_R load_slew362 (.A(net364),
    .Y(net362));
 AND3x4_ASAP7_75t_R _19046_ (.A(_00285_),
    .B(_01357_),
    .C(_01727_),
    .Y(_13771_));
 AND2x6_ASAP7_75t_R _19047_ (.A(_00284_),
    .B(_13771_),
    .Y(_13772_));
 BUFx16f_ASAP7_75t_R load_slew361 (.A(net362),
    .Y(net361));
 BUFx16f_ASAP7_75t_R load_slew360 (.A(net363),
    .Y(net360));
 CKINVDCx20_ASAP7_75t_R _19050_ (.A(_00285_),
    .Y(_13775_));
 BUFx16f_ASAP7_75t_R max_cap359 (.A(net360),
    .Y(net359));
 BUFx16f_ASAP7_75t_R load_slew358 (.A(net359),
    .Y(net358));
 NAND2x2_ASAP7_75t_R _19053_ (.A(_01357_),
    .B(_01727_),
    .Y(_13778_));
 BUFx16f_ASAP7_75t_R max_cap357 (.A(net358),
    .Y(net357));
 AO221x1_ASAP7_75t_R _19055_ (.A1(_13775_),
    .A2(_00291_),
    .B1(_01451_),
    .B2(_13778_),
    .C(_13538_),
    .Y(_13780_));
 AOI21x1_ASAP7_75t_R _19056_ (.A1(_13442_),
    .A2(_13772_),
    .B(_13780_),
    .Y(_13781_));
 OA21x2_ASAP7_75t_R _19057_ (.A1(_00284_),
    .A2(_13767_),
    .B(_13781_),
    .Y(_13782_));
 AOI21x1_ASAP7_75t_R _19058_ (.A1(_13538_),
    .A2(_13623_),
    .B(_13782_),
    .Y(_17755_));
 INVx1_ASAP7_75t_R _19059_ (.A(_17755_),
    .Y(_16715_));
 INVx2_ASAP7_75t_R _19060_ (.A(_01720_),
    .Y(\cs_registers_i.pc_id_i[1] ));
 BUFx16f_ASAP7_75t_R load_slew356 (.A(net357),
    .Y(net356));
 OR3x4_ASAP7_75t_R _19062_ (.A(_00172_),
    .B(_13470_),
    .C(_13463_),
    .Y(_13784_));
 NAND2x1_ASAP7_75t_R _19063_ (.A(_13487_),
    .B(_13784_),
    .Y(_13785_));
 OR2x2_ASAP7_75t_R _19064_ (.A(_13463_),
    .B(_13503_),
    .Y(_13786_));
 OR3x1_ASAP7_75t_R _19065_ (.A(_13479_),
    .B(_13467_),
    .C(_13470_),
    .Y(_13787_));
 AND4x2_ASAP7_75t_R _19066_ (.A(_13487_),
    .B(_13786_),
    .C(_13784_),
    .D(_13787_),
    .Y(_13788_));
 OR4x1_ASAP7_75t_R _19067_ (.A(_00278_),
    .B(_00168_),
    .C(_13460_),
    .D(_00175_),
    .Y(_13789_));
 OR3x1_ASAP7_75t_R _19068_ (.A(_13480_),
    .B(_00172_),
    .C(_13486_),
    .Y(_13790_));
 OR3x1_ASAP7_75t_R _19069_ (.A(_00163_),
    .B(_00165_),
    .C(_01746_),
    .Y(_13791_));
 AO21x1_ASAP7_75t_R _19070_ (.A1(_13789_),
    .A2(_13790_),
    .B(_13791_),
    .Y(_13792_));
 AO211x2_ASAP7_75t_R _19071_ (.A1(_13559_),
    .A2(_13547_),
    .B(_13510_),
    .C(_13507_),
    .Y(_13793_));
 AOI221x1_ASAP7_75t_R _19072_ (.A1(_13570_),
    .A2(_13785_),
    .B1(_13788_),
    .B2(_13792_),
    .C(_13793_),
    .Y(_13794_));
 BUFx16f_ASAP7_75t_R load_slew355 (.A(net358),
    .Y(net355));
 BUFx16f_ASAP7_75t_R load_slew354 (.A(net355),
    .Y(net354));
 NAND2x2_ASAP7_75t_R _19075_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(_13794_),
    .Y(_13797_));
 BUFx12f_ASAP7_75t_R load_slew353 (.A(net354),
    .Y(net353));
 BUFx16f_ASAP7_75t_R load_slew352 (.A(net365),
    .Y(net352));
 BUFx16f_ASAP7_75t_R load_slew351 (.A(net352),
    .Y(net351));
 NOR3x2_ASAP7_75t_R _19079_ (.B(_00163_),
    .C(_01746_),
    .Y(_13801_),
    .A(_00278_));
 AND4x2_ASAP7_75t_R _19080_ (.A(_13460_),
    .B(_13456_),
    .C(_13476_),
    .D(_13801_),
    .Y(_13802_));
 NAND3x2_ASAP7_75t_R _19081_ (.B(_00281_),
    .C(_00282_),
    .Y(_13803_),
    .A(_00279_));
 NAND2x2_ASAP7_75t_R _19082_ (.A(_13802_),
    .B(_13803_),
    .Y(_13804_));
 OR3x1_ASAP7_75t_R _19083_ (.A(net2212),
    .B(_13794_),
    .C(_13804_),
    .Y(_13805_));
 AO221x2_ASAP7_75t_R _19084_ (.A1(_13570_),
    .A2(_13802_),
    .B1(_13803_),
    .B2(_13547_),
    .C(_13504_),
    .Y(_13806_));
 AND2x6_ASAP7_75t_R _19085_ (.A(_13445_),
    .B(_13449_),
    .Y(_13807_));
 OAI21x1_ASAP7_75t_R _19086_ (.A1(_13788_),
    .A2(_13806_),
    .B(_13807_),
    .Y(_13808_));
 AOI21x1_ASAP7_75t_R _19087_ (.A1(_13797_),
    .A2(_13805_),
    .B(_13808_),
    .Y(_13809_));
 AND2x6_ASAP7_75t_R _19088_ (.A(_13808_),
    .B(_13794_),
    .Y(_13810_));
 BUFx16f_ASAP7_75t_R wire350 (.A(net351),
    .Y(net350));
 BUFx16f_ASAP7_75t_R load_slew349 (.A(net351),
    .Y(net349));
 INVx1_ASAP7_75t_R _19091_ (.A(_01640_),
    .Y(_13813_));
 AO32x2_ASAP7_75t_R _19092_ (.A1(_13711_),
    .A2(_13766_),
    .A3(_13810_),
    .B1(_13450_),
    .B2(_13813_),
    .Y(_13814_));
 NOR2x2_ASAP7_75t_R _19093_ (.A(_13809_),
    .B(_13814_),
    .Y(_18332_));
 AND2x6_ASAP7_75t_R _19094_ (.A(_01357_),
    .B(_01727_),
    .Y(_13815_));
 BUFx16f_ASAP7_75t_R load_slew348 (.A(net367),
    .Y(net348));
 AND2x6_ASAP7_75t_R _19096_ (.A(_13534_),
    .B(_13537_),
    .Y(_13817_));
 BUFx16f_ASAP7_75t_R load_slew347 (.A(net348),
    .Y(net347));
 BUFx16f_ASAP7_75t_R load_slew346 (.A(net2143),
    .Y(net346));
 BUFx16f_ASAP7_75t_R max_cap345 (.A(net368),
    .Y(net345));
 BUFx16f_ASAP7_75t_R load_slew344 (.A(net368),
    .Y(net344));
 OA21x2_ASAP7_75t_R _19101_ (.A1(_00291_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_13822_));
 AOI21x1_ASAP7_75t_R _19102_ (.A1(_13538_),
    .A2(_18332_),
    .B(_13822_),
    .Y(_17756_));
 INVx1_ASAP7_75t_R _19103_ (.A(_17756_),
    .Y(_16716_));
 INVx1_ASAP7_75t_R _19104_ (.A(_00301_),
    .Y(_13823_));
 BUFx16f_ASAP7_75t_R load_slew343 (.A(net368),
    .Y(net343));
 NAND2x1_ASAP7_75t_R _19106_ (.A(net2298),
    .B(_00299_),
    .Y(_13825_));
 BUFx16f_ASAP7_75t_R max_cap342 (.A(net345),
    .Y(net342));
 OA211x2_ASAP7_75t_R _19108_ (.A1(net2248),
    .A2(_13823_),
    .B(_13825_),
    .C(net375),
    .Y(_13827_));
 INVx1_ASAP7_75t_R _19109_ (.A(_00302_),
    .Y(_13828_));
 NAND2x1_ASAP7_75t_R _19110_ (.A(net2248),
    .B(_00300_),
    .Y(_13829_));
 OA211x2_ASAP7_75t_R _19111_ (.A1(net2248),
    .A2(_13828_),
    .B(_13829_),
    .C(net323),
    .Y(_13830_));
 OR3x1_ASAP7_75t_R _19112_ (.A(_13350_),
    .B(_13827_),
    .C(_13830_),
    .Y(_13831_));
 BUFx16f_ASAP7_75t_R max_cap341 (.A(net342),
    .Y(net341));
 INVx1_ASAP7_75t_R _19114_ (.A(_00305_),
    .Y(_13833_));
 NAND2x1_ASAP7_75t_R _19115_ (.A(net2299),
    .B(_00303_),
    .Y(_13834_));
 OA211x2_ASAP7_75t_R _19116_ (.A1(net2297),
    .A2(_13833_),
    .B(_13834_),
    .C(net376),
    .Y(_13835_));
 INVx1_ASAP7_75t_R _19117_ (.A(_00306_),
    .Y(_13836_));
 NAND2x1_ASAP7_75t_R _19118_ (.A(net368),
    .B(_00304_),
    .Y(_13837_));
 OA211x2_ASAP7_75t_R _19119_ (.A1(net2297),
    .A2(_13836_),
    .B(_13837_),
    .C(net323),
    .Y(_13838_));
 OR3x1_ASAP7_75t_R _19120_ (.A(net2359),
    .B(_13835_),
    .C(_13838_),
    .Y(_13839_));
 AO21x1_ASAP7_75t_R _19121_ (.A1(_13831_),
    .A2(_13839_),
    .B(net329),
    .Y(_13840_));
 BUFx12f_ASAP7_75t_R load_slew340 (.A(net342),
    .Y(net340));
 AND2x2_ASAP7_75t_R _19123_ (.A(net345),
    .B(_00295_),
    .Y(_13842_));
 AO21x1_ASAP7_75t_R _19124_ (.A1(net326),
    .A2(_00297_),
    .B(_13842_),
    .Y(_13843_));
 AND2x2_ASAP7_75t_R _19125_ (.A(net2143),
    .B(_00296_),
    .Y(_13844_));
 AO21x1_ASAP7_75t_R _19126_ (.A1(net326),
    .A2(_00298_),
    .B(_13844_),
    .Y(_13845_));
 AOI22x1_ASAP7_75t_R _19127_ (.A1(_13366_),
    .A2(_13843_),
    .B1(_13845_),
    .B2(_13402_),
    .Y(_13846_));
 INVx1_ASAP7_75t_R _19128_ (.A(_00293_),
    .Y(_13847_));
 INVx1_ASAP7_75t_R _19129_ (.A(_01709_),
    .Y(_13848_));
 NOR2x1_ASAP7_75t_R _19130_ (.A(net345),
    .B(_00294_),
    .Y(_13849_));
 AO21x1_ASAP7_75t_R _19131_ (.A1(net345),
    .A2(_13848_),
    .B(_13849_),
    .Y(_13850_));
 NAND2x2_ASAP7_75t_R _19132_ (.A(net2358),
    .B(net333),
    .Y(_13851_));
 BUFx16f_ASAP7_75t_R load_slew339 (.A(net341),
    .Y(net339));
 AO221x1_ASAP7_75t_R _19134_ (.A1(_13847_),
    .A2(net2244),
    .B1(_13850_),
    .B2(net323),
    .C(_13851_),
    .Y(_13853_));
 BUFx12f_ASAP7_75t_R load_slew338 (.A(_01744_),
    .Y(net338));
 OA211x2_ASAP7_75t_R _19136_ (.A1(_13373_),
    .A2(_13846_),
    .B(_13853_),
    .C(net328),
    .Y(_13855_));
 INVx1_ASAP7_75t_R _19137_ (.A(_00321_),
    .Y(_13856_));
 NAND2x1_ASAP7_75t_R _19138_ (.A(net368),
    .B(_00319_),
    .Y(_13857_));
 OA211x2_ASAP7_75t_R _19139_ (.A1(net368),
    .A2(_13856_),
    .B(_13857_),
    .C(_13350_),
    .Y(_13858_));
 INVx1_ASAP7_75t_R _19140_ (.A(_00317_),
    .Y(_13859_));
 NAND2x1_ASAP7_75t_R _19141_ (.A(net368),
    .B(_00315_),
    .Y(_13860_));
 OA211x2_ASAP7_75t_R _19142_ (.A1(net368),
    .A2(_13859_),
    .B(_13860_),
    .C(net338),
    .Y(_13861_));
 OR3x1_ASAP7_75t_R _19143_ (.A(net323),
    .B(_13858_),
    .C(_13861_),
    .Y(_13862_));
 BUFx16f_ASAP7_75t_R load_slew337 (.A(net338),
    .Y(net337));
 INVx1_ASAP7_75t_R _19145_ (.A(_00322_),
    .Y(_13864_));
 NAND2x1_ASAP7_75t_R _19146_ (.A(net368),
    .B(_00320_),
    .Y(_13865_));
 OA211x2_ASAP7_75t_R _19147_ (.A1(net368),
    .A2(_13864_),
    .B(_13865_),
    .C(_13350_),
    .Y(_13866_));
 INVx1_ASAP7_75t_R _19148_ (.A(_00318_),
    .Y(_13867_));
 NAND2x1_ASAP7_75t_R _19149_ (.A(net368),
    .B(_00316_),
    .Y(_13868_));
 OA211x2_ASAP7_75t_R _19150_ (.A1(net368),
    .A2(_13867_),
    .B(_13868_),
    .C(net338),
    .Y(_13869_));
 OR3x1_ASAP7_75t_R _19151_ (.A(net376),
    .B(_13866_),
    .C(_13869_),
    .Y(_13870_));
 INVx1_ASAP7_75t_R _19152_ (.A(_00313_),
    .Y(_13871_));
 NAND2x1_ASAP7_75t_R _19153_ (.A(net2144),
    .B(_00311_),
    .Y(_13872_));
 OA211x2_ASAP7_75t_R _19154_ (.A1(net2143),
    .A2(_13871_),
    .B(_13872_),
    .C(_13350_),
    .Y(_13873_));
 INVx1_ASAP7_75t_R _19155_ (.A(_00309_),
    .Y(_13874_));
 NAND2x1_ASAP7_75t_R _19156_ (.A(net342),
    .B(_00307_),
    .Y(_13875_));
 OA211x2_ASAP7_75t_R _19157_ (.A1(net342),
    .A2(_13874_),
    .B(_13875_),
    .C(net337),
    .Y(_13876_));
 OR3x1_ASAP7_75t_R _19158_ (.A(net323),
    .B(_13873_),
    .C(_13876_),
    .Y(_13877_));
 INVx1_ASAP7_75t_R _19159_ (.A(_00314_),
    .Y(_13878_));
 NAND2x1_ASAP7_75t_R _19160_ (.A(net346),
    .B(_00312_),
    .Y(_13879_));
 OA211x2_ASAP7_75t_R _19161_ (.A1(net2143),
    .A2(_13878_),
    .B(_13879_),
    .C(_13350_),
    .Y(_13880_));
 INVx1_ASAP7_75t_R _19162_ (.A(_00310_),
    .Y(_13881_));
 NAND2x1_ASAP7_75t_R _19163_ (.A(net2143),
    .B(_00308_),
    .Y(_13882_));
 OA211x2_ASAP7_75t_R _19164_ (.A1(net2143),
    .A2(_13881_),
    .B(_13882_),
    .C(net337),
    .Y(_13883_));
 OR3x1_ASAP7_75t_R _19165_ (.A(net375),
    .B(_13880_),
    .C(_13883_),
    .Y(_13884_));
 AO33x2_ASAP7_75t_R _19166_ (.A1(_13439_),
    .A2(_13862_),
    .A3(_13870_),
    .B1(_13877_),
    .B2(_13884_),
    .B3(_13356_),
    .Y(_13885_));
 AO21x2_ASAP7_75t_R _19167_ (.A1(_13840_),
    .A2(_13855_),
    .B(_13885_),
    .Y(_13886_));
 BUFx12f_ASAP7_75t_R load_slew336 (.A(net337),
    .Y(net336));
 AND2x6_ASAP7_75t_R _19169_ (.A(_13807_),
    .B(_13513_),
    .Y(_13888_));
 AND4x1_ASAP7_75t_R _19170_ (.A(net323),
    .B(_13521_),
    .C(_13495_),
    .D(_13888_),
    .Y(_13889_));
 INVx2_ASAP7_75t_R _19171_ (.A(_00323_),
    .Y(_13890_));
 OA211x2_ASAP7_75t_R _19172_ (.A1(_13518_),
    .A2(_13519_),
    .B(_13478_),
    .C(_13482_),
    .Y(_13891_));
 AND3x1_ASAP7_75t_R _19173_ (.A(_13890_),
    .B(_13888_),
    .C(_13891_),
    .Y(_13892_));
 AOI211x1_ASAP7_75t_R _19174_ (.A1(_13474_),
    .A2(_13886_),
    .B(_13889_),
    .C(_13892_),
    .Y(_13893_));
 CKINVDCx20_ASAP7_75t_R _19175_ (.A(net303),
    .Y(_13894_));
 BUFx12f_ASAP7_75t_R load_slew335 (.A(net336),
    .Y(net335));
 BUFx16f_ASAP7_75t_R wire334 (.A(net335),
    .Y(net334));
 BUFx6f_ASAP7_75t_R load_slew333 (.A(_00245_),
    .Y(net333));
 BUFx16f_ASAP7_75t_R load_slew332 (.A(_00245_),
    .Y(net332));
 BUFx16f_ASAP7_75t_R load_slew331 (.A(net332),
    .Y(net331));
 BUFx16f_ASAP7_75t_R load_slew330 (.A(net331),
    .Y(net330));
 BUFx16f_ASAP7_75t_R load_slew329 (.A(net333),
    .Y(net329));
 BUFx12f_ASAP7_75t_R load_slew328 (.A(_00244_),
    .Y(net328));
 BUFx16f_ASAP7_75t_R wire327 (.A(net328),
    .Y(net327));
 BUFx16f_ASAP7_75t_R max_length326 (.A(_13359_),
    .Y(net326));
 INVx1_ASAP7_75t_R _19186_ (.A(_00294_),
    .Y(_13903_));
 BUFx16f_ASAP7_75t_R max_length325 (.A(_13376_),
    .Y(net325));
 BUFx16f_ASAP7_75t_R max_length324 (.A(net325),
    .Y(net324));
 NAND2x1_ASAP7_75t_R _19189_ (.A(net417),
    .B(_01709_),
    .Y(_13906_));
 BUFx16f_ASAP7_75t_R max_length323 (.A(_13376_),
    .Y(net323));
 BUFx12f_ASAP7_75t_R load_slew322 (.A(_13402_),
    .Y(net322));
 OA211x2_ASAP7_75t_R _19192_ (.A1(net417),
    .A2(_13903_),
    .B(_13906_),
    .C(_13649_),
    .Y(_13909_));
 AO21x1_ASAP7_75t_R _19193_ (.A1(_13847_),
    .A2(_13687_),
    .B(_13909_),
    .Y(_13910_));
 BUFx16f_ASAP7_75t_R wire321 (.A(_13630_),
    .Y(net321));
 BUFx16f_ASAP7_75t_R max_length320 (.A(net321),
    .Y(net320));
 BUFx16f_ASAP7_75t_R max_length319 (.A(_13649_),
    .Y(net319));
 NAND2x1_ASAP7_75t_R _19197_ (.A(net417),
    .B(_00308_),
    .Y(_13914_));
 OA211x2_ASAP7_75t_R _19198_ (.A1(net417),
    .A2(_13881_),
    .B(_13914_),
    .C(_13649_),
    .Y(_13915_));
 BUFx16f_ASAP7_75t_R max_length318 (.A(net319),
    .Y(net318));
 BUFx16f_ASAP7_75t_R wire317 (.A(_13649_),
    .Y(net317));
 NAND2x1_ASAP7_75t_R _19201_ (.A(net417),
    .B(_00307_),
    .Y(_13918_));
 OA211x2_ASAP7_75t_R _19202_ (.A1(net417),
    .A2(_13874_),
    .B(_13918_),
    .C(net2261),
    .Y(_13919_));
 OR3x1_ASAP7_75t_R _19203_ (.A(_00286_),
    .B(_13915_),
    .C(_13919_),
    .Y(_13920_));
 OA211x2_ASAP7_75t_R _19204_ (.A1(_13626_),
    .A2(_13910_),
    .B(_13920_),
    .C(net387),
    .Y(_13921_));
 BUFx16f_ASAP7_75t_R wire316 (.A(_13675_),
    .Y(net316));
 BUFx16f_ASAP7_75t_R load_slew315 (.A(_14005_),
    .Y(net315));
 BUFx10_ASAP7_75t_R load_slew314 (.A(_02290_),
    .Y(net314));
 BUFx6f_ASAP7_75t_R max_cap313 (.A(net314),
    .Y(net313));
 BUFx12f_ASAP7_75t_R max_length312 (.A(_14015_),
    .Y(net312));
 INVx1_ASAP7_75t_R _19210_ (.A(_00298_),
    .Y(_13927_));
 BUFx16f_ASAP7_75t_R load_slew311 (.A(_14184_),
    .Y(net311));
 NAND2x1_ASAP7_75t_R _19212_ (.A(net417),
    .B(_00296_),
    .Y(_13929_));
 BUFx12f_ASAP7_75t_R max_cap310 (.A(_05570_),
    .Y(net310));
 OA211x2_ASAP7_75t_R _19214_ (.A1(net417),
    .A2(_13927_),
    .B(_13929_),
    .C(_13649_),
    .Y(_13931_));
 BUFx16f_ASAP7_75t_R load_slew309 (.A(_13538_),
    .Y(net309));
 BUFx16f_ASAP7_75t_R load_slew308 (.A(net309),
    .Y(net308));
 INVx1_ASAP7_75t_R _19217_ (.A(_00297_),
    .Y(_13934_));
 BUFx12f_ASAP7_75t_R load_slew307 (.A(_02286_),
    .Y(net307));
 NAND2x1_ASAP7_75t_R _19219_ (.A(net417),
    .B(_00295_),
    .Y(_13936_));
 OA211x2_ASAP7_75t_R _19220_ (.A1(net417),
    .A2(_13934_),
    .B(_13936_),
    .C(_00290_),
    .Y(_13937_));
 OR3x1_ASAP7_75t_R _19221_ (.A(_13626_),
    .B(_13931_),
    .C(_13937_),
    .Y(_13938_));
 NAND2x1_ASAP7_75t_R _19222_ (.A(net417),
    .B(_00312_),
    .Y(_13939_));
 OA211x2_ASAP7_75t_R _19223_ (.A1(net417),
    .A2(_13878_),
    .B(_13939_),
    .C(_13649_),
    .Y(_13940_));
 BUFx12f_ASAP7_75t_R load_slew306 (.A(_02289_),
    .Y(net306));
 NAND2x1_ASAP7_75t_R _19225_ (.A(net417),
    .B(_00311_),
    .Y(_13942_));
 OA211x2_ASAP7_75t_R _19226_ (.A1(net417),
    .A2(_13871_),
    .B(_13942_),
    .C(net2261),
    .Y(_13943_));
 OR3x1_ASAP7_75t_R _19227_ (.A(net378),
    .B(_13940_),
    .C(_13943_),
    .Y(_13944_));
 AND3x1_ASAP7_75t_R _19228_ (.A(_13630_),
    .B(_13938_),
    .C(_13944_),
    .Y(_13945_));
 OR3x2_ASAP7_75t_R _19229_ (.A(_13636_),
    .B(_13921_),
    .C(_13945_),
    .Y(_13946_));
 BUFx16f_ASAP7_75t_R load_slew305 (.A(_13893_),
    .Y(net305));
 NAND2x1_ASAP7_75t_R _19231_ (.A(_00289_),
    .B(_00304_),
    .Y(_13948_));
 OA211x2_ASAP7_75t_R _19232_ (.A1(net2210),
    .A2(_13836_),
    .B(_13948_),
    .C(_13649_),
    .Y(_13949_));
 NAND2x1_ASAP7_75t_R _19233_ (.A(net2378),
    .B(_00303_),
    .Y(_13950_));
 OA211x2_ASAP7_75t_R _19234_ (.A1(net2210),
    .A2(_13833_),
    .B(_13950_),
    .C(_00290_),
    .Y(_13951_));
 OR3x1_ASAP7_75t_R _19235_ (.A(_13626_),
    .B(_13949_),
    .C(_13951_),
    .Y(_13952_));
 BUFx12f_ASAP7_75t_R load_slew304 (.A(net305),
    .Y(net304));
 NAND2x1_ASAP7_75t_R _19237_ (.A(net418),
    .B(_00320_),
    .Y(_13954_));
 OA211x2_ASAP7_75t_R _19238_ (.A1(net418),
    .A2(_13864_),
    .B(_13954_),
    .C(_13649_),
    .Y(_13955_));
 NAND2x1_ASAP7_75t_R _19239_ (.A(net418),
    .B(_00319_),
    .Y(_13956_));
 OA211x2_ASAP7_75t_R _19240_ (.A1(net418),
    .A2(_13856_),
    .B(_13956_),
    .C(_00290_),
    .Y(_13957_));
 OR3x1_ASAP7_75t_R _19241_ (.A(_00286_),
    .B(_13955_),
    .C(_13957_),
    .Y(_13958_));
 AND3x1_ASAP7_75t_R _19242_ (.A(_13630_),
    .B(_13952_),
    .C(_13958_),
    .Y(_13959_));
 BUFx16f_ASAP7_75t_R load_slew303 (.A(net304),
    .Y(net303));
 BUFx12f_ASAP7_75t_R load_slew302 (.A(_14296_),
    .Y(net302));
 BUFx16f_ASAP7_75t_R load_slew301 (.A(_06273_),
    .Y(net301));
 BUFx16f_ASAP7_75t_R load_slew300 (.A(net301),
    .Y(net300));
 NAND2x1_ASAP7_75t_R _19247_ (.A(net2378),
    .B(_00300_),
    .Y(_13964_));
 OA211x2_ASAP7_75t_R _19248_ (.A1(net2210),
    .A2(_13828_),
    .B(_13964_),
    .C(_13649_),
    .Y(_13965_));
 BUFx16f_ASAP7_75t_R wire299 (.A(_06296_),
    .Y(net299));
 BUFx6f_ASAP7_75t_R load_slew298 (.A(\ex_block_i.alu_adder_result_ex_o[0] ),
    .Y(net298));
 NAND2x1_ASAP7_75t_R _19251_ (.A(net2378),
    .B(_00299_),
    .Y(_13968_));
 OA211x2_ASAP7_75t_R _19252_ (.A1(net2210),
    .A2(_13823_),
    .B(_13968_),
    .C(_00290_),
    .Y(_13969_));
 OR3x1_ASAP7_75t_R _19253_ (.A(_13626_),
    .B(_13965_),
    .C(_13969_),
    .Y(_13970_));
 BUFx6f_ASAP7_75t_R load_slew297 (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .Y(net297));
 NAND2x1_ASAP7_75t_R _19255_ (.A(net427),
    .B(_00317_),
    .Y(_13972_));
 OA211x2_ASAP7_75t_R _19256_ (.A1(net427),
    .A2(_13867_),
    .B(_13972_),
    .C(_13675_),
    .Y(_13973_));
 INVx1_ASAP7_75t_R _19257_ (.A(_00316_),
    .Y(_13974_));
 NAND2x1_ASAP7_75t_R _19258_ (.A(net427),
    .B(_00315_),
    .Y(_13975_));
 BUFx6f_ASAP7_75t_R load_slew296 (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .Y(net296));
 OA211x2_ASAP7_75t_R _19260_ (.A1(net427),
    .A2(_13974_),
    .B(_13975_),
    .C(net418),
    .Y(_13977_));
 OR3x1_ASAP7_75t_R _19261_ (.A(_00286_),
    .B(_13973_),
    .C(_13977_),
    .Y(_13978_));
 AND3x1_ASAP7_75t_R _19262_ (.A(net2300),
    .B(_13970_),
    .C(_13978_),
    .Y(_13979_));
 OR3x2_ASAP7_75t_R _19263_ (.A(net382),
    .B(_13959_),
    .C(_13979_),
    .Y(_13980_));
 AND2x4_ASAP7_75t_R _19264_ (.A(_13946_),
    .B(_13980_),
    .Y(_13981_));
 BUFx6f_ASAP7_75t_R load_slew295 (.A(net2194),
    .Y(net295));
 BUFx12f_ASAP7_75t_R wire294 (.A(_02537_),
    .Y(net294));
 BUFx6f_ASAP7_75t_R load_slew293 (.A(net174),
    .Y(net293));
 AOI22x1_ASAP7_75t_R _19268_ (.A1(_13775_),
    .A2(_00324_),
    .B1(_01452_),
    .B2(_13778_),
    .Y(_13985_));
 NAND2x2_ASAP7_75t_R _19269_ (.A(_00284_),
    .B(_13771_),
    .Y(_13986_));
 BUFx12f_ASAP7_75t_R wire292 (.A(_18555_),
    .Y(net292));
 OA211x2_ASAP7_75t_R _19271_ (.A1(_00284_),
    .A2(_13981_),
    .B(_13985_),
    .C(_13986_),
    .Y(_13988_));
 AO21x1_ASAP7_75t_R _19272_ (.A1(_13772_),
    .A2(_13886_),
    .B(_13988_),
    .Y(_13989_));
 BUFx12f_ASAP7_75t_R max_cap291 (.A(net292),
    .Y(net291));
 XNOR2x1_ASAP7_75t_R _19274_ (.B(_13893_),
    .Y(_13991_),
    .A(_13620_));
 AND2x2_ASAP7_75t_R _19275_ (.A(_13538_),
    .B(_13991_),
    .Y(_13992_));
 AO21x1_ASAP7_75t_R _19276_ (.A1(_13817_),
    .A2(_13989_),
    .B(_13992_),
    .Y(_16718_));
 OA21x2_ASAP7_75t_R _19277_ (.A1(_13788_),
    .A2(_13806_),
    .B(_13807_),
    .Y(_13993_));
 BUFx12f_ASAP7_75t_R max_cap290 (.A(_06981_),
    .Y(net290));
 BUFx6f_ASAP7_75t_R wire289 (.A(net176),
    .Y(net289));
 INVx1_ASAP7_75t_R _19280_ (.A(_01641_),
    .Y(_13996_));
 AO32x1_ASAP7_75t_R _19281_ (.A1(net319),
    .A2(_13802_),
    .A3(_13993_),
    .B1(_13996_),
    .B2(_13450_),
    .Y(_13997_));
 AND3x2_ASAP7_75t_R _19282_ (.A(_13810_),
    .B(_13946_),
    .C(_13980_),
    .Y(_13998_));
 OR2x2_ASAP7_75t_R _19283_ (.A(_13997_),
    .B(_13998_),
    .Y(_13999_));
 BUFx16f_ASAP7_75t_R wire288 (.A(_06987_),
    .Y(net288));
 INVx2_ASAP7_75t_R _19285_ (.A(_13999_),
    .Y(_18326_));
 BUFx16f_ASAP7_75t_R load_slew287 (.A(_09831_),
    .Y(net287));
 OR3x1_ASAP7_75t_R _19287_ (.A(_00324_),
    .B(_13538_),
    .C(_13815_),
    .Y(_14001_));
 OA21x2_ASAP7_75t_R _19288_ (.A1(_13817_),
    .A2(_18326_),
    .B(_14001_),
    .Y(_16719_));
 OA211x2_ASAP7_75t_R _19289_ (.A1(_13577_),
    .A2(_13607_),
    .B(_13538_),
    .C(_13618_),
    .Y(_14002_));
 BUFx16f_ASAP7_75t_R load_slew286 (.A(_09873_),
    .Y(net286));
 BUFx16f_ASAP7_75t_R wire285 (.A(net286),
    .Y(net285));
 BUFx16f_ASAP7_75t_R load_slew284 (.A(_09915_),
    .Y(net284));
 NAND2x2_ASAP7_75t_R _19293_ (.A(net385),
    .B(net379),
    .Y(_14005_));
 BUFx16f_ASAP7_75t_R wire283 (.A(net284),
    .Y(net283));
 BUFx16f_ASAP7_75t_R load_slew282 (.A(_09996_),
    .Y(net282));
 NAND2x2_ASAP7_75t_R _19296_ (.A(net423),
    .B(net316),
    .Y(_14008_));
 BUFx16f_ASAP7_75t_R wire281 (.A(net282),
    .Y(net281));
 BUFx16f_ASAP7_75t_R load_slew280 (.A(_10037_),
    .Y(net280));
 AND2x2_ASAP7_75t_R _19299_ (.A(net399),
    .B(_01697_),
    .Y(_14011_));
 AO21x1_ASAP7_75t_R _19300_ (.A1(net316),
    .A2(_00326_),
    .B(_14011_),
    .Y(_14012_));
 BUFx16f_ASAP7_75t_R load_slew279 (.A(net280),
    .Y(net279));
 OAI22x1_ASAP7_75t_R _19302_ (.A1(_00325_),
    .A2(net2293),
    .B1(_14012_),
    .B2(net421),
    .Y(_14014_));
 NAND2x2_ASAP7_75t_R _19303_ (.A(net320),
    .B(net379),
    .Y(_14015_));
 BUFx16f_ASAP7_75t_R load_slew278 (.A(_10078_),
    .Y(net278));
 BUFx16f_ASAP7_75t_R wire277 (.A(net278),
    .Y(net277));
 BUFx16f_ASAP7_75t_R load_slew276 (.A(_10162_),
    .Y(net276));
 INVx1_ASAP7_75t_R _19307_ (.A(_00329_),
    .Y(_14019_));
 NAND2x1_ASAP7_75t_R _19308_ (.A(net399),
    .B(_00327_),
    .Y(_14020_));
 OA211x2_ASAP7_75t_R _19309_ (.A1(net399),
    .A2(_14019_),
    .B(_14020_),
    .C(net421),
    .Y(_14021_));
 INVx1_ASAP7_75t_R _19310_ (.A(_00330_),
    .Y(_14022_));
 NAND2x1_ASAP7_75t_R _19311_ (.A(net399),
    .B(_00328_),
    .Y(_14023_));
 OA211x2_ASAP7_75t_R _19312_ (.A1(net399),
    .A2(_14022_),
    .B(_14023_),
    .C(net317),
    .Y(_14024_));
 OR3x1_ASAP7_75t_R _19313_ (.A(net312),
    .B(_14021_),
    .C(_14024_),
    .Y(_14025_));
 OA21x2_ASAP7_75t_R _19314_ (.A1(_14005_),
    .A2(_14014_),
    .B(_14025_),
    .Y(_14026_));
 INVx1_ASAP7_75t_R _19315_ (.A(_00345_),
    .Y(_14027_));
 BUFx16f_ASAP7_75t_R wire275 (.A(_10162_),
    .Y(net275));
 NAND2x1_ASAP7_75t_R _19317_ (.A(net404),
    .B(_00343_),
    .Y(_14029_));
 OA211x2_ASAP7_75t_R _19318_ (.A1(net404),
    .A2(_14027_),
    .B(_14029_),
    .C(net321),
    .Y(_14030_));
 BUFx16f_ASAP7_75t_R load_slew274 (.A(_10214_),
    .Y(net274));
 BUFx16f_ASAP7_75t_R wire273 (.A(net274),
    .Y(net273));
 INVx1_ASAP7_75t_R _19321_ (.A(_00341_),
    .Y(_14033_));
 BUFx16f_ASAP7_75t_R load_slew272 (.A(_10271_),
    .Y(net272));
 BUFx16f_ASAP7_75t_R load_slew271 (.A(net272),
    .Y(net271));
 NAND2x1_ASAP7_75t_R _19324_ (.A(net404),
    .B(_00339_),
    .Y(_14036_));
 BUFx16f_ASAP7_75t_R load_slew270 (.A(_10434_),
    .Y(net270));
 OA211x2_ASAP7_75t_R _19326_ (.A1(net404),
    .A2(_14033_),
    .B(_14036_),
    .C(net383),
    .Y(_14038_));
 OR3x1_ASAP7_75t_R _19327_ (.A(net317),
    .B(_14030_),
    .C(_14038_),
    .Y(_14039_));
 INVx1_ASAP7_75t_R _19328_ (.A(_00346_),
    .Y(_14040_));
 NAND2x1_ASAP7_75t_R _19329_ (.A(net404),
    .B(_00344_),
    .Y(_14041_));
 OA211x2_ASAP7_75t_R _19330_ (.A1(net404),
    .A2(_14040_),
    .B(_14041_),
    .C(net321),
    .Y(_14042_));
 INVx1_ASAP7_75t_R _19331_ (.A(_00342_),
    .Y(_14043_));
 NAND2x1_ASAP7_75t_R _19332_ (.A(net404),
    .B(_00340_),
    .Y(_14044_));
 OA211x2_ASAP7_75t_R _19333_ (.A1(net404),
    .A2(_14043_),
    .B(_14044_),
    .C(net383),
    .Y(_14045_));
 OR3x1_ASAP7_75t_R _19334_ (.A(net421),
    .B(_14042_),
    .C(_14045_),
    .Y(_14046_));
 BUFx16f_ASAP7_75t_R load_slew269 (.A(net270),
    .Y(net269));
 BUFx16f_ASAP7_75t_R load_slew268 (.A(_10596_),
    .Y(net268));
 NAND2x1_ASAP7_75t_R _19337_ (.A(net380),
    .B(_13626_),
    .Y(_14049_));
 AO21x1_ASAP7_75t_R _19338_ (.A1(_14039_),
    .A2(_14046_),
    .B(_14049_),
    .Y(_14050_));
 BUFx16f_ASAP7_75t_R load_slew267 (.A(net268),
    .Y(net267));
 INVx1_ASAP7_75t_R _19340_ (.A(_00333_),
    .Y(_14052_));
 BUFx16f_ASAP7_75t_R load_slew266 (.A(_10784_),
    .Y(net266));
 BUFx16f_ASAP7_75t_R load_slew265 (.A(net266),
    .Y(net265));
 NAND2x1_ASAP7_75t_R _19343_ (.A(net403),
    .B(_00331_),
    .Y(_14055_));
 BUFx16f_ASAP7_75t_R load_slew264 (.A(_10946_),
    .Y(net264));
 OA211x2_ASAP7_75t_R _19345_ (.A1(net403),
    .A2(_14052_),
    .B(_14055_),
    .C(net420),
    .Y(_14057_));
 BUFx16f_ASAP7_75t_R wire263 (.A(net264),
    .Y(net263));
 INVx1_ASAP7_75t_R _19347_ (.A(_00334_),
    .Y(_14059_));
 NAND2x1_ASAP7_75t_R _19348_ (.A(net403),
    .B(_00332_),
    .Y(_14060_));
 BUFx6f_ASAP7_75t_R load_slew262 (.A(net152),
    .Y(net262));
 OA211x2_ASAP7_75t_R _19350_ (.A1(net403),
    .A2(_14059_),
    .B(_14060_),
    .C(net317),
    .Y(_14062_));
 OR3x1_ASAP7_75t_R _19351_ (.A(net321),
    .B(_14057_),
    .C(_14062_),
    .Y(_14063_));
 BUFx6f_ASAP7_75t_R load_slew261 (.A(net160),
    .Y(net261));
 BUFx6f_ASAP7_75t_R load_slew260 (.A(_00785_),
    .Y(net260));
 INVx1_ASAP7_75t_R _19354_ (.A(_00337_),
    .Y(_14066_));
 NAND2x1_ASAP7_75t_R _19355_ (.A(net403),
    .B(_00335_),
    .Y(_14067_));
 OA211x2_ASAP7_75t_R _19356_ (.A1(net403),
    .A2(_14066_),
    .B(_14067_),
    .C(net420),
    .Y(_14068_));
 INVx1_ASAP7_75t_R _19357_ (.A(_00338_),
    .Y(_14069_));
 BUFx6f_ASAP7_75t_R wire259 (.A(net158),
    .Y(net259));
 BUFx6f_ASAP7_75t_R wire258 (.A(net162),
    .Y(net258));
 NAND2x1_ASAP7_75t_R _19360_ (.A(net403),
    .B(_00336_),
    .Y(_14072_));
 BUFx16f_ASAP7_75t_R max_cap257 (.A(_07825_),
    .Y(net257));
 OA211x2_ASAP7_75t_R _19362_ (.A1(net403),
    .A2(_14069_),
    .B(_14072_),
    .C(net317),
    .Y(_14074_));
 OR3x1_ASAP7_75t_R _19363_ (.A(net384),
    .B(_14068_),
    .C(_14074_),
    .Y(_14075_));
 AO21x1_ASAP7_75t_R _19364_ (.A1(_14063_),
    .A2(_14075_),
    .B(_13626_),
    .Y(_14076_));
 BUFx16f_ASAP7_75t_R max_cap256 (.A(_07866_),
    .Y(net256));
 INVx1_ASAP7_75t_R _19366_ (.A(_00354_),
    .Y(_14078_));
 NAND2x1_ASAP7_75t_R _19367_ (.A(net403),
    .B(_00352_),
    .Y(_14079_));
 BUFx16f_ASAP7_75t_R load_slew255 (.A(_09319_),
    .Y(net255));
 OA211x2_ASAP7_75t_R _19369_ (.A1(net403),
    .A2(_14078_),
    .B(_14079_),
    .C(net321),
    .Y(_14081_));
 INVx1_ASAP7_75t_R _19370_ (.A(_00350_),
    .Y(_14082_));
 NAND2x1_ASAP7_75t_R _19371_ (.A(net403),
    .B(_00348_),
    .Y(_14083_));
 BUFx16f_ASAP7_75t_R wire254 (.A(net255),
    .Y(net254));
 OA211x2_ASAP7_75t_R _19373_ (.A1(net403),
    .A2(_14082_),
    .B(_14083_),
    .C(net384),
    .Y(_14085_));
 OR3x1_ASAP7_75t_R _19374_ (.A(net420),
    .B(_14081_),
    .C(_14085_),
    .Y(_14086_));
 BUFx12f_ASAP7_75t_R max_cap253 (.A(_12481_),
    .Y(net253));
 BUFx12f_ASAP7_75t_R max_cap252 (.A(_07760_),
    .Y(net252));
 BUFx6f_ASAP7_75t_R max_cap251 (.A(_08026_),
    .Y(net251));
 INVx1_ASAP7_75t_R _19378_ (.A(_00353_),
    .Y(_14090_));
 NAND2x1_ASAP7_75t_R _19379_ (.A(net403),
    .B(_00351_),
    .Y(_14091_));
 OA211x2_ASAP7_75t_R _19380_ (.A1(net403),
    .A2(_14090_),
    .B(_14091_),
    .C(net321),
    .Y(_14092_));
 INVx1_ASAP7_75t_R _19381_ (.A(_00349_),
    .Y(_14093_));
 NAND2x1_ASAP7_75t_R _19382_ (.A(net403),
    .B(_00347_),
    .Y(_14094_));
 OA211x2_ASAP7_75t_R _19383_ (.A1(net403),
    .A2(_14093_),
    .B(_14094_),
    .C(net384),
    .Y(_14095_));
 OR3x1_ASAP7_75t_R _19384_ (.A(net317),
    .B(_14092_),
    .C(_14095_),
    .Y(_14096_));
 AO21x1_ASAP7_75t_R _19385_ (.A1(_14086_),
    .A2(_14096_),
    .B(net377),
    .Y(_14097_));
 AO21x1_ASAP7_75t_R _19386_ (.A1(_14076_),
    .A2(_14097_),
    .B(net380),
    .Y(_14098_));
 OA211x2_ASAP7_75t_R _19387_ (.A1(_13626_),
    .A2(_14026_),
    .B(_14050_),
    .C(_14098_),
    .Y(_14099_));
 BUFx16f_ASAP7_75t_R max_cap250 (.A(_08593_),
    .Y(net250));
 BUFx2_ASAP7_75t_R output249 (.A(net249),
    .Y(instr_req_o));
 BUFx2_ASAP7_75t_R output248 (.A(net248),
    .Y(instr_addr_o[9]));
 NAND2x2_ASAP7_75t_R _19391_ (.A(_13993_),
    .B(_13794_),
    .Y(_14103_));
 OAI22x1_ASAP7_75t_R _19392_ (.A1(_01629_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00199_),
    .Y(_14104_));
 AOI21x1_ASAP7_75t_R _19393_ (.A1(_13810_),
    .A2(_14099_),
    .B(_14104_),
    .Y(_18385_));
 BUFx2_ASAP7_75t_R output247 (.A(net247),
    .Y(instr_addr_o[8]));
 BUFx2_ASAP7_75t_R output246 (.A(net246),
    .Y(instr_addr_o[7]));
 NAND2x1_ASAP7_75t_R _19396_ (.A(net2257),
    .B(_00370_),
    .Y(_14107_));
 BUFx2_ASAP7_75t_R output245 (.A(net245),
    .Y(instr_addr_o[6]));
 NAND2x1_ASAP7_75t_R _19398_ (.A(net2278),
    .B(_00372_),
    .Y(_14109_));
 NAND2x1_ASAP7_75t_R _19399_ (.A(net2257),
    .B(_00369_),
    .Y(_14110_));
 NAND2x1_ASAP7_75t_R _19400_ (.A(net2278),
    .B(_00371_),
    .Y(_14111_));
 AO33x2_ASAP7_75t_R _19401_ (.A1(_13377_),
    .A2(_14107_),
    .A3(_14109_),
    .B1(_14110_),
    .B2(_14111_),
    .B3(_13357_),
    .Y(_14112_));
 BUFx2_ASAP7_75t_R output244 (.A(net244),
    .Y(instr_addr_o[5]));
 INVx1_ASAP7_75t_R _19403_ (.A(_00373_),
    .Y(_14114_));
 BUFx2_ASAP7_75t_R output243 (.A(net243),
    .Y(instr_addr_o[4]));
 NOR2x1_ASAP7_75t_R _19405_ (.A(net363),
    .B(_00375_),
    .Y(_14116_));
 AO21x1_ASAP7_75t_R _19406_ (.A1(net2333),
    .A2(_14114_),
    .B(_14116_),
    .Y(_14117_));
 INVx1_ASAP7_75t_R _19407_ (.A(_00376_),
    .Y(_14118_));
 NAND2x1_ASAP7_75t_R _19408_ (.A(net2257),
    .B(_00374_),
    .Y(_14119_));
 OA211x2_ASAP7_75t_R _19409_ (.A1(net2259),
    .A2(_14118_),
    .B(net322),
    .C(_14119_),
    .Y(_14120_));
 AO21x1_ASAP7_75t_R _19410_ (.A1(_13366_),
    .A2(_14117_),
    .B(_14120_),
    .Y(_14121_));
 OA21x2_ASAP7_75t_R _19411_ (.A1(_14112_),
    .A2(_14121_),
    .B(_13356_),
    .Y(_14122_));
 NAND2x1_ASAP7_75t_R _19412_ (.A(net374),
    .B(_00377_),
    .Y(_14123_));
 NAND2x1_ASAP7_75t_R _19413_ (.A(net325),
    .B(_00378_),
    .Y(_14124_));
 AND2x6_ASAP7_75t_R _19414_ (.A(net367),
    .B(net336),
    .Y(_14125_));
 AND2x4_ASAP7_75t_R _19415_ (.A(net326),
    .B(net336),
    .Y(_14126_));
 INVx1_ASAP7_75t_R _19416_ (.A(_00380_),
    .Y(_14127_));
 NAND2x1_ASAP7_75t_R _19417_ (.A(net374),
    .B(_00379_),
    .Y(_14128_));
 OA21x2_ASAP7_75t_R _19418_ (.A1(net374),
    .A2(_14127_),
    .B(_14128_),
    .Y(_14129_));
 AO32x1_ASAP7_75t_R _19419_ (.A1(_14123_),
    .A2(_14124_),
    .A3(_14125_),
    .B1(_14126_),
    .B2(_14129_),
    .Y(_14130_));
 BUFx2_ASAP7_75t_R output242 (.A(net242),
    .Y(instr_addr_o[3]));
 INVx1_ASAP7_75t_R _19421_ (.A(_00383_),
    .Y(_14132_));
 NAND2x1_ASAP7_75t_R _19422_ (.A(net2257),
    .B(_00381_),
    .Y(_14133_));
 OA21x2_ASAP7_75t_R _19423_ (.A1(net2259),
    .A2(_14132_),
    .B(_14133_),
    .Y(_14134_));
 INVx1_ASAP7_75t_R _19424_ (.A(_00384_),
    .Y(_14135_));
 NAND2x1_ASAP7_75t_R _19425_ (.A(net2257),
    .B(_00382_),
    .Y(_14136_));
 OA211x2_ASAP7_75t_R _19426_ (.A1(net2265),
    .A2(_14135_),
    .B(net322),
    .C(_14136_),
    .Y(_14137_));
 AO21x1_ASAP7_75t_R _19427_ (.A1(_13366_),
    .A2(_14134_),
    .B(_14137_),
    .Y(_14138_));
 OA21x2_ASAP7_75t_R _19428_ (.A1(_14130_),
    .A2(_14138_),
    .B(_13439_),
    .Y(_14139_));
 INVx1_ASAP7_75t_R _19429_ (.A(_00363_),
    .Y(_14140_));
 NAND2x1_ASAP7_75t_R _19430_ (.A(net2257),
    .B(_00361_),
    .Y(_14141_));
 OA21x2_ASAP7_75t_R _19431_ (.A1(net364),
    .A2(_14140_),
    .B(_14141_),
    .Y(_14142_));
 INVx1_ASAP7_75t_R _19432_ (.A(_00367_),
    .Y(_14143_));
 NAND2x1_ASAP7_75t_R _19433_ (.A(net2257),
    .B(_00365_),
    .Y(_14144_));
 OA21x2_ASAP7_75t_R _19434_ (.A1(net2265),
    .A2(_14143_),
    .B(_14144_),
    .Y(_14145_));
 INVx1_ASAP7_75t_R _19435_ (.A(_00368_),
    .Y(_14146_));
 NAND2x1_ASAP7_75t_R _19436_ (.A(net2257),
    .B(_00366_),
    .Y(_14147_));
 OA211x2_ASAP7_75t_R _19437_ (.A1(net364),
    .A2(_14146_),
    .B(net322),
    .C(_14147_),
    .Y(_14148_));
 AO221x1_ASAP7_75t_R _19438_ (.A1(_13357_),
    .A2(_14142_),
    .B1(_14145_),
    .B2(_13366_),
    .C(_14148_),
    .Y(_14149_));
 BUFx2_ASAP7_75t_R output241 (.A(net241),
    .Y(instr_addr_o[31]));
 INVx1_ASAP7_75t_R _19440_ (.A(_00364_),
    .Y(_14151_));
 NAND2x1_ASAP7_75t_R _19441_ (.A(net2257),
    .B(_00362_),
    .Y(_14152_));
 OA21x2_ASAP7_75t_R _19442_ (.A1(net2265),
    .A2(_14151_),
    .B(_14152_),
    .Y(_14153_));
 AO21x1_ASAP7_75t_R _19443_ (.A1(_13377_),
    .A2(_14153_),
    .B(net329),
    .Y(_14154_));
 AND2x2_ASAP7_75t_R _19444_ (.A(net2259),
    .B(_00357_),
    .Y(_14155_));
 AO21x1_ASAP7_75t_R _19445_ (.A1(_13359_),
    .A2(_00359_),
    .B(_14155_),
    .Y(_14156_));
 BUFx2_ASAP7_75t_R output240 (.A(net240),
    .Y(instr_addr_o[30]));
 AND2x2_ASAP7_75t_R _19447_ (.A(net2259),
    .B(_00358_),
    .Y(_14158_));
 AO21x1_ASAP7_75t_R _19448_ (.A1(_13359_),
    .A2(_00360_),
    .B(_14158_),
    .Y(_14159_));
 BUFx2_ASAP7_75t_R output239 (.A(net239),
    .Y(instr_addr_o[2]));
 AOI22x1_ASAP7_75t_R _19450_ (.A1(_13366_),
    .A2(_14156_),
    .B1(_14159_),
    .B2(net322),
    .Y(_14161_));
 INVx1_ASAP7_75t_R _19451_ (.A(_00356_),
    .Y(_14162_));
 NAND2x1_ASAP7_75t_R _19452_ (.A(net2259),
    .B(_01707_),
    .Y(_14163_));
 OA211x2_ASAP7_75t_R _19453_ (.A1(net2265),
    .A2(_14162_),
    .B(_14163_),
    .C(net325),
    .Y(_14164_));
 INVx1_ASAP7_75t_R _19454_ (.A(_00355_),
    .Y(_14165_));
 AND3x1_ASAP7_75t_R _19455_ (.A(net374),
    .B(net2260),
    .C(_14165_),
    .Y(_14166_));
 OA31x2_ASAP7_75t_R _19456_ (.A1(_13851_),
    .A2(_14164_),
    .A3(_14166_),
    .B1(net327),
    .Y(_14167_));
 OA221x2_ASAP7_75t_R _19457_ (.A1(_14149_),
    .A2(_14154_),
    .B1(_14161_),
    .B2(_13373_),
    .C(_14167_),
    .Y(_14168_));
 OR3x4_ASAP7_75t_R _19458_ (.A(_14122_),
    .B(_14139_),
    .C(_14168_),
    .Y(_14169_));
 BUFx2_ASAP7_75t_R output238 (.A(net238),
    .Y(instr_addr_o[29]));
 AND3x1_ASAP7_75t_R _19460_ (.A(_00385_),
    .B(_13505_),
    .C(_13891_),
    .Y(_14171_));
 BUFx2_ASAP7_75t_R output237 (.A(net237),
    .Y(instr_addr_o[28]));
 AND2x2_ASAP7_75t_R _19462_ (.A(_13807_),
    .B(_13473_),
    .Y(_14173_));
 OAI21x1_ASAP7_75t_R _19463_ (.A1(net2361),
    .A2(_13520_),
    .B(_14173_),
    .Y(_14174_));
 BUFx2_ASAP7_75t_R output236 (.A(net236),
    .Y(instr_addr_o[27]));
 INVx3_ASAP7_75t_R _19465_ (.A(_00187_),
    .Y(_14176_));
 AND3x2_ASAP7_75t_R _19466_ (.A(_13807_),
    .B(_13481_),
    .C(_13513_),
    .Y(_14177_));
 AND3x1_ASAP7_75t_R _19467_ (.A(_14176_),
    .B(_13520_),
    .C(_14177_),
    .Y(_14178_));
 OA33x2_ASAP7_75t_R _19468_ (.A1(_13450_),
    .A2(_13473_),
    .A3(_14169_),
    .B1(_14171_),
    .B2(_14174_),
    .B3(_14178_),
    .Y(_14179_));
 CKINVDCx12_ASAP7_75t_R _19469_ (.A(_14179_),
    .Y(_14180_));
 BUFx2_ASAP7_75t_R output235 (.A(net235),
    .Y(instr_addr_o[26]));
 BUFx2_ASAP7_75t_R output234 (.A(net234),
    .Y(instr_addr_o[25]));
 INVx4_ASAP7_75t_R _19472_ (.A(_00191_),
    .Y(_14182_));
 AND2x2_ASAP7_75t_R _19473_ (.A(_13520_),
    .B(_14177_),
    .Y(_14183_));
 NAND2x2_ASAP7_75t_R _19474_ (.A(net372),
    .B(_13359_),
    .Y(_14184_));
 AND2x2_ASAP7_75t_R _19475_ (.A(net345),
    .B(_01706_),
    .Y(_14185_));
 AO21x1_ASAP7_75t_R _19476_ (.A1(net326),
    .A2(_00387_),
    .B(_14185_),
    .Y(_14186_));
 OAI22x1_ASAP7_75t_R _19477_ (.A1(_00386_),
    .A2(net311),
    .B1(_14186_),
    .B2(net376),
    .Y(_14187_));
 AND2x2_ASAP7_75t_R _19478_ (.A(net344),
    .B(_00388_),
    .Y(_14188_));
 AO21x1_ASAP7_75t_R _19479_ (.A1(net326),
    .A2(_00390_),
    .B(_14188_),
    .Y(_14189_));
 AND2x2_ASAP7_75t_R _19480_ (.A(net344),
    .B(_00389_),
    .Y(_14190_));
 AO21x1_ASAP7_75t_R _19481_ (.A1(net326),
    .A2(_00391_),
    .B(_14190_),
    .Y(_14191_));
 AOI22x1_ASAP7_75t_R _19482_ (.A1(_13366_),
    .A2(_14189_),
    .B1(_14191_),
    .B2(_13402_),
    .Y(_14192_));
 OA21x2_ASAP7_75t_R _19483_ (.A1(_13350_),
    .A2(_14187_),
    .B(_14192_),
    .Y(_14193_));
 INVx1_ASAP7_75t_R _19484_ (.A(_00403_),
    .Y(_14194_));
 NAND2x1_ASAP7_75t_R _19485_ (.A(net341),
    .B(_00401_),
    .Y(_14195_));
 OA21x2_ASAP7_75t_R _19486_ (.A1(net341),
    .A2(_14194_),
    .B(_14195_),
    .Y(_14196_));
 INVx1_ASAP7_75t_R _19487_ (.A(_00402_),
    .Y(_14197_));
 NAND2x1_ASAP7_75t_R _19488_ (.A(net341),
    .B(_00400_),
    .Y(_14198_));
 OA211x2_ASAP7_75t_R _19489_ (.A1(net341),
    .A2(_14197_),
    .B(_13357_),
    .C(_14198_),
    .Y(_14199_));
 INVx1_ASAP7_75t_R _19490_ (.A(_00407_),
    .Y(_14200_));
 NAND2x1_ASAP7_75t_R _19491_ (.A(net341),
    .B(_00405_),
    .Y(_14201_));
 OA211x2_ASAP7_75t_R _19492_ (.A1(net341),
    .A2(_14200_),
    .B(_13402_),
    .C(_14201_),
    .Y(_14202_));
 AOI211x1_ASAP7_75t_R _19493_ (.A1(_13377_),
    .A2(_14196_),
    .B(_14199_),
    .C(_14202_),
    .Y(_14203_));
 NAND2x1_ASAP7_75t_R _19494_ (.A(net376),
    .B(_13350_),
    .Y(_14204_));
 AND2x2_ASAP7_75t_R _19495_ (.A(net341),
    .B(_00404_),
    .Y(_14205_));
 AO21x1_ASAP7_75t_R _19496_ (.A1(net326),
    .A2(_00406_),
    .B(_14205_),
    .Y(_14206_));
 OA21x2_ASAP7_75t_R _19497_ (.A1(_14204_),
    .A2(_14206_),
    .B(_13356_),
    .Y(_14207_));
 INVx1_ASAP7_75t_R _19498_ (.A(_00395_),
    .Y(_14208_));
 NAND2x1_ASAP7_75t_R _19499_ (.A(net368),
    .B(_00393_),
    .Y(_14209_));
 OA21x2_ASAP7_75t_R _19500_ (.A1(net368),
    .A2(_14208_),
    .B(_14209_),
    .Y(_14210_));
 INVx1_ASAP7_75t_R _19501_ (.A(_00399_),
    .Y(_14211_));
 NAND2x1_ASAP7_75t_R _19502_ (.A(net368),
    .B(_00397_),
    .Y(_14212_));
 OA211x2_ASAP7_75t_R _19503_ (.A1(net368),
    .A2(_14211_),
    .B(_13402_),
    .C(_14212_),
    .Y(_14213_));
 INVx1_ASAP7_75t_R _19504_ (.A(_00394_),
    .Y(_14214_));
 NAND2x1_ASAP7_75t_R _19505_ (.A(net368),
    .B(_00392_),
    .Y(_14215_));
 OA211x2_ASAP7_75t_R _19506_ (.A1(net368),
    .A2(_14214_),
    .B(_13357_),
    .C(_14215_),
    .Y(_14216_));
 AOI211x1_ASAP7_75t_R _19507_ (.A1(_13377_),
    .A2(_14210_),
    .B(_14213_),
    .C(_14216_),
    .Y(_14217_));
 AND2x2_ASAP7_75t_R _19508_ (.A(net344),
    .B(_00396_),
    .Y(_14218_));
 AO21x1_ASAP7_75t_R _19509_ (.A1(net326),
    .A2(_00398_),
    .B(_14218_),
    .Y(_14219_));
 OA21x2_ASAP7_75t_R _19510_ (.A1(_14204_),
    .A2(_14219_),
    .B(_13375_),
    .Y(_14220_));
 AOI22x1_ASAP7_75t_R _19511_ (.A1(_14203_),
    .A2(_14207_),
    .B1(_14217_),
    .B2(_14220_),
    .Y(_14221_));
 AND2x2_ASAP7_75t_R _19512_ (.A(net368),
    .B(_00408_),
    .Y(_14222_));
 AO21x1_ASAP7_75t_R _19513_ (.A1(net326),
    .A2(_00410_),
    .B(_14222_),
    .Y(_14223_));
 AND2x2_ASAP7_75t_R _19514_ (.A(net344),
    .B(_00412_),
    .Y(_14224_));
 AO21x1_ASAP7_75t_R _19515_ (.A1(net326),
    .A2(_00414_),
    .B(_14224_),
    .Y(_14225_));
 AO22x1_ASAP7_75t_R _19516_ (.A1(_13357_),
    .A2(_14223_),
    .B1(_14225_),
    .B2(_13366_),
    .Y(_14226_));
 AND2x2_ASAP7_75t_R _19517_ (.A(net344),
    .B(_00413_),
    .Y(_14227_));
 AO21x1_ASAP7_75t_R _19518_ (.A1(net326),
    .A2(_00415_),
    .B(_14227_),
    .Y(_14228_));
 AND2x2_ASAP7_75t_R _19519_ (.A(net368),
    .B(_00409_),
    .Y(_14229_));
 AO21x1_ASAP7_75t_R _19520_ (.A1(net326),
    .A2(_00411_),
    .B(_14229_),
    .Y(_14230_));
 AO22x1_ASAP7_75t_R _19521_ (.A1(_13402_),
    .A2(_14228_),
    .B1(_14230_),
    .B2(_13377_),
    .Y(_14231_));
 OAI21x1_ASAP7_75t_R _19522_ (.A1(_14226_),
    .A2(_14231_),
    .B(_13439_),
    .Y(_14232_));
 OA211x2_ASAP7_75t_R _19523_ (.A1(_13410_),
    .A2(_14193_),
    .B(_14221_),
    .C(_14232_),
    .Y(_14233_));
 BUFx2_ASAP7_75t_R output233 (.A(net233),
    .Y(instr_addr_o[24]));
 BUFx2_ASAP7_75t_R output232 (.A(net232),
    .Y(instr_addr_o[23]));
 AND2x2_ASAP7_75t_R _19526_ (.A(_13373_),
    .B(_13473_),
    .Y(_14236_));
 AND2x2_ASAP7_75t_R _19527_ (.A(_13495_),
    .B(_14236_),
    .Y(_14237_));
 AOI221x1_ASAP7_75t_R _19528_ (.A1(_14182_),
    .A2(_14183_),
    .B1(_14233_),
    .B2(_13474_),
    .C(_14237_),
    .Y(_14238_));
 CKINVDCx12_ASAP7_75t_R _19529_ (.A(_14238_),
    .Y(_14239_));
 BUFx2_ASAP7_75t_R output231 (.A(net231),
    .Y(instr_addr_o[22]));
 BUFx2_ASAP7_75t_R output230 (.A(net230),
    .Y(instr_addr_o[21]));
 BUFx2_ASAP7_75t_R output229 (.A(net229),
    .Y(instr_addr_o[20]));
 INVx1_ASAP7_75t_R _19533_ (.A(_00428_),
    .Y(_14241_));
 NAND2x1_ASAP7_75t_R _19534_ (.A(net361),
    .B(_00426_),
    .Y(_14242_));
 OA211x2_ASAP7_75t_R _19535_ (.A1(net361),
    .A2(_14241_),
    .B(_13366_),
    .C(_14242_),
    .Y(_14243_));
 AND2x2_ASAP7_75t_R _19536_ (.A(net361),
    .B(_00422_),
    .Y(_14244_));
 AO21x1_ASAP7_75t_R _19537_ (.A1(_13359_),
    .A2(_00424_),
    .B(_14244_),
    .Y(_14245_));
 OR2x2_ASAP7_75t_R _19538_ (.A(net361),
    .B(_00425_),
    .Y(_14246_));
 OA211x2_ASAP7_75t_R _19539_ (.A1(_13359_),
    .A2(_00423_),
    .B(_14246_),
    .C(net324),
    .Y(_14247_));
 AOI211x1_ASAP7_75t_R _19540_ (.A1(net373),
    .A2(_14245_),
    .B(_14247_),
    .C(_13350_),
    .Y(_14248_));
 INVx1_ASAP7_75t_R _19541_ (.A(_00429_),
    .Y(_14249_));
 NAND2x1_ASAP7_75t_R _19542_ (.A(net361),
    .B(_00427_),
    .Y(_14250_));
 OA211x2_ASAP7_75t_R _19543_ (.A1(net361),
    .A2(_14249_),
    .B(net322),
    .C(_14250_),
    .Y(_14251_));
 OR4x2_ASAP7_75t_R _19544_ (.A(net329),
    .B(_14243_),
    .C(_14248_),
    .D(_14251_),
    .Y(_14252_));
 AND2x2_ASAP7_75t_R _19545_ (.A(net2267),
    .B(_00418_),
    .Y(_14253_));
 AO21x1_ASAP7_75t_R _19546_ (.A1(net2260),
    .A2(_00420_),
    .B(_14253_),
    .Y(_14254_));
 AND2x2_ASAP7_75t_R _19547_ (.A(net2258),
    .B(_00419_),
    .Y(_14255_));
 AO21x1_ASAP7_75t_R _19548_ (.A1(net2260),
    .A2(_00421_),
    .B(_14255_),
    .Y(_14256_));
 AOI22x1_ASAP7_75t_R _19549_ (.A1(_13366_),
    .A2(_14254_),
    .B1(_14256_),
    .B2(net322),
    .Y(_14257_));
 INVx1_ASAP7_75t_R _19550_ (.A(_00416_),
    .Y(_14258_));
 INVx1_ASAP7_75t_R _19551_ (.A(_00417_),
    .Y(_14259_));
 NAND2x1_ASAP7_75t_R _19552_ (.A(net357),
    .B(_01705_),
    .Y(_14260_));
 OA21x2_ASAP7_75t_R _19553_ (.A1(net357),
    .A2(_14259_),
    .B(_14260_),
    .Y(_14261_));
 AO221x1_ASAP7_75t_R _19554_ (.A1(_14258_),
    .A2(net2227),
    .B1(_14261_),
    .B2(net324),
    .C(_13851_),
    .Y(_14262_));
 OA211x2_ASAP7_75t_R _19555_ (.A1(_13373_),
    .A2(_14257_),
    .B(_14262_),
    .C(net327),
    .Y(_14263_));
 INVx1_ASAP7_75t_R _19556_ (.A(_00436_),
    .Y(_14264_));
 NAND2x1_ASAP7_75t_R _19557_ (.A(net2258),
    .B(_00434_),
    .Y(_14265_));
 OA211x2_ASAP7_75t_R _19558_ (.A1(net2268),
    .A2(_14264_),
    .B(_14265_),
    .C(_13350_),
    .Y(_14266_));
 INVx1_ASAP7_75t_R _19559_ (.A(_00432_),
    .Y(_14267_));
 NAND2x1_ASAP7_75t_R _19560_ (.A(net2258),
    .B(_00430_),
    .Y(_14268_));
 OA211x2_ASAP7_75t_R _19561_ (.A1(net2267),
    .A2(_14267_),
    .B(_14268_),
    .C(net334),
    .Y(_14269_));
 OR3x1_ASAP7_75t_R _19562_ (.A(net324),
    .B(_14266_),
    .C(_14269_),
    .Y(_14270_));
 AND2x2_ASAP7_75t_R _19563_ (.A(net2258),
    .B(_00435_),
    .Y(_14271_));
 AO21x1_ASAP7_75t_R _19564_ (.A1(net2260),
    .A2(_00437_),
    .B(_14271_),
    .Y(_14272_));
 AND2x2_ASAP7_75t_R _19565_ (.A(net2258),
    .B(_00431_),
    .Y(_14273_));
 AO21x1_ASAP7_75t_R _19566_ (.A1(net2260),
    .A2(_00433_),
    .B(_14273_),
    .Y(_14274_));
 NAND2x2_ASAP7_75t_R _19567_ (.A(net329),
    .B(_13355_),
    .Y(_14275_));
 AOI221x1_ASAP7_75t_R _19568_ (.A1(net322),
    .A2(_14272_),
    .B1(_14274_),
    .B2(_13377_),
    .C(_14275_),
    .Y(_14276_));
 INVx1_ASAP7_75t_R _19569_ (.A(_00439_),
    .Y(_14277_));
 NAND2x1_ASAP7_75t_R _19570_ (.A(net372),
    .B(_00438_),
    .Y(_14278_));
 OA211x2_ASAP7_75t_R _19571_ (.A1(net372),
    .A2(_14277_),
    .B(_14125_),
    .C(_14278_),
    .Y(_14279_));
 INVx1_ASAP7_75t_R _19572_ (.A(_00440_),
    .Y(_14280_));
 NAND2x1_ASAP7_75t_R _19573_ (.A(net324),
    .B(_00441_),
    .Y(_14281_));
 OA211x2_ASAP7_75t_R _19574_ (.A1(net324),
    .A2(_14280_),
    .B(net2222),
    .C(_14281_),
    .Y(_14282_));
 INVx1_ASAP7_75t_R _19575_ (.A(_00444_),
    .Y(_14283_));
 NAND2x1_ASAP7_75t_R _19576_ (.A(net2258),
    .B(_00442_),
    .Y(_14284_));
 OA211x2_ASAP7_75t_R _19577_ (.A1(net2267),
    .A2(_14283_),
    .B(_13366_),
    .C(_14284_),
    .Y(_14285_));
 INVx1_ASAP7_75t_R _19578_ (.A(_00445_),
    .Y(_14286_));
 NAND2x1_ASAP7_75t_R _19579_ (.A(net2258),
    .B(_00443_),
    .Y(_14287_));
 OA211x2_ASAP7_75t_R _19580_ (.A1(net2267),
    .A2(_14286_),
    .B(net322),
    .C(_14287_),
    .Y(_14288_));
 OR4x1_ASAP7_75t_R _19581_ (.A(_14279_),
    .B(_14282_),
    .C(_14285_),
    .D(_14288_),
    .Y(_14289_));
 AO222x2_ASAP7_75t_R _19582_ (.A1(_14252_),
    .A2(_14263_),
    .B1(_14270_),
    .B2(_14276_),
    .C1(_14289_),
    .C2(_13439_),
    .Y(_14290_));
 BUFx2_ASAP7_75t_R output228 (.A(net228),
    .Y(instr_addr_o[19]));
 BUFx2_ASAP7_75t_R output227 (.A(net227),
    .Y(instr_addr_o[18]));
 INVx3_ASAP7_75t_R _19585_ (.A(_00194_),
    .Y(_14293_));
 AND3x4_ASAP7_75t_R _19586_ (.A(_14293_),
    .B(_13520_),
    .C(_14177_),
    .Y(_14294_));
 AND3x1_ASAP7_75t_R _19587_ (.A(_13355_),
    .B(_13521_),
    .C(_13495_),
    .Y(_14295_));
 AOI211x1_ASAP7_75t_R _19588_ (.A1(_13474_),
    .A2(net2218),
    .B(_14294_),
    .C(_14295_),
    .Y(_14296_));
 CKINVDCx10_ASAP7_75t_R _19589_ (.A(net302),
    .Y(_14297_));
 BUFx2_ASAP7_75t_R output226 (.A(net226),
    .Y(instr_addr_o[17]));
 BUFx2_ASAP7_75t_R output225 (.A(net225),
    .Y(instr_addr_o[16]));
 BUFx2_ASAP7_75t_R output224 (.A(net224),
    .Y(instr_addr_o[15]));
 BUFx2_ASAP7_75t_R output223 (.A(net223),
    .Y(instr_addr_o[14]));
 INVx1_ASAP7_75t_R _19594_ (.A(_02054_),
    .Y(\cs_registers_i.mhpmcounter[2][44] ));
 INVx1_ASAP7_75t_R _19595_ (.A(_02160_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[44] ));
 BUFx2_ASAP7_75t_R output222 (.A(net222),
    .Y(instr_addr_o[13]));
 INVx1_ASAP7_75t_R _19597_ (.A(_00463_),
    .Y(_14301_));
 NAND2x1_ASAP7_75t_R _19598_ (.A(net362),
    .B(_00461_),
    .Y(_14302_));
 OA211x2_ASAP7_75t_R _19599_ (.A1(net362),
    .A2(_14301_),
    .B(_13377_),
    .C(_14302_),
    .Y(_14303_));
 BUFx2_ASAP7_75t_R output221 (.A(net221),
    .Y(instr_addr_o[12]));
 INVx1_ASAP7_75t_R _19601_ (.A(_00467_),
    .Y(_14305_));
 NAND2x1_ASAP7_75t_R _19602_ (.A(net362),
    .B(_00465_),
    .Y(_14306_));
 OA211x2_ASAP7_75t_R _19603_ (.A1(net362),
    .A2(_14305_),
    .B(net322),
    .C(_14306_),
    .Y(_14307_));
 BUFx2_ASAP7_75t_R output220 (.A(net220),
    .Y(instr_addr_o[11]));
 INVx1_ASAP7_75t_R _19605_ (.A(_00466_),
    .Y(_14309_));
 NAND2x1_ASAP7_75t_R _19606_ (.A(net362),
    .B(_00464_),
    .Y(_14310_));
 OA211x2_ASAP7_75t_R _19607_ (.A1(net362),
    .A2(_14309_),
    .B(_13366_),
    .C(_14310_),
    .Y(_14311_));
 INVx1_ASAP7_75t_R _19608_ (.A(_00462_),
    .Y(_14312_));
 NAND2x1_ASAP7_75t_R _19609_ (.A(net362),
    .B(_00460_),
    .Y(_14313_));
 OA211x2_ASAP7_75t_R _19610_ (.A1(net362),
    .A2(_14312_),
    .B(_13357_),
    .C(_14313_),
    .Y(_14314_));
 OR4x1_ASAP7_75t_R _19611_ (.A(_14303_),
    .B(_14307_),
    .C(_14311_),
    .D(_14314_),
    .Y(_14315_));
 INVx1_ASAP7_75t_R _19612_ (.A(_00471_),
    .Y(_14316_));
 NAND2x1_ASAP7_75t_R _19613_ (.A(net361),
    .B(_00469_),
    .Y(_14317_));
 OA211x2_ASAP7_75t_R _19614_ (.A1(net361),
    .A2(_14316_),
    .B(_13377_),
    .C(_14317_),
    .Y(_14318_));
 INVx1_ASAP7_75t_R _19615_ (.A(_00475_),
    .Y(_14319_));
 NAND2x1_ASAP7_75t_R _19616_ (.A(net361),
    .B(_00473_),
    .Y(_14320_));
 OA211x2_ASAP7_75t_R _19617_ (.A1(net361),
    .A2(_14319_),
    .B(net322),
    .C(_14320_),
    .Y(_14321_));
 INVx1_ASAP7_75t_R _19618_ (.A(_00470_),
    .Y(_14322_));
 NAND2x1_ASAP7_75t_R _19619_ (.A(net361),
    .B(_00468_),
    .Y(_14323_));
 OA211x2_ASAP7_75t_R _19620_ (.A1(net361),
    .A2(_14322_),
    .B(_13357_),
    .C(_14323_),
    .Y(_14324_));
 INVx1_ASAP7_75t_R _19621_ (.A(_00474_),
    .Y(_14325_));
 NAND2x1_ASAP7_75t_R _19622_ (.A(net361),
    .B(_00472_),
    .Y(_14326_));
 OA211x2_ASAP7_75t_R _19623_ (.A1(net361),
    .A2(_14325_),
    .B(_13366_),
    .C(_14326_),
    .Y(_14327_));
 OR4x1_ASAP7_75t_R _19624_ (.A(_14318_),
    .B(_14321_),
    .C(_14324_),
    .D(_14327_),
    .Y(_14328_));
 BUFx2_ASAP7_75t_R output219 (.A(net219),
    .Y(instr_addr_o[10]));
 INVx1_ASAP7_75t_R _19626_ (.A(_00458_),
    .Y(_14330_));
 NAND2x1_ASAP7_75t_R _19627_ (.A(net361),
    .B(_00456_),
    .Y(_14331_));
 OA21x2_ASAP7_75t_R _19628_ (.A1(net361),
    .A2(_14330_),
    .B(_14331_),
    .Y(_14332_));
 INVx1_ASAP7_75t_R _19629_ (.A(_00454_),
    .Y(_14333_));
 NAND2x1_ASAP7_75t_R _19630_ (.A(net361),
    .B(_00452_),
    .Y(_14334_));
 OA211x2_ASAP7_75t_R _19631_ (.A1(net361),
    .A2(_14333_),
    .B(_13357_),
    .C(_14334_),
    .Y(_14335_));
 AO21x1_ASAP7_75t_R _19632_ (.A1(_13366_),
    .A2(_14332_),
    .B(_14335_),
    .Y(_14336_));
 INVx1_ASAP7_75t_R _19633_ (.A(_00459_),
    .Y(_14337_));
 NAND2x1_ASAP7_75t_R _19634_ (.A(net361),
    .B(_00457_),
    .Y(_14338_));
 OA211x2_ASAP7_75t_R _19635_ (.A1(net361),
    .A2(_14337_),
    .B(net322),
    .C(_14338_),
    .Y(_14339_));
 INVx1_ASAP7_75t_R _19636_ (.A(_00455_),
    .Y(_14340_));
 NAND2x1_ASAP7_75t_R _19637_ (.A(net361),
    .B(_00453_),
    .Y(_14341_));
 OA211x2_ASAP7_75t_R _19638_ (.A1(net361),
    .A2(_14340_),
    .B(_13377_),
    .C(_14341_),
    .Y(_14342_));
 OR4x1_ASAP7_75t_R _19639_ (.A(net329),
    .B(_14336_),
    .C(_14339_),
    .D(_14342_),
    .Y(_14343_));
 AND2x2_ASAP7_75t_R _19640_ (.A(net362),
    .B(_00448_),
    .Y(_14344_));
 AO21x1_ASAP7_75t_R _19641_ (.A1(net2260),
    .A2(_00450_),
    .B(_14344_),
    .Y(_14345_));
 AND2x2_ASAP7_75t_R _19642_ (.A(net362),
    .B(_00449_),
    .Y(_14346_));
 AO21x1_ASAP7_75t_R _19643_ (.A1(net2260),
    .A2(_00451_),
    .B(_14346_),
    .Y(_14347_));
 AOI22x1_ASAP7_75t_R _19644_ (.A1(_13366_),
    .A2(_14345_),
    .B1(_14347_),
    .B2(net322),
    .Y(_14348_));
 INVx1_ASAP7_75t_R _19645_ (.A(_00446_),
    .Y(_14349_));
 INVx1_ASAP7_75t_R _19646_ (.A(_00447_),
    .Y(_14350_));
 NAND2x1_ASAP7_75t_R _19647_ (.A(net362),
    .B(_01704_),
    .Y(_14351_));
 OA21x2_ASAP7_75t_R _19648_ (.A1(net362),
    .A2(_14350_),
    .B(_14351_),
    .Y(_14352_));
 AO221x1_ASAP7_75t_R _19649_ (.A1(_14349_),
    .A2(net2229),
    .B1(_14352_),
    .B2(net324),
    .C(_13851_),
    .Y(_14353_));
 OA211x2_ASAP7_75t_R _19650_ (.A1(_13373_),
    .A2(_14348_),
    .B(_14353_),
    .C(net327),
    .Y(_14354_));
 AO222x2_ASAP7_75t_R _19651_ (.A1(_13356_),
    .A2(_14315_),
    .B1(_14328_),
    .B2(_13439_),
    .C1(_14343_),
    .C2(_14354_),
    .Y(_14355_));
 OA21x2_ASAP7_75t_R _19652_ (.A1(_13450_),
    .A2(_13473_),
    .B(_13481_),
    .Y(_14356_));
 OA211x2_ASAP7_75t_R _19653_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14356_),
    .C(_13528_),
    .Y(_14357_));
 AO21x2_ASAP7_75t_R _19654_ (.A1(_13474_),
    .A2(_14355_),
    .B(_14357_),
    .Y(_14358_));
 INVx13_ASAP7_75t_R _19655_ (.A(_14358_),
    .Y(_14359_));
 BUFx2_ASAP7_75t_R output218 (.A(net218),
    .Y(data_we_o));
 BUFx2_ASAP7_75t_R output217 (.A(net217),
    .Y(data_wdata_o[9]));
 BUFx2_ASAP7_75t_R output216 (.A(net216),
    .Y(data_wdata_o[8]));
 CKINVDCx5p33_ASAP7_75t_R _19659_ (.A(_00283_),
    .Y(_14362_));
 OA211x2_ASAP7_75t_R _19660_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14362_),
    .C(_13481_),
    .Y(_14363_));
 BUFx2_ASAP7_75t_R output215 (.A(net215),
    .Y(data_wdata_o[7]));
 BUFx2_ASAP7_75t_R output214 (.A(net214),
    .Y(data_wdata_o[6]));
 INVx1_ASAP7_75t_R _19663_ (.A(_00488_),
    .Y(_14366_));
 NAND2x1_ASAP7_75t_R _19664_ (.A(net362),
    .B(_00486_),
    .Y(_14367_));
 OA21x2_ASAP7_75t_R _19665_ (.A1(net362),
    .A2(_14366_),
    .B(_14367_),
    .Y(_14368_));
 INVx1_ASAP7_75t_R _19666_ (.A(_00484_),
    .Y(_14369_));
 NAND2x1_ASAP7_75t_R _19667_ (.A(net362),
    .B(_00482_),
    .Y(_14370_));
 OA21x2_ASAP7_75t_R _19668_ (.A1(net362),
    .A2(_14369_),
    .B(_14370_),
    .Y(_14371_));
 AO221x1_ASAP7_75t_R _19669_ (.A1(_13366_),
    .A2(_14368_),
    .B1(_14371_),
    .B2(_13357_),
    .C(net329),
    .Y(_14372_));
 INVx1_ASAP7_75t_R _19670_ (.A(_00489_),
    .Y(_14373_));
 NAND2x1_ASAP7_75t_R _19671_ (.A(net334),
    .B(_00485_),
    .Y(_14374_));
 OA211x2_ASAP7_75t_R _19672_ (.A1(net334),
    .A2(_14373_),
    .B(_14374_),
    .C(net2260),
    .Y(_14375_));
 INVx1_ASAP7_75t_R _19673_ (.A(_00487_),
    .Y(_14376_));
 NAND2x1_ASAP7_75t_R _19674_ (.A(net334),
    .B(_00483_),
    .Y(_14377_));
 OA211x2_ASAP7_75t_R _19675_ (.A1(net334),
    .A2(_14376_),
    .B(_14377_),
    .C(net362),
    .Y(_14378_));
 OA21x2_ASAP7_75t_R _19676_ (.A1(_14375_),
    .A2(_14378_),
    .B(net325),
    .Y(_14379_));
 INVx1_ASAP7_75t_R _19677_ (.A(_00480_),
    .Y(_14380_));
 NAND2x1_ASAP7_75t_R _19678_ (.A(net362),
    .B(_00478_),
    .Y(_14381_));
 OA211x2_ASAP7_75t_R _19679_ (.A1(net362),
    .A2(_14380_),
    .B(_14381_),
    .C(net373),
    .Y(_14382_));
 NAND2x2_ASAP7_75t_R _19680_ (.A(_13350_),
    .B(net329),
    .Y(_14383_));
 INVx1_ASAP7_75t_R _19681_ (.A(_00481_),
    .Y(_14384_));
 NAND2x1_ASAP7_75t_R _19682_ (.A(net362),
    .B(_00479_),
    .Y(_14385_));
 OA211x2_ASAP7_75t_R _19683_ (.A1(net362),
    .A2(_14384_),
    .B(_14385_),
    .C(net325),
    .Y(_14386_));
 OR3x1_ASAP7_75t_R _19684_ (.A(_14382_),
    .B(_14383_),
    .C(_14386_),
    .Y(_14387_));
 INVx1_ASAP7_75t_R _19685_ (.A(_00476_),
    .Y(_14388_));
 AND3x1_ASAP7_75t_R _19686_ (.A(net373),
    .B(net2260),
    .C(_14388_),
    .Y(_14389_));
 INVx1_ASAP7_75t_R _19687_ (.A(_00477_),
    .Y(_14390_));
 NAND2x1_ASAP7_75t_R _19688_ (.A(net362),
    .B(_01703_),
    .Y(_14391_));
 OA211x2_ASAP7_75t_R _19689_ (.A1(net362),
    .A2(_14390_),
    .B(_14391_),
    .C(net324),
    .Y(_14392_));
 OA31x2_ASAP7_75t_R _19690_ (.A1(_13851_),
    .A2(_14389_),
    .A3(_14392_),
    .B1(net327),
    .Y(_14393_));
 OA211x2_ASAP7_75t_R _19691_ (.A1(_14372_),
    .A2(_14379_),
    .B(_14387_),
    .C(_14393_),
    .Y(_14394_));
 INVx1_ASAP7_75t_R _19692_ (.A(_00496_),
    .Y(_14395_));
 NAND2x1_ASAP7_75t_R _19693_ (.A(net2266),
    .B(_00494_),
    .Y(_14396_));
 OA211x2_ASAP7_75t_R _19694_ (.A1(net2266),
    .A2(_14395_),
    .B(_14396_),
    .C(net373),
    .Y(_14397_));
 INVx1_ASAP7_75t_R _19695_ (.A(_00497_),
    .Y(_14398_));
 NAND2x1_ASAP7_75t_R _19696_ (.A(net2266),
    .B(_00495_),
    .Y(_14399_));
 OA211x2_ASAP7_75t_R _19697_ (.A1(net2266),
    .A2(_14398_),
    .B(_14399_),
    .C(net325),
    .Y(_14400_));
 OR3x1_ASAP7_75t_R _19698_ (.A(net334),
    .B(_14397_),
    .C(_14400_),
    .Y(_14401_));
 AND2x2_ASAP7_75t_R _19699_ (.A(net2266),
    .B(_00491_),
    .Y(_14402_));
 AO21x1_ASAP7_75t_R _19700_ (.A1(_13359_),
    .A2(_00493_),
    .B(_14402_),
    .Y(_14403_));
 AND2x2_ASAP7_75t_R _19701_ (.A(net2266),
    .B(_00490_),
    .Y(_14404_));
 AO21x1_ASAP7_75t_R _19702_ (.A1(net2260),
    .A2(_00492_),
    .B(_14404_),
    .Y(_14405_));
 AOI221x1_ASAP7_75t_R _19703_ (.A1(_13377_),
    .A2(_14403_),
    .B1(_14405_),
    .B2(_13357_),
    .C(_14275_),
    .Y(_14406_));
 OR3x4_ASAP7_75t_R _19704_ (.A(net336),
    .B(net329),
    .C(net328),
    .Y(_14407_));
 AOI221x1_ASAP7_75t_R _19705_ (.A1(_00502_),
    .A2(_13390_),
    .B1(net2217),
    .B2(_00504_),
    .C(_14407_),
    .Y(_14408_));
 AND2x2_ASAP7_75t_R _19706_ (.A(net362),
    .B(_00503_),
    .Y(_14409_));
 AO21x1_ASAP7_75t_R _19707_ (.A1(net2260),
    .A2(_00505_),
    .B(_14409_),
    .Y(_14410_));
 NAND2x1_ASAP7_75t_R _19708_ (.A(net325),
    .B(_14410_),
    .Y(_14411_));
 INVx1_ASAP7_75t_R _19709_ (.A(_00501_),
    .Y(_14412_));
 NAND2x1_ASAP7_75t_R _19710_ (.A(net2257),
    .B(_00499_),
    .Y(_14413_));
 OA211x2_ASAP7_75t_R _19711_ (.A1(net2259),
    .A2(_14412_),
    .B(_14413_),
    .C(net325),
    .Y(_14414_));
 INVx1_ASAP7_75t_R _19712_ (.A(_00500_),
    .Y(_14415_));
 NAND2x1_ASAP7_75t_R _19713_ (.A(net2258),
    .B(_00498_),
    .Y(_14416_));
 OA211x2_ASAP7_75t_R _19714_ (.A1(net2266),
    .A2(_14415_),
    .B(_14416_),
    .C(net373),
    .Y(_14417_));
 OA211x2_ASAP7_75t_R _19715_ (.A1(_14414_),
    .A2(_14417_),
    .B(net334),
    .C(_13439_),
    .Y(_14418_));
 AO221x2_ASAP7_75t_R _19716_ (.A1(_14401_),
    .A2(_14406_),
    .B1(_14408_),
    .B2(_14411_),
    .C(_14418_),
    .Y(_14419_));
 OR2x6_ASAP7_75t_R _19717_ (.A(_14394_),
    .B(_14419_),
    .Y(_14420_));
 BUFx2_ASAP7_75t_R output213 (.A(net213),
    .Y(data_wdata_o[5]));
 AND2x2_ASAP7_75t_R _19719_ (.A(_13474_),
    .B(_14420_),
    .Y(_14422_));
 AO21x2_ASAP7_75t_R _19720_ (.A1(_13521_),
    .A2(_14363_),
    .B(_14422_),
    .Y(_18353_));
 INVx1_ASAP7_75t_R _19721_ (.A(_18353_),
    .Y(_18355_));
 INVx3_ASAP7_75t_R _19722_ (.A(_01742_),
    .Y(_14423_));
 OA21x2_ASAP7_75t_R _19723_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14356_),
    .Y(_14424_));
 INVx1_ASAP7_75t_R _19724_ (.A(_00518_),
    .Y(_14425_));
 NAND2x1_ASAP7_75t_R _19725_ (.A(net2276),
    .B(_00516_),
    .Y(_14426_));
 OA21x2_ASAP7_75t_R _19726_ (.A1(net2269),
    .A2(_14425_),
    .B(_14426_),
    .Y(_14427_));
 INVx1_ASAP7_75t_R _19727_ (.A(_00514_),
    .Y(_14428_));
 NAND2x1_ASAP7_75t_R _19728_ (.A(net2276),
    .B(_00512_),
    .Y(_14429_));
 OA21x2_ASAP7_75t_R _19729_ (.A1(net2269),
    .A2(_14428_),
    .B(_14429_),
    .Y(_14430_));
 AO221x1_ASAP7_75t_R _19730_ (.A1(_13366_),
    .A2(_14427_),
    .B1(_14430_),
    .B2(_13357_),
    .C(net329),
    .Y(_14431_));
 INVx1_ASAP7_75t_R _19731_ (.A(_00519_),
    .Y(_14432_));
 NAND2x1_ASAP7_75t_R _19732_ (.A(net336),
    .B(_00515_),
    .Y(_14433_));
 OA211x2_ASAP7_75t_R _19733_ (.A1(net336),
    .A2(_14432_),
    .B(_14433_),
    .C(net326),
    .Y(_14434_));
 INVx1_ASAP7_75t_R _19734_ (.A(_00517_),
    .Y(_14435_));
 NAND2x1_ASAP7_75t_R _19735_ (.A(net336),
    .B(_00513_),
    .Y(_14436_));
 OA211x2_ASAP7_75t_R _19736_ (.A1(net336),
    .A2(_14435_),
    .B(_14436_),
    .C(net2269),
    .Y(_14437_));
 OA21x2_ASAP7_75t_R _19737_ (.A1(_14434_),
    .A2(_14437_),
    .B(net323),
    .Y(_14438_));
 INVx1_ASAP7_75t_R _19738_ (.A(_00510_),
    .Y(_14439_));
 NAND2x1_ASAP7_75t_R _19739_ (.A(net2357),
    .B(_00508_),
    .Y(_14440_));
 OA211x2_ASAP7_75t_R _19740_ (.A1(net2269),
    .A2(_14439_),
    .B(_14440_),
    .C(net374),
    .Y(_14441_));
 INVx1_ASAP7_75t_R _19741_ (.A(_00511_),
    .Y(_14442_));
 NAND2x1_ASAP7_75t_R _19742_ (.A(net365),
    .B(_00509_),
    .Y(_14443_));
 OA211x2_ASAP7_75t_R _19743_ (.A1(net2269),
    .A2(_14442_),
    .B(_14443_),
    .C(net323),
    .Y(_14444_));
 OR3x1_ASAP7_75t_R _19744_ (.A(_14383_),
    .B(_14441_),
    .C(_14444_),
    .Y(_14445_));
 INVx1_ASAP7_75t_R _19745_ (.A(_00506_),
    .Y(_14446_));
 AND3x1_ASAP7_75t_R _19746_ (.A(net374),
    .B(net326),
    .C(_14446_),
    .Y(_14447_));
 INVx1_ASAP7_75t_R _19747_ (.A(_00507_),
    .Y(_14448_));
 NAND2x1_ASAP7_75t_R _19748_ (.A(net2357),
    .B(_01702_),
    .Y(_14449_));
 OA211x2_ASAP7_75t_R _19749_ (.A1(net2269),
    .A2(_14448_),
    .B(_14449_),
    .C(net323),
    .Y(_14450_));
 OA31x2_ASAP7_75t_R _19750_ (.A1(_13851_),
    .A2(_14447_),
    .A3(_14450_),
    .B1(net327),
    .Y(_14451_));
 OA211x2_ASAP7_75t_R _19751_ (.A1(_14431_),
    .A2(_14438_),
    .B(_14445_),
    .C(_14451_),
    .Y(_14452_));
 INVx1_ASAP7_75t_R _19752_ (.A(_00527_),
    .Y(_14453_));
 NAND2x1_ASAP7_75t_R _19753_ (.A(net2257),
    .B(_00525_),
    .Y(_14454_));
 OA211x2_ASAP7_75t_R _19754_ (.A1(net2259),
    .A2(_14453_),
    .B(_14454_),
    .C(net323),
    .Y(_14455_));
 INVx1_ASAP7_75t_R _19755_ (.A(_00526_),
    .Y(_14456_));
 NAND2x1_ASAP7_75t_R _19756_ (.A(net2257),
    .B(_00524_),
    .Y(_14457_));
 OA211x2_ASAP7_75t_R _19757_ (.A1(net2259),
    .A2(_14456_),
    .B(_14457_),
    .C(net374),
    .Y(_14458_));
 OR3x1_ASAP7_75t_R _19758_ (.A(net336),
    .B(_14455_),
    .C(_14458_),
    .Y(_14459_));
 AND2x2_ASAP7_75t_R _19759_ (.A(net2257),
    .B(_00521_),
    .Y(_14460_));
 AO21x1_ASAP7_75t_R _19760_ (.A1(net2278),
    .A2(_00523_),
    .B(_14460_),
    .Y(_14461_));
 AND2x2_ASAP7_75t_R _19761_ (.A(net2276),
    .B(_00520_),
    .Y(_14462_));
 AO21x1_ASAP7_75t_R _19762_ (.A1(net2278),
    .A2(_00522_),
    .B(_14462_),
    .Y(_14463_));
 AOI221x1_ASAP7_75t_R _19763_ (.A1(_13377_),
    .A2(_14461_),
    .B1(_14463_),
    .B2(_13357_),
    .C(_14275_),
    .Y(_14464_));
 BUFx2_ASAP7_75t_R output212 (.A(net212),
    .Y(data_wdata_o[4]));
 AND2x2_ASAP7_75t_R _19765_ (.A(net2276),
    .B(_00529_),
    .Y(_14466_));
 AO21x1_ASAP7_75t_R _19766_ (.A1(net2278),
    .A2(_00531_),
    .B(_14466_),
    .Y(_14467_));
 NAND2x1_ASAP7_75t_R _19767_ (.A(net323),
    .B(_14467_),
    .Y(_14468_));
 NAND2x1_ASAP7_75t_R _19768_ (.A(net336),
    .B(_13439_),
    .Y(_14469_));
 AOI221x1_ASAP7_75t_R _19769_ (.A1(_00528_),
    .A2(_13390_),
    .B1(net2227),
    .B2(_00530_),
    .C(_14469_),
    .Y(_14470_));
 INVx1_ASAP7_75t_R _19770_ (.A(_00535_),
    .Y(_14471_));
 NAND2x1_ASAP7_75t_R _19771_ (.A(net2357),
    .B(_00533_),
    .Y(_14472_));
 OA211x2_ASAP7_75t_R _19772_ (.A1(net2269),
    .A2(_14471_),
    .B(_14472_),
    .C(net323),
    .Y(_14473_));
 INVx1_ASAP7_75t_R _19773_ (.A(_00534_),
    .Y(_14474_));
 NAND2x1_ASAP7_75t_R _19774_ (.A(net2357),
    .B(_00532_),
    .Y(_14475_));
 OA211x2_ASAP7_75t_R _19775_ (.A1(net2269),
    .A2(_14474_),
    .B(_14475_),
    .C(net374),
    .Y(_14476_));
 OA211x2_ASAP7_75t_R _19776_ (.A1(_14473_),
    .A2(_14476_),
    .B(_13350_),
    .C(_13439_),
    .Y(_14477_));
 AO221x2_ASAP7_75t_R _19777_ (.A1(_14459_),
    .A2(_14464_),
    .B1(_14468_),
    .B2(_14470_),
    .C(_14477_),
    .Y(_14478_));
 OR2x6_ASAP7_75t_R _19778_ (.A(_14452_),
    .B(_14478_),
    .Y(_14479_));
 BUFx2_ASAP7_75t_R output211 (.A(net211),
    .Y(data_wdata_o[3]));
 AO22x2_ASAP7_75t_R _19780_ (.A1(_14423_),
    .A2(_14424_),
    .B1(_14479_),
    .B2(_13474_),
    .Y(_14481_));
 BUFx2_ASAP7_75t_R output210 (.A(net210),
    .Y(data_wdata_o[31]));
 INVx2_ASAP7_75t_R _19782_ (.A(_14481_),
    .Y(_18360_));
 INVx1_ASAP7_75t_R _19783_ (.A(_00549_),
    .Y(_14482_));
 NAND2x1_ASAP7_75t_R _19784_ (.A(net352),
    .B(_00547_),
    .Y(_14483_));
 OA211x2_ASAP7_75t_R _19785_ (.A1(net352),
    .A2(_14482_),
    .B(_14483_),
    .C(net323),
    .Y(_14484_));
 INVx1_ASAP7_75t_R _19786_ (.A(_00548_),
    .Y(_14485_));
 NAND2x1_ASAP7_75t_R _19787_ (.A(net352),
    .B(_00546_),
    .Y(_14486_));
 OA211x2_ASAP7_75t_R _19788_ (.A1(net352),
    .A2(_14485_),
    .B(_14486_),
    .C(net374),
    .Y(_14487_));
 BUFx2_ASAP7_75t_R output209 (.A(net209),
    .Y(data_wdata_o[30]));
 OA21x2_ASAP7_75t_R _19790_ (.A1(_14484_),
    .A2(_14487_),
    .B(_13350_),
    .Y(_14489_));
 INVx1_ASAP7_75t_R _19791_ (.A(_00544_),
    .Y(_14490_));
 NAND2x1_ASAP7_75t_R _19792_ (.A(net323),
    .B(_00545_),
    .Y(_14491_));
 OA211x2_ASAP7_75t_R _19793_ (.A1(net323),
    .A2(_14490_),
    .B(_14126_),
    .C(_14491_),
    .Y(_14492_));
 BUFx2_ASAP7_75t_R output208 (.A(net208),
    .Y(data_wdata_o[2]));
 INVx1_ASAP7_75t_R _19795_ (.A(_00543_),
    .Y(_14494_));
 NAND2x1_ASAP7_75t_R _19796_ (.A(net374),
    .B(_00542_),
    .Y(_14495_));
 OA211x2_ASAP7_75t_R _19797_ (.A1(net374),
    .A2(_14494_),
    .B(_14125_),
    .C(_14495_),
    .Y(_14496_));
 OR4x1_ASAP7_75t_R _19798_ (.A(net329),
    .B(_14489_),
    .C(_14492_),
    .D(_14496_),
    .Y(_14497_));
 BUFx2_ASAP7_75t_R output207 (.A(net207),
    .Y(data_wdata_o[29]));
 AND2x2_ASAP7_75t_R _19800_ (.A(net2257),
    .B(_00538_),
    .Y(_14499_));
 AO21x1_ASAP7_75t_R _19801_ (.A1(net2278),
    .A2(_00540_),
    .B(_14499_),
    .Y(_14500_));
 AND2x2_ASAP7_75t_R _19802_ (.A(net352),
    .B(_00539_),
    .Y(_14501_));
 AO21x1_ASAP7_75t_R _19803_ (.A1(net2278),
    .A2(_00541_),
    .B(_14501_),
    .Y(_14502_));
 AOI22x1_ASAP7_75t_R _19804_ (.A1(_13366_),
    .A2(_14500_),
    .B1(_14502_),
    .B2(net322),
    .Y(_14503_));
 INVx1_ASAP7_75t_R _19805_ (.A(_00536_),
    .Y(_14504_));
 INVx1_ASAP7_75t_R _19806_ (.A(_00537_),
    .Y(_14505_));
 NAND2x1_ASAP7_75t_R _19807_ (.A(net352),
    .B(_01701_),
    .Y(_14506_));
 OA21x2_ASAP7_75t_R _19808_ (.A1(net352),
    .A2(_14505_),
    .B(_14506_),
    .Y(_14507_));
 AO221x1_ASAP7_75t_R _19809_ (.A1(_14504_),
    .A2(net2242),
    .B1(_14507_),
    .B2(net323),
    .C(_13851_),
    .Y(_14508_));
 OA211x2_ASAP7_75t_R _19810_ (.A1(_13373_),
    .A2(_14503_),
    .B(_14508_),
    .C(net327),
    .Y(_14509_));
 INVx1_ASAP7_75t_R _19811_ (.A(_00564_),
    .Y(_14510_));
 NAND2x1_ASAP7_75t_R _19812_ (.A(net352),
    .B(_00562_),
    .Y(_14511_));
 OA211x2_ASAP7_75t_R _19813_ (.A1(net351),
    .A2(_14510_),
    .B(_14511_),
    .C(_13350_),
    .Y(_14512_));
 INVx1_ASAP7_75t_R _19814_ (.A(_00560_),
    .Y(_14513_));
 NAND2x1_ASAP7_75t_R _19815_ (.A(net351),
    .B(_00558_),
    .Y(_14514_));
 OA211x2_ASAP7_75t_R _19816_ (.A1(net351),
    .A2(_14513_),
    .B(_14514_),
    .C(net335),
    .Y(_14515_));
 OR3x1_ASAP7_75t_R _19817_ (.A(net325),
    .B(_14512_),
    .C(_14515_),
    .Y(_14516_));
 INVx1_ASAP7_75t_R _19818_ (.A(_00565_),
    .Y(_14517_));
 NAND2x1_ASAP7_75t_R _19819_ (.A(net351),
    .B(_00563_),
    .Y(_14518_));
 OA211x2_ASAP7_75t_R _19820_ (.A1(net351),
    .A2(_14517_),
    .B(_14518_),
    .C(_13350_),
    .Y(_14519_));
 INVx1_ASAP7_75t_R _19821_ (.A(_00561_),
    .Y(_14520_));
 NAND2x1_ASAP7_75t_R _19822_ (.A(net351),
    .B(_00559_),
    .Y(_14521_));
 OA211x2_ASAP7_75t_R _19823_ (.A1(net351),
    .A2(_14520_),
    .B(_14521_),
    .C(net335),
    .Y(_14522_));
 OR3x1_ASAP7_75t_R _19824_ (.A(net374),
    .B(_14519_),
    .C(_14522_),
    .Y(_14523_));
 INVx1_ASAP7_75t_R _19825_ (.A(_00556_),
    .Y(_14524_));
 NAND2x1_ASAP7_75t_R _19826_ (.A(net351),
    .B(_00554_),
    .Y(_14525_));
 OA211x2_ASAP7_75t_R _19827_ (.A1(net351),
    .A2(_14524_),
    .B(_14525_),
    .C(_13350_),
    .Y(_14526_));
 INVx1_ASAP7_75t_R _19828_ (.A(_00552_),
    .Y(_14527_));
 NAND2x1_ASAP7_75t_R _19829_ (.A(net351),
    .B(_00550_),
    .Y(_14528_));
 OA211x2_ASAP7_75t_R _19830_ (.A1(net351),
    .A2(_14527_),
    .B(_14528_),
    .C(net335),
    .Y(_14529_));
 OR3x1_ASAP7_75t_R _19831_ (.A(net325),
    .B(_14526_),
    .C(_14529_),
    .Y(_14530_));
 INVx1_ASAP7_75t_R _19832_ (.A(_00557_),
    .Y(_14531_));
 NAND2x1_ASAP7_75t_R _19833_ (.A(net352),
    .B(_00555_),
    .Y(_14532_));
 OA211x2_ASAP7_75t_R _19834_ (.A1(net352),
    .A2(_14531_),
    .B(_14532_),
    .C(_13350_),
    .Y(_14533_));
 INVx1_ASAP7_75t_R _19835_ (.A(_00553_),
    .Y(_14534_));
 NAND2x1_ASAP7_75t_R _19836_ (.A(net352),
    .B(_00551_),
    .Y(_14535_));
 OA211x2_ASAP7_75t_R _19837_ (.A1(net352),
    .A2(_14534_),
    .B(_14535_),
    .C(net335),
    .Y(_14536_));
 OR3x1_ASAP7_75t_R _19838_ (.A(net374),
    .B(_14533_),
    .C(_14536_),
    .Y(_14537_));
 AO33x2_ASAP7_75t_R _19839_ (.A1(_13439_),
    .A2(_14516_),
    .A3(_14523_),
    .B1(_14530_),
    .B2(_14537_),
    .B3(_13356_),
    .Y(_14538_));
 AO21x2_ASAP7_75t_R _19840_ (.A1(_14497_),
    .A2(_14509_),
    .B(_14538_),
    .Y(_14539_));
 INVx2_ASAP7_75t_R _19841_ (.A(_14539_),
    .Y(_14540_));
 BUFx2_ASAP7_75t_R output206 (.A(net206),
    .Y(data_wdata_o[28]));
 NAND2x1_ASAP7_75t_R _19843_ (.A(_13807_),
    .B(_13513_),
    .Y(_14542_));
 AO21x2_ASAP7_75t_R _19844_ (.A1(_13520_),
    .A2(_14542_),
    .B(_13497_),
    .Y(_14543_));
 OR3x1_ASAP7_75t_R _19845_ (.A(_01741_),
    .B(_13474_),
    .C(_14543_),
    .Y(_14544_));
 OAI21x1_ASAP7_75t_R _19846_ (.A1(_13521_),
    .A2(_14540_),
    .B(_14544_),
    .Y(_18363_));
 INVx1_ASAP7_75t_R _19847_ (.A(_18363_),
    .Y(_18365_));
 BUFx2_ASAP7_75t_R output205 (.A(net205),
    .Y(data_wdata_o[27]));
 INVx1_ASAP7_75t_R _19849_ (.A(_01740_),
    .Y(_14546_));
 BUFx2_ASAP7_75t_R output204 (.A(net204),
    .Y(data_wdata_o[26]));
 BUFx2_ASAP7_75t_R output203 (.A(net203),
    .Y(data_wdata_o[25]));
 INVx1_ASAP7_75t_R _19852_ (.A(_00578_),
    .Y(_14549_));
 NAND2x1_ASAP7_75t_R _19853_ (.A(net344),
    .B(_00576_),
    .Y(_14550_));
 OA211x2_ASAP7_75t_R _19854_ (.A1(net344),
    .A2(_14549_),
    .B(_13366_),
    .C(_14550_),
    .Y(_14551_));
 INVx1_ASAP7_75t_R _19855_ (.A(_00574_),
    .Y(_14552_));
 NAND2x1_ASAP7_75t_R _19856_ (.A(net368),
    .B(_00572_),
    .Y(_14553_));
 OA211x2_ASAP7_75t_R _19857_ (.A1(net344),
    .A2(_14552_),
    .B(_13357_),
    .C(_14553_),
    .Y(_14554_));
 INVx1_ASAP7_75t_R _19858_ (.A(_00579_),
    .Y(_14555_));
 NAND2x1_ASAP7_75t_R _19859_ (.A(net338),
    .B(_00575_),
    .Y(_14556_));
 OA211x2_ASAP7_75t_R _19860_ (.A1(net338),
    .A2(_14555_),
    .B(_14556_),
    .C(net326),
    .Y(_14557_));
 INVx1_ASAP7_75t_R _19861_ (.A(_00577_),
    .Y(_14558_));
 NAND2x1_ASAP7_75t_R _19862_ (.A(net338),
    .B(_00573_),
    .Y(_14559_));
 OA211x2_ASAP7_75t_R _19863_ (.A1(net338),
    .A2(_14558_),
    .B(_14559_),
    .C(net344),
    .Y(_14560_));
 OA21x2_ASAP7_75t_R _19864_ (.A1(_14557_),
    .A2(_14560_),
    .B(_13376_),
    .Y(_14561_));
 OR4x2_ASAP7_75t_R _19865_ (.A(_00245_),
    .B(_14551_),
    .C(_14554_),
    .D(_14561_),
    .Y(_14562_));
 AND2x2_ASAP7_75t_R _19866_ (.A(net2248),
    .B(_00568_),
    .Y(_14563_));
 AO21x1_ASAP7_75t_R _19867_ (.A1(net2278),
    .A2(_00570_),
    .B(_14563_),
    .Y(_14564_));
 AND2x2_ASAP7_75t_R _19868_ (.A(net346),
    .B(_00569_),
    .Y(_14565_));
 AO21x1_ASAP7_75t_R _19869_ (.A1(net2278),
    .A2(_00571_),
    .B(_14565_),
    .Y(_14566_));
 AOI22x1_ASAP7_75t_R _19870_ (.A1(_13366_),
    .A2(_14564_),
    .B1(_14566_),
    .B2(_13402_),
    .Y(_14567_));
 INVx1_ASAP7_75t_R _19871_ (.A(_00566_),
    .Y(_14568_));
 AND2x2_ASAP7_75t_R _19872_ (.A(net346),
    .B(_01700_),
    .Y(_14569_));
 AOI21x1_ASAP7_75t_R _19873_ (.A1(net2278),
    .A2(_00567_),
    .B(_14569_),
    .Y(_14570_));
 AO221x1_ASAP7_75t_R _19874_ (.A1(_14568_),
    .A2(net2242),
    .B1(_14570_),
    .B2(net323),
    .C(_13851_),
    .Y(_14571_));
 OA211x2_ASAP7_75t_R _19875_ (.A1(_13373_),
    .A2(_14567_),
    .B(_14571_),
    .C(net328),
    .Y(_14572_));
 INVx1_ASAP7_75t_R _19876_ (.A(_00587_),
    .Y(_14573_));
 NAND2x1_ASAP7_75t_R _19877_ (.A(net346),
    .B(_00585_),
    .Y(_14574_));
 OA211x2_ASAP7_75t_R _19878_ (.A1(net346),
    .A2(_14573_),
    .B(_13402_),
    .C(_14574_),
    .Y(_14575_));
 INVx1_ASAP7_75t_R _19879_ (.A(_00582_),
    .Y(_14576_));
 NAND2x1_ASAP7_75t_R _19880_ (.A(net346),
    .B(_00580_),
    .Y(_14577_));
 OA211x2_ASAP7_75t_R _19881_ (.A1(net346),
    .A2(_14576_),
    .B(_13357_),
    .C(_14577_),
    .Y(_14578_));
 INVx1_ASAP7_75t_R _19882_ (.A(_00586_),
    .Y(_14579_));
 NAND2x1_ASAP7_75t_R _19883_ (.A(net346),
    .B(_00584_),
    .Y(_14580_));
 OA211x2_ASAP7_75t_R _19884_ (.A1(net346),
    .A2(_14579_),
    .B(_13366_),
    .C(_14580_),
    .Y(_14581_));
 INVx1_ASAP7_75t_R _19885_ (.A(_00583_),
    .Y(_14582_));
 NAND2x1_ASAP7_75t_R _19886_ (.A(net346),
    .B(_00581_),
    .Y(_14583_));
 OA211x2_ASAP7_75t_R _19887_ (.A1(net346),
    .A2(_14582_),
    .B(_13377_),
    .C(_14583_),
    .Y(_14584_));
 OR4x1_ASAP7_75t_R _19888_ (.A(_14575_),
    .B(_14578_),
    .C(_14581_),
    .D(_14584_),
    .Y(_14585_));
 NAND2x1_ASAP7_75t_R _19889_ (.A(net323),
    .B(_00589_),
    .Y(_14586_));
 NAND2x1_ASAP7_75t_R _19890_ (.A(net374),
    .B(_00588_),
    .Y(_14587_));
 INVx1_ASAP7_75t_R _19891_ (.A(_00590_),
    .Y(_14588_));
 NOR2x1_ASAP7_75t_R _19892_ (.A(net374),
    .B(_00591_),
    .Y(_14589_));
 AO21x1_ASAP7_75t_R _19893_ (.A1(net374),
    .A2(_14588_),
    .B(_14589_),
    .Y(_14590_));
 AO32x1_ASAP7_75t_R _19894_ (.A1(_14125_),
    .A2(_14586_),
    .A3(_14587_),
    .B1(_14590_),
    .B2(_14126_),
    .Y(_14591_));
 AND2x2_ASAP7_75t_R _19895_ (.A(net2269),
    .B(_00593_),
    .Y(_14592_));
 AO21x1_ASAP7_75t_R _19896_ (.A1(net2278),
    .A2(_00595_),
    .B(_14592_),
    .Y(_14593_));
 AO21x1_ASAP7_75t_R _19897_ (.A1(_00592_),
    .A2(_13390_),
    .B(_14407_),
    .Y(_14594_));
 AOI221x1_ASAP7_75t_R _19898_ (.A1(_00594_),
    .A2(net2242),
    .B1(_14593_),
    .B2(net323),
    .C(_14594_),
    .Y(_14595_));
 AO21x1_ASAP7_75t_R _19899_ (.A1(_13439_),
    .A2(_14591_),
    .B(_14595_),
    .Y(_14596_));
 AO221x2_ASAP7_75t_R _19900_ (.A1(_14562_),
    .A2(_14572_),
    .B1(_14585_),
    .B2(_13356_),
    .C(_14596_),
    .Y(_14597_));
 BUFx2_ASAP7_75t_R output202 (.A(net202),
    .Y(data_wdata_o[24]));
 AO22x2_ASAP7_75t_R _19902_ (.A1(_14546_),
    .A2(_14424_),
    .B1(_14597_),
    .B2(_13474_),
    .Y(_14599_));
 BUFx2_ASAP7_75t_R output201 (.A(net201),
    .Y(data_wdata_o[23]));
 INVx1_ASAP7_75t_R _19904_ (.A(_14599_),
    .Y(_18370_));
 INVx1_ASAP7_75t_R _19905_ (.A(_00608_),
    .Y(_14600_));
 NAND2x1_ASAP7_75t_R _19906_ (.A(net361),
    .B(_00606_),
    .Y(_14601_));
 OA211x2_ASAP7_75t_R _19907_ (.A1(net361),
    .A2(_14600_),
    .B(_13366_),
    .C(_14601_),
    .Y(_14602_));
 AND2x2_ASAP7_75t_R _19908_ (.A(net361),
    .B(_00602_),
    .Y(_14603_));
 AO21x1_ASAP7_75t_R _19909_ (.A1(_13359_),
    .A2(_00604_),
    .B(_14603_),
    .Y(_14604_));
 OR2x2_ASAP7_75t_R _19910_ (.A(net361),
    .B(_00605_),
    .Y(_14605_));
 OA211x2_ASAP7_75t_R _19911_ (.A1(_13359_),
    .A2(_00603_),
    .B(_14605_),
    .C(net325),
    .Y(_14606_));
 AOI211x1_ASAP7_75t_R _19912_ (.A1(net373),
    .A2(_14604_),
    .B(_14606_),
    .C(_13350_),
    .Y(_14607_));
 INVx1_ASAP7_75t_R _19913_ (.A(_00609_),
    .Y(_14608_));
 NAND2x1_ASAP7_75t_R _19914_ (.A(net361),
    .B(_00607_),
    .Y(_14609_));
 OA211x2_ASAP7_75t_R _19915_ (.A1(net361),
    .A2(_14608_),
    .B(net322),
    .C(_14609_),
    .Y(_14610_));
 OR4x2_ASAP7_75t_R _19916_ (.A(net329),
    .B(_14602_),
    .C(_14607_),
    .D(_14610_),
    .Y(_14611_));
 BUFx2_ASAP7_75t_R output200 (.A(net200),
    .Y(data_wdata_o[22]));
 BUFx2_ASAP7_75t_R output199 (.A(net199),
    .Y(data_wdata_o[21]));
 AND2x2_ASAP7_75t_R _19919_ (.A(net362),
    .B(_01699_),
    .Y(_14614_));
 AO21x1_ASAP7_75t_R _19920_ (.A1(net2260),
    .A2(_00597_),
    .B(_14614_),
    .Y(_14615_));
 BUFx2_ASAP7_75t_R output198 (.A(net198),
    .Y(data_wdata_o[20]));
 OAI22x1_ASAP7_75t_R _19922_ (.A1(_00596_),
    .A2(_14184_),
    .B1(_14615_),
    .B2(net373),
    .Y(_14617_));
 INVx1_ASAP7_75t_R _19923_ (.A(_00601_),
    .Y(_14618_));
 NAND2x1_ASAP7_75t_R _19924_ (.A(net362),
    .B(_00599_),
    .Y(_14619_));
 OA211x2_ASAP7_75t_R _19925_ (.A1(net362),
    .A2(_14618_),
    .B(_14619_),
    .C(net325),
    .Y(_14620_));
 INVx1_ASAP7_75t_R _19926_ (.A(_00600_),
    .Y(_14621_));
 NAND2x1_ASAP7_75t_R _19927_ (.A(net362),
    .B(_00598_),
    .Y(_14622_));
 OA211x2_ASAP7_75t_R _19928_ (.A1(net362),
    .A2(_14621_),
    .B(_14622_),
    .C(net373),
    .Y(_14623_));
 OR3x1_ASAP7_75t_R _19929_ (.A(_14383_),
    .B(_14620_),
    .C(_14623_),
    .Y(_14624_));
 OA211x2_ASAP7_75t_R _19930_ (.A1(_13851_),
    .A2(_14617_),
    .B(_14624_),
    .C(net327),
    .Y(_14625_));
 INVx1_ASAP7_75t_R _19931_ (.A(_00617_),
    .Y(_14626_));
 NAND2x1_ASAP7_75t_R _19932_ (.A(net361),
    .B(_00615_),
    .Y(_14627_));
 OA211x2_ASAP7_75t_R _19933_ (.A1(net361),
    .A2(_14626_),
    .B(_14627_),
    .C(net325),
    .Y(_14628_));
 INVx1_ASAP7_75t_R _19934_ (.A(_00616_),
    .Y(_14629_));
 NAND2x1_ASAP7_75t_R _19935_ (.A(net362),
    .B(_00614_),
    .Y(_14630_));
 OA211x2_ASAP7_75t_R _19936_ (.A1(net362),
    .A2(_14629_),
    .B(_14630_),
    .C(net373),
    .Y(_14631_));
 OR3x1_ASAP7_75t_R _19937_ (.A(net334),
    .B(_14628_),
    .C(_14631_),
    .Y(_14632_));
 AND2x2_ASAP7_75t_R _19938_ (.A(net362),
    .B(_00611_),
    .Y(_14633_));
 AO21x1_ASAP7_75t_R _19939_ (.A1(_13359_),
    .A2(_00613_),
    .B(_14633_),
    .Y(_14634_));
 AND2x2_ASAP7_75t_R _19940_ (.A(net362),
    .B(_00610_),
    .Y(_14635_));
 AO21x1_ASAP7_75t_R _19941_ (.A1(_13359_),
    .A2(_00612_),
    .B(_14635_),
    .Y(_14636_));
 AOI22x1_ASAP7_75t_R _19942_ (.A1(_13377_),
    .A2(_14634_),
    .B1(_14636_),
    .B2(_13357_),
    .Y(_14637_));
 INVx1_ASAP7_75t_R _19943_ (.A(_00624_),
    .Y(_14638_));
 NAND2x1_ASAP7_75t_R _19944_ (.A(net361),
    .B(_00622_),
    .Y(_14639_));
 OA211x2_ASAP7_75t_R _19945_ (.A1(net361),
    .A2(_14638_),
    .B(_14639_),
    .C(net373),
    .Y(_14640_));
 INVx1_ASAP7_75t_R _19946_ (.A(_00625_),
    .Y(_14641_));
 NAND2x1_ASAP7_75t_R _19947_ (.A(net361),
    .B(_00623_),
    .Y(_14642_));
 OA211x2_ASAP7_75t_R _19948_ (.A1(net361),
    .A2(_14641_),
    .B(_14642_),
    .C(net325),
    .Y(_14643_));
 OR3x1_ASAP7_75t_R _19949_ (.A(net334),
    .B(_14640_),
    .C(_14643_),
    .Y(_14644_));
 AND2x2_ASAP7_75t_R _19950_ (.A(net361),
    .B(_00619_),
    .Y(_14645_));
 AO21x1_ASAP7_75t_R _19951_ (.A1(_13359_),
    .A2(_00621_),
    .B(_14645_),
    .Y(_14646_));
 AND2x2_ASAP7_75t_R _19952_ (.A(net361),
    .B(_00618_),
    .Y(_14647_));
 AO21x1_ASAP7_75t_R _19953_ (.A1(_13359_),
    .A2(_00620_),
    .B(_14647_),
    .Y(_14648_));
 AOI22x1_ASAP7_75t_R _19954_ (.A1(_13377_),
    .A2(_14646_),
    .B1(_14648_),
    .B2(_13357_),
    .Y(_14649_));
 AO33x2_ASAP7_75t_R _19955_ (.A1(_13356_),
    .A2(_14632_),
    .A3(_14637_),
    .B1(_14644_),
    .B2(_14649_),
    .B3(_13439_),
    .Y(_14650_));
 AOI21x1_ASAP7_75t_R _19956_ (.A1(_14611_),
    .A2(_14625_),
    .B(_14650_),
    .Y(_14651_));
 INVx3_ASAP7_75t_R _19957_ (.A(_14651_),
    .Y(_14652_));
 AO22x2_ASAP7_75t_R _19958_ (.A1(_13595_),
    .A2(_14424_),
    .B1(_14652_),
    .B2(_13474_),
    .Y(_14653_));
 BUFx2_ASAP7_75t_R output197 (.A(net197),
    .Y(data_wdata_o[1]));
 INVx2_ASAP7_75t_R _19960_ (.A(_14653_),
    .Y(_18375_));
 INVx1_ASAP7_75t_R _19961_ (.A(_00634_),
    .Y(_14654_));
 NAND2x1_ASAP7_75t_R _19962_ (.A(net2258),
    .B(_00632_),
    .Y(_14655_));
 OA211x2_ASAP7_75t_R _19963_ (.A1(net2258),
    .A2(_14654_),
    .B(_13357_),
    .C(_14655_),
    .Y(_14656_));
 INVx1_ASAP7_75t_R _19964_ (.A(_00635_),
    .Y(_14657_));
 NAND2x1_ASAP7_75t_R _19965_ (.A(net2258),
    .B(_00633_),
    .Y(_14658_));
 OA211x2_ASAP7_75t_R _19966_ (.A1(net2267),
    .A2(_14657_),
    .B(_13377_),
    .C(_14658_),
    .Y(_14659_));
 INVx1_ASAP7_75t_R _19967_ (.A(_00638_),
    .Y(_14660_));
 NAND2x1_ASAP7_75t_R _19968_ (.A(net2258),
    .B(_00636_),
    .Y(_14661_));
 OA211x2_ASAP7_75t_R _19969_ (.A1(net2266),
    .A2(_14660_),
    .B(_13366_),
    .C(_14661_),
    .Y(_14662_));
 INVx1_ASAP7_75t_R _19970_ (.A(_00639_),
    .Y(_14663_));
 NAND2x1_ASAP7_75t_R _19971_ (.A(net2258),
    .B(_00637_),
    .Y(_14664_));
 OA211x2_ASAP7_75t_R _19972_ (.A1(net360),
    .A2(_14663_),
    .B(net322),
    .C(_14664_),
    .Y(_14665_));
 OR5x2_ASAP7_75t_R _19973_ (.A(net330),
    .B(_14656_),
    .C(_14659_),
    .D(_14662_),
    .E(_14665_),
    .Y(_14666_));
 AND2x2_ASAP7_75t_R _19974_ (.A(net2258),
    .B(_00628_),
    .Y(_14667_));
 AO21x1_ASAP7_75t_R _19975_ (.A1(net2278),
    .A2(_00630_),
    .B(_14667_),
    .Y(_14668_));
 AND2x2_ASAP7_75t_R _19976_ (.A(net2258),
    .B(_00629_),
    .Y(_14669_));
 AO21x1_ASAP7_75t_R _19977_ (.A1(net2260),
    .A2(_00631_),
    .B(_14669_),
    .Y(_14670_));
 AOI22x1_ASAP7_75t_R _19978_ (.A1(_13366_),
    .A2(_14668_),
    .B1(_14670_),
    .B2(net322),
    .Y(_14671_));
 INVx1_ASAP7_75t_R _19979_ (.A(_00626_),
    .Y(_14672_));
 INVx1_ASAP7_75t_R _19980_ (.A(_00627_),
    .Y(_14673_));
 NAND2x1_ASAP7_75t_R _19981_ (.A(net2333),
    .B(_01698_),
    .Y(_14674_));
 OA21x2_ASAP7_75t_R _19982_ (.A1(net2333),
    .A2(_14673_),
    .B(_14674_),
    .Y(_14675_));
 AO221x1_ASAP7_75t_R _19983_ (.A1(_14672_),
    .A2(net2227),
    .B1(_14675_),
    .B2(net325),
    .C(_13851_),
    .Y(_14676_));
 OA211x2_ASAP7_75t_R _19984_ (.A1(_13373_),
    .A2(_14671_),
    .B(_14676_),
    .C(net327),
    .Y(_14677_));
 INVx1_ASAP7_75t_R _19985_ (.A(_00650_),
    .Y(_14678_));
 NOR2x1_ASAP7_75t_R _19986_ (.A(net373),
    .B(_00651_),
    .Y(_14679_));
 AO21x1_ASAP7_75t_R _19987_ (.A1(net373),
    .A2(_14678_),
    .B(_14679_),
    .Y(_14680_));
 INVx1_ASAP7_75t_R _19988_ (.A(_00649_),
    .Y(_14681_));
 NAND2x1_ASAP7_75t_R _19989_ (.A(net373),
    .B(_00648_),
    .Y(_14682_));
 OA211x2_ASAP7_75t_R _19990_ (.A1(net373),
    .A2(_14681_),
    .B(_14125_),
    .C(_14682_),
    .Y(_14683_));
 AO21x1_ASAP7_75t_R _19991_ (.A1(net2222),
    .A2(_14680_),
    .B(_14683_),
    .Y(_14684_));
 AND2x2_ASAP7_75t_R _19992_ (.A(net2257),
    .B(_00653_),
    .Y(_14685_));
 AO21x1_ASAP7_75t_R _19993_ (.A1(net2278),
    .A2(_00655_),
    .B(_14685_),
    .Y(_14686_));
 AO21x1_ASAP7_75t_R _19994_ (.A1(_00652_),
    .A2(_13390_),
    .B(_14407_),
    .Y(_14687_));
 AOI221x1_ASAP7_75t_R _19995_ (.A1(_00654_),
    .A2(net2227),
    .B1(_14686_),
    .B2(net325),
    .C(_14687_),
    .Y(_14688_));
 AO21x1_ASAP7_75t_R _19996_ (.A1(_13439_),
    .A2(_14684_),
    .B(_14688_),
    .Y(_14689_));
 NAND2x1_ASAP7_75t_R _19997_ (.A(net2333),
    .B(_00645_),
    .Y(_14690_));
 NAND2x1_ASAP7_75t_R _19998_ (.A(net2278),
    .B(_00647_),
    .Y(_14691_));
 NAND2x1_ASAP7_75t_R _19999_ (.A(net2333),
    .B(_00641_),
    .Y(_14692_));
 NAND2x1_ASAP7_75t_R _20000_ (.A(net2278),
    .B(_00643_),
    .Y(_14693_));
 AO33x2_ASAP7_75t_R _20001_ (.A1(net322),
    .A2(_14690_),
    .A3(_14691_),
    .B1(_14692_),
    .B2(_14693_),
    .B3(_13377_),
    .Y(_14694_));
 INVx1_ASAP7_75t_R _20002_ (.A(_00644_),
    .Y(_14695_));
 NOR2x1_ASAP7_75t_R _20003_ (.A(net2333),
    .B(_00646_),
    .Y(_14696_));
 AO21x1_ASAP7_75t_R _20004_ (.A1(net2333),
    .A2(_14695_),
    .B(_14696_),
    .Y(_14697_));
 INVx1_ASAP7_75t_R _20005_ (.A(_00642_),
    .Y(_14698_));
 NAND2x1_ASAP7_75t_R _20006_ (.A(net2333),
    .B(_00640_),
    .Y(_14699_));
 OA211x2_ASAP7_75t_R _20007_ (.A1(net2333),
    .A2(_14698_),
    .B(_13357_),
    .C(_14699_),
    .Y(_14700_));
 AO21x1_ASAP7_75t_R _20008_ (.A1(_13366_),
    .A2(_14697_),
    .B(_14700_),
    .Y(_14701_));
 OA21x2_ASAP7_75t_R _20009_ (.A1(_14694_),
    .A2(_14701_),
    .B(_13356_),
    .Y(_14702_));
 AOI211x1_ASAP7_75t_R _20010_ (.A1(_14666_),
    .A2(_14677_),
    .B(_14689_),
    .C(_14702_),
    .Y(_14703_));
 INVx3_ASAP7_75t_R _20011_ (.A(_00280_),
    .Y(_14704_));
 AND3x1_ASAP7_75t_R _20012_ (.A(_13890_),
    .B(_13476_),
    .C(_13465_),
    .Y(_14705_));
 AO31x2_ASAP7_75t_R _20013_ (.A1(_14704_),
    .A2(_13478_),
    .A3(_13482_),
    .B(_14705_),
    .Y(_14706_));
 AND3x1_ASAP7_75t_R _20014_ (.A(_13807_),
    .B(_13473_),
    .C(_13513_),
    .Y(_14707_));
 AND2x2_ASAP7_75t_R _20015_ (.A(net323),
    .B(_13505_),
    .Y(_14708_));
 AOI22x1_ASAP7_75t_R _20016_ (.A1(_14706_),
    .A2(_14707_),
    .B1(_14708_),
    .B2(_13495_),
    .Y(_14709_));
 OA21x2_ASAP7_75t_R _20017_ (.A1(_13521_),
    .A2(_14703_),
    .B(_14709_),
    .Y(_14710_));
 BUFx2_ASAP7_75t_R output196 (.A(net196),
    .Y(data_wdata_o[19]));
 INVx4_ASAP7_75t_R _20019_ (.A(_14710_),
    .Y(_18380_));
 INVx1_ASAP7_75t_R _20020_ (.A(_01476_),
    .Y(\cs_registers_i.mhpmcounter[2][12] ));
 INVx1_ASAP7_75t_R _20021_ (.A(_01507_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[12] ));
 INVx2_ASAP7_75t_R _20022_ (.A(_18385_),
    .Y(_18383_));
 AND5x2_ASAP7_75t_R _20023_ (.A(net2264),
    .B(net2213),
    .C(net2302),
    .D(_00287_),
    .E(net378),
    .Y(_14711_));
 AND2x2_ASAP7_75t_R _20024_ (.A(_13559_),
    .B(_14711_),
    .Y(_14712_));
 OR3x4_ASAP7_75t_R _20025_ (.A(_00281_),
    .B(_13784_),
    .C(_14712_),
    .Y(_17812_));
 INVx1_ASAP7_75t_R _20026_ (.A(_17812_),
    .Y(_17816_));
 NOR3x2_ASAP7_75t_R _20027_ (.B(_13784_),
    .C(_14711_),
    .Y(_14713_),
    .A(_00282_));
 CKINVDCx9p33_ASAP7_75t_R _20028_ (.A(_14713_),
    .Y(_14714_));
 BUFx2_ASAP7_75t_R output195 (.A(net195),
    .Y(data_wdata_o[18]));
 INVx2_ASAP7_75t_R _20030_ (.A(_00196_),
    .Y(\cs_registers_i.pc_id_i[11] ));
 BUFx2_ASAP7_75t_R output194 (.A(net194),
    .Y(data_wdata_o[17]));
 INVx1_ASAP7_75t_R _20032_ (.A(_00646_),
    .Y(_14716_));
 BUFx2_ASAP7_75t_R output193 (.A(net193),
    .Y(data_wdata_o[16]));
 NAND2x1_ASAP7_75t_R _20034_ (.A(net407),
    .B(_00644_),
    .Y(_14718_));
 OA211x2_ASAP7_75t_R _20035_ (.A1(net407),
    .A2(_14716_),
    .B(_14718_),
    .C(net320),
    .Y(_14719_));
 BUFx2_ASAP7_75t_R output192 (.A(net192),
    .Y(data_wdata_o[15]));
 BUFx2_ASAP7_75t_R output191 (.A(net191),
    .Y(data_wdata_o[14]));
 NAND2x1_ASAP7_75t_R _20038_ (.A(net407),
    .B(_00640_),
    .Y(_14722_));
 OA211x2_ASAP7_75t_R _20039_ (.A1(net407),
    .A2(_14698_),
    .B(_14722_),
    .C(net385),
    .Y(_14723_));
 OR3x1_ASAP7_75t_R _20040_ (.A(net318),
    .B(_14719_),
    .C(_14723_),
    .Y(_14724_));
 BUFx2_ASAP7_75t_R output190 (.A(net190),
    .Y(data_wdata_o[13]));
 INVx1_ASAP7_75t_R _20042_ (.A(_00647_),
    .Y(_14726_));
 NAND2x1_ASAP7_75t_R _20043_ (.A(net407),
    .B(_00645_),
    .Y(_14727_));
 OA211x2_ASAP7_75t_R _20044_ (.A1(net401),
    .A2(_14726_),
    .B(_14727_),
    .C(net320),
    .Y(_14728_));
 INVx1_ASAP7_75t_R _20045_ (.A(_00643_),
    .Y(_14729_));
 NAND2x1_ASAP7_75t_R _20046_ (.A(net407),
    .B(_00641_),
    .Y(_14730_));
 OA211x2_ASAP7_75t_R _20047_ (.A1(net407),
    .A2(_14729_),
    .B(_14730_),
    .C(net385),
    .Y(_14731_));
 OR3x1_ASAP7_75t_R _20048_ (.A(net422),
    .B(_14728_),
    .C(_14731_),
    .Y(_14732_));
 BUFx2_ASAP7_75t_R output189 (.A(net189),
    .Y(data_wdata_o[12]));
 INVx1_ASAP7_75t_R _20050_ (.A(_00630_),
    .Y(_14734_));
 NAND2x1_ASAP7_75t_R _20051_ (.A(net401),
    .B(_00628_),
    .Y(_14735_));
 OA211x2_ASAP7_75t_R _20052_ (.A1(net401),
    .A2(_14734_),
    .B(_14735_),
    .C(net422),
    .Y(_14736_));
 INVx1_ASAP7_75t_R _20053_ (.A(_00631_),
    .Y(_14737_));
 NAND2x1_ASAP7_75t_R _20054_ (.A(net400),
    .B(_00629_),
    .Y(_14738_));
 OA211x2_ASAP7_75t_R _20055_ (.A1(net400),
    .A2(_14737_),
    .B(_14738_),
    .C(net317),
    .Y(_14739_));
 OR3x1_ASAP7_75t_R _20056_ (.A(net312),
    .B(_14736_),
    .C(_14739_),
    .Y(_14740_));
 NAND2x1_ASAP7_75t_R _20057_ (.A(net401),
    .B(_01698_),
    .Y(_14741_));
 OA211x2_ASAP7_75t_R _20058_ (.A1(net401),
    .A2(_14673_),
    .B(_14741_),
    .C(net318),
    .Y(_14742_));
 BUFx2_ASAP7_75t_R output188 (.A(net188),
    .Y(data_wdata_o[11]));
 BUFx2_ASAP7_75t_R output187 (.A(net187),
    .Y(data_wdata_o[10]));
 NOR2x1_ASAP7_75t_R _20061_ (.A(net401),
    .B(_00626_),
    .Y(_14745_));
 BUFx2_ASAP7_75t_R output186 (.A(net186),
    .Y(data_wdata_o[0]));
 AO21x1_ASAP7_75t_R _20063_ (.A1(net422),
    .A2(_14745_),
    .B(net315),
    .Y(_14747_));
 OA21x2_ASAP7_75t_R _20064_ (.A1(_14742_),
    .A2(_14747_),
    .B(net377),
    .Y(_14748_));
 AO32x1_ASAP7_75t_R _20065_ (.A1(_13626_),
    .A2(_14724_),
    .A3(_14732_),
    .B1(_14740_),
    .B2(_14748_),
    .Y(_14749_));
 BUFx2_ASAP7_75t_R output185 (.A(net185),
    .Y(data_req_o));
 BUFx2_ASAP7_75t_R output184 (.A(net184),
    .Y(data_be_o[3]));
 NAND2x1_ASAP7_75t_R _20068_ (.A(net400),
    .B(_00633_),
    .Y(_14752_));
 OA211x2_ASAP7_75t_R _20069_ (.A1(net400),
    .A2(_14657_),
    .B(_14752_),
    .C(net318),
    .Y(_14753_));
 NAND2x1_ASAP7_75t_R _20070_ (.A(net400),
    .B(_00632_),
    .Y(_14754_));
 OA211x2_ASAP7_75t_R _20071_ (.A1(net400),
    .A2(_14654_),
    .B(_14754_),
    .C(net421),
    .Y(_14755_));
 OR3x1_ASAP7_75t_R _20072_ (.A(net320),
    .B(_14753_),
    .C(_14755_),
    .Y(_14756_));
 NAND2x1_ASAP7_75t_R _20073_ (.A(net401),
    .B(_00637_),
    .Y(_14757_));
 OA211x2_ASAP7_75t_R _20074_ (.A1(net401),
    .A2(_14663_),
    .B(_14757_),
    .C(net318),
    .Y(_14758_));
 NAND2x1_ASAP7_75t_R _20075_ (.A(net401),
    .B(_00636_),
    .Y(_14759_));
 OA211x2_ASAP7_75t_R _20076_ (.A1(net401),
    .A2(_14660_),
    .B(_14759_),
    .C(net421),
    .Y(_14760_));
 OR3x1_ASAP7_75t_R _20077_ (.A(net384),
    .B(_14758_),
    .C(_14760_),
    .Y(_14761_));
 AND2x2_ASAP7_75t_R _20078_ (.A(_14756_),
    .B(_14761_),
    .Y(_14762_));
 AND2x2_ASAP7_75t_R _20079_ (.A(_14740_),
    .B(_14748_),
    .Y(_14763_));
 BUFx2_ASAP7_75t_R output183 (.A(net183),
    .Y(data_be_o[2]));
 BUFx2_ASAP7_75t_R output182 (.A(net182),
    .Y(data_be_o[1]));
 NOR2x1_ASAP7_75t_R _20082_ (.A(net384),
    .B(_00654_),
    .Y(_14766_));
 AO21x1_ASAP7_75t_R _20083_ (.A1(net384),
    .A2(_14678_),
    .B(_14766_),
    .Y(_14767_));
 INVx1_ASAP7_75t_R _20084_ (.A(_00655_),
    .Y(_14768_));
 NAND2x1_ASAP7_75t_R _20085_ (.A(net384),
    .B(_00651_),
    .Y(_14769_));
 BUFx2_ASAP7_75t_R output181 (.A(net181),
    .Y(data_be_o[0]));
 BUFx2_ASAP7_75t_R output180 (.A(net2203),
    .Y(data_addr_o[9]));
 OA211x2_ASAP7_75t_R _20088_ (.A1(net384),
    .A2(_14768_),
    .B(_14769_),
    .C(net318),
    .Y(_14772_));
 AO21x1_ASAP7_75t_R _20089_ (.A1(net422),
    .A2(_14767_),
    .B(_14772_),
    .Y(_14773_));
 INVx1_ASAP7_75t_R _20090_ (.A(_00653_),
    .Y(_14774_));
 NAND2x1_ASAP7_75t_R _20091_ (.A(net422),
    .B(_00652_),
    .Y(_14775_));
 OA211x2_ASAP7_75t_R _20092_ (.A1(net422),
    .A2(_14774_),
    .B(_14775_),
    .C(net320),
    .Y(_14776_));
 NAND2x1_ASAP7_75t_R _20093_ (.A(net422),
    .B(_00648_),
    .Y(_14777_));
 OA211x2_ASAP7_75t_R _20094_ (.A1(net422),
    .A2(_14681_),
    .B(_14777_),
    .C(net384),
    .Y(_14778_));
 OR3x1_ASAP7_75t_R _20095_ (.A(net316),
    .B(_14776_),
    .C(_14778_),
    .Y(_14779_));
 NOR2x2_ASAP7_75t_R _20096_ (.A(net382),
    .B(net378),
    .Y(_14780_));
 BUFx2_ASAP7_75t_R output179 (.A(net179),
    .Y(data_addr_o[8]));
 OA211x2_ASAP7_75t_R _20098_ (.A1(net408),
    .A2(_14773_),
    .B(_14779_),
    .C(_14780_),
    .Y(_14782_));
 AO221x2_ASAP7_75t_R _20099_ (.A1(net379),
    .A2(_14749_),
    .B1(_14762_),
    .B2(_14763_),
    .C(_14782_),
    .Y(_14783_));
 BUFx2_ASAP7_75t_R output178 (.A(net178),
    .Y(data_addr_o[7]));
 BUFx2_ASAP7_75t_R output177 (.A(net177),
    .Y(data_addr_o[6]));
 INVx1_ASAP7_75t_R _20102_ (.A(_01630_),
    .Y(_14786_));
 AO32x2_ASAP7_75t_R _20103_ (.A1(\cs_registers_i.pc_id_i[11] ),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_14786_),
    .B2(_13450_),
    .Y(_14787_));
 AOI21x1_ASAP7_75t_R _20104_ (.A1(_13810_),
    .A2(_14783_),
    .B(_14787_),
    .Y(_18379_));
 INVx1_ASAP7_75t_R _20105_ (.A(_01487_),
    .Y(\cs_registers_i.mhpmcounter[2][1] ));
 INVx1_ASAP7_75t_R _20106_ (.A(_01518_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[1] ));
 INVx1_ASAP7_75t_R _20107_ (.A(_18332_),
    .Y(_18330_));
 INVx1_ASAP7_75t_R _20108_ (.A(_02066_),
    .Y(\cs_registers_i.mhpmcounter[2][32] ));
 INVx1_ASAP7_75t_R _20109_ (.A(_02172_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[32] ));
 INVx1_ASAP7_75t_R _20110_ (.A(_01732_),
    .Y(_14788_));
 BUFx2_ASAP7_75t_R output176 (.A(net289),
    .Y(data_addr_o[5]));
 BUFx2_ASAP7_75t_R output175 (.A(net175),
    .Y(data_addr_o[4]));
 INVx5_ASAP7_75t_R _20113_ (.A(_01717_),
    .Y(_14791_));
 BUFx2_ASAP7_75t_R output174 (.A(net293),
    .Y(data_addr_o[3]));
 INVx3_ASAP7_75t_R _20115_ (.A(_01715_),
    .Y(_14793_));
 AND3x4_ASAP7_75t_R _20116_ (.A(_01714_),
    .B(_14793_),
    .C(_01716_),
    .Y(_14794_));
 BUFx2_ASAP7_75t_R output173 (.A(net173),
    .Y(data_addr_o[31]));
 AND2x6_ASAP7_75t_R _20118_ (.A(_14791_),
    .B(_14794_),
    .Y(_14796_));
 AND3x4_ASAP7_75t_R _20119_ (.A(_13459_),
    .B(_01721_),
    .C(_14796_),
    .Y(_14797_));
 BUFx2_ASAP7_75t_R output172 (.A(net172),
    .Y(data_addr_o[30]));
 OR5x2_ASAP7_75t_R _20121_ (.A(net323),
    .B(net2277),
    .C(_01740_),
    .D(_01741_),
    .E(_13851_),
    .Y(_14799_));
 BUFx2_ASAP7_75t_R output171 (.A(net171),
    .Y(data_addr_o[2]));
 INVx1_ASAP7_75t_R _20123_ (.A(_01741_),
    .Y(_14801_));
 NAND2x1_ASAP7_75t_R _20124_ (.A(_01740_),
    .B(_14801_),
    .Y(_14802_));
 NAND2x2_ASAP7_75t_R _20125_ (.A(net323),
    .B(net2277),
    .Y(_14803_));
 OR3x1_ASAP7_75t_R _20126_ (.A(_14383_),
    .B(_14802_),
    .C(_14803_),
    .Y(_14804_));
 OR4x1_ASAP7_75t_R _20127_ (.A(_00244_),
    .B(_01739_),
    .C(_01742_),
    .D(_01743_),
    .Y(_14805_));
 OR3x2_ASAP7_75t_R _20128_ (.A(_14704_),
    .B(_14362_),
    .C(_14805_),
    .Y(_14806_));
 AND4x2_ASAP7_75t_R _20129_ (.A(_00244_),
    .B(_00280_),
    .C(_01739_),
    .D(_01743_),
    .Y(_14807_));
 NAND2x2_ASAP7_75t_R _20130_ (.A(_13531_),
    .B(_14807_),
    .Y(_14808_));
 OA21x2_ASAP7_75t_R _20131_ (.A1(_14799_),
    .A2(_14806_),
    .B(_14808_),
    .Y(_14809_));
 AOI21x1_ASAP7_75t_R _20132_ (.A1(_14799_),
    .A2(_14804_),
    .B(_14809_),
    .Y(_14810_));
 AND2x2_ASAP7_75t_R _20133_ (.A(_00281_),
    .B(_00282_),
    .Y(_14811_));
 AND5x2_ASAP7_75t_R _20134_ (.A(_13460_),
    .B(_13456_),
    .C(_13476_),
    .D(_13801_),
    .E(_14811_),
    .Y(_14812_));
 AND2x2_ASAP7_75t_R _20135_ (.A(_13531_),
    .B(_14807_),
    .Y(_14813_));
 AND4x1_ASAP7_75t_R _20136_ (.A(net333),
    .B(_01740_),
    .C(_01741_),
    .D(_14125_),
    .Y(_14814_));
 NAND2x1_ASAP7_75t_R _20137_ (.A(_14813_),
    .B(_14814_),
    .Y(_14815_));
 NAND2x1_ASAP7_75t_R _20138_ (.A(_14812_),
    .B(_14815_),
    .Y(_14816_));
 AO22x1_ASAP7_75t_R _20139_ (.A1(_00279_),
    .A2(_13595_),
    .B1(_01743_),
    .B2(_13559_),
    .Y(_14817_));
 NAND2x1_ASAP7_75t_R _20140_ (.A(_13483_),
    .B(_14817_),
    .Y(_14818_));
 AND2x2_ASAP7_75t_R _20141_ (.A(_01739_),
    .B(_13592_),
    .Y(_14819_));
 AO221x1_ASAP7_75t_R _20142_ (.A1(_13611_),
    .A2(_14818_),
    .B1(_14819_),
    .B2(_13600_),
    .C(_13612_),
    .Y(_14820_));
 OAI21x1_ASAP7_75t_R _20143_ (.A1(_14810_),
    .A2(_14816_),
    .B(_14820_),
    .Y(_14821_));
 NAND3x1_ASAP7_75t_R _20144_ (.A(_13496_),
    .B(_00172_),
    .C(_13550_),
    .Y(_14822_));
 NAND2x1_ASAP7_75t_R _20145_ (.A(_00165_),
    .B(_13456_),
    .Y(_14823_));
 AO21x1_ASAP7_75t_R _20146_ (.A1(_13496_),
    .A2(_00172_),
    .B(_13479_),
    .Y(_14824_));
 AO21x1_ASAP7_75t_R _20147_ (.A1(_14823_),
    .A2(_14824_),
    .B(_13480_),
    .Y(_14825_));
 AND2x2_ASAP7_75t_R _20148_ (.A(_13496_),
    .B(_00168_),
    .Y(_14826_));
 AO32x1_ASAP7_75t_R _20149_ (.A1(_13587_),
    .A2(_14826_),
    .A3(_13558_),
    .B1(_13547_),
    .B2(_13570_),
    .Y(_14827_));
 AND4x2_ASAP7_75t_R _20150_ (.A(_00278_),
    .B(_00172_),
    .C(_13489_),
    .D(_13476_),
    .Y(_14828_));
 NAND2x1_ASAP7_75t_R _20151_ (.A(_00282_),
    .B(_00175_),
    .Y(_14829_));
 AO21x1_ASAP7_75t_R _20152_ (.A1(_13570_),
    .A2(_14829_),
    .B(_13592_),
    .Y(_14830_));
 AO21x1_ASAP7_75t_R _20153_ (.A1(_14828_),
    .A2(_14830_),
    .B(_13467_),
    .Y(_14831_));
 AO211x2_ASAP7_75t_R _20154_ (.A1(_14822_),
    .A2(_14825_),
    .B(_14827_),
    .C(_14831_),
    .Y(_14832_));
 NOR2x1_ASAP7_75t_R _20155_ (.A(_13616_),
    .B(_13580_),
    .Y(_14833_));
 AND2x6_ASAP7_75t_R _20156_ (.A(_00187_),
    .B(_00191_),
    .Y(_14834_));
 AND4x2_ASAP7_75t_R _20157_ (.A(_00279_),
    .B(_00323_),
    .C(_00184_),
    .D(_00194_),
    .Y(_14835_));
 NAND3x2_ASAP7_75t_R _20158_ (.B(_14834_),
    .C(_14835_),
    .Y(_14836_),
    .A(_14711_));
 INVx1_ASAP7_75t_R _20159_ (.A(_01847_),
    .Y(_14837_));
 AO221x1_ASAP7_75t_R _20160_ (.A1(_13574_),
    .A2(_14833_),
    .B1(_14812_),
    .B2(_14836_),
    .C(_14837_),
    .Y(_14838_));
 NOR2x1_ASAP7_75t_R _20161_ (.A(_13570_),
    .B(_13786_),
    .Y(_14839_));
 OA21x2_ASAP7_75t_R _20162_ (.A1(_13547_),
    .A2(_14839_),
    .B(_13559_),
    .Y(_14840_));
 OR3x2_ASAP7_75t_R _20163_ (.A(_14832_),
    .B(_14838_),
    .C(_14840_),
    .Y(_14841_));
 NOR2x2_ASAP7_75t_R _20164_ (.A(_14821_),
    .B(_14841_),
    .Y(_14842_));
 AND3x4_ASAP7_75t_R _20165_ (.A(_13817_),
    .B(_14797_),
    .C(_14842_),
    .Y(_14843_));
 BUFx2_ASAP7_75t_R output170 (.A(net2142),
    .Y(data_addr_o[29]));
 NAND2x2_ASAP7_75t_R _20167_ (.A(_00279_),
    .B(_14843_),
    .Y(_14845_));
 BUFx2_ASAP7_75t_R output169 (.A(net169),
    .Y(data_addr_o[28]));
 BUFx2_ASAP7_75t_R output168 (.A(net2156),
    .Y(data_addr_o[27]));
 BUFx2_ASAP7_75t_R output167 (.A(net167),
    .Y(data_addr_o[26]));
 BUFx2_ASAP7_75t_R output166 (.A(net2176),
    .Y(data_addr_o[25]));
 BUFx2_ASAP7_75t_R output165 (.A(net165),
    .Y(data_addr_o[24]));
 AO21x1_ASAP7_75t_R _20173_ (.A1(_13534_),
    .A2(_13803_),
    .B(_01874_),
    .Y(_14851_));
 AOI211x1_ASAP7_75t_R _20174_ (.A1(_01314_),
    .A2(_14851_),
    .B(_14845_),
    .C(_14362_),
    .Y(_14852_));
 AO21x1_ASAP7_75t_R _20175_ (.A1(_14788_),
    .A2(_14845_),
    .B(_14852_),
    .Y(_00000_));
 INVx2_ASAP7_75t_R _20176_ (.A(_00162_),
    .Y(\cs_registers_i.pc_id_i[2] ));
 OR3x1_ASAP7_75t_R _20177_ (.A(net2302),
    .B(_13784_),
    .C(_13808_),
    .Y(_14853_));
 OA21x2_ASAP7_75t_R _20178_ (.A1(_01639_),
    .A2(_13807_),
    .B(_14853_),
    .Y(_14854_));
 BUFx2_ASAP7_75t_R output164 (.A(net2178),
    .Y(data_addr_o[23]));
 BUFx2_ASAP7_75t_R output163 (.A(net163),
    .Y(data_addr_o[22]));
 NAND2x1_ASAP7_75t_R _20181_ (.A(net408),
    .B(_00374_),
    .Y(_14857_));
 BUFx2_ASAP7_75t_R output162 (.A(net258),
    .Y(data_addr_o[21]));
 BUFx2_ASAP7_75t_R output161 (.A(net161),
    .Y(data_addr_o[20]));
 OA211x2_ASAP7_75t_R _20184_ (.A1(net408),
    .A2(_14118_),
    .B(_14857_),
    .C(net318),
    .Y(_14860_));
 BUFx2_ASAP7_75t_R output160 (.A(net261),
    .Y(data_addr_o[19]));
 BUFx2_ASAP7_75t_R output159 (.A(net159),
    .Y(data_addr_o[18]));
 BUFx2_ASAP7_75t_R output158 (.A(net259),
    .Y(data_addr_o[17]));
 INVx1_ASAP7_75t_R _20188_ (.A(_00375_),
    .Y(_14864_));
 NAND2x1_ASAP7_75t_R _20189_ (.A(net408),
    .B(_00373_),
    .Y(_14865_));
 OA211x2_ASAP7_75t_R _20190_ (.A1(net408),
    .A2(_14864_),
    .B(_14865_),
    .C(net425),
    .Y(_14866_));
 OR3x1_ASAP7_75t_R _20191_ (.A(net385),
    .B(_14860_),
    .C(_14866_),
    .Y(_14867_));
 BUFx2_ASAP7_75t_R output157 (.A(net157),
    .Y(data_addr_o[16]));
 BUFx2_ASAP7_75t_R output156 (.A(net156),
    .Y(data_addr_o[15]));
 INVx1_ASAP7_75t_R _20194_ (.A(_00372_),
    .Y(_14870_));
 BUFx2_ASAP7_75t_R output155 (.A(net155),
    .Y(data_addr_o[14]));
 NAND2x1_ASAP7_75t_R _20196_ (.A(net409),
    .B(_00370_),
    .Y(_14872_));
 OA211x2_ASAP7_75t_R _20197_ (.A1(net409),
    .A2(_14870_),
    .B(_14872_),
    .C(net318),
    .Y(_14873_));
 INVx1_ASAP7_75t_R _20198_ (.A(_00371_),
    .Y(_14874_));
 NAND2x1_ASAP7_75t_R _20199_ (.A(net409),
    .B(_00369_),
    .Y(_14875_));
 OA211x2_ASAP7_75t_R _20200_ (.A1(net409),
    .A2(_14874_),
    .B(_14875_),
    .C(net422),
    .Y(_14876_));
 OR3x1_ASAP7_75t_R _20201_ (.A(net320),
    .B(_14873_),
    .C(_14876_),
    .Y(_14877_));
 INVx1_ASAP7_75t_R _20202_ (.A(_00359_),
    .Y(_14878_));
 NAND2x1_ASAP7_75t_R _20203_ (.A(net408),
    .B(_00357_),
    .Y(_14879_));
 OA211x2_ASAP7_75t_R _20204_ (.A1(net408),
    .A2(_14878_),
    .B(_14879_),
    .C(net422),
    .Y(_14880_));
 BUFx2_ASAP7_75t_R output154 (.A(net154),
    .Y(data_addr_o[13]));
 INVx1_ASAP7_75t_R _20206_ (.A(_00360_),
    .Y(_14882_));
 NAND2x1_ASAP7_75t_R _20207_ (.A(net408),
    .B(_00358_),
    .Y(_14883_));
 BUFx2_ASAP7_75t_R output153 (.A(net153),
    .Y(data_addr_o[12]));
 OA211x2_ASAP7_75t_R _20209_ (.A1(net408),
    .A2(_14882_),
    .B(_14883_),
    .C(net318),
    .Y(_14885_));
 OR3x1_ASAP7_75t_R _20210_ (.A(net312),
    .B(_14880_),
    .C(_14885_),
    .Y(_14886_));
 BUFx2_ASAP7_75t_R output152 (.A(net262),
    .Y(data_addr_o[11]));
 NAND2x1_ASAP7_75t_R _20212_ (.A(net422),
    .B(_00355_),
    .Y(_14888_));
 OA211x2_ASAP7_75t_R _20213_ (.A1(net422),
    .A2(_14162_),
    .B(_14888_),
    .C(net316),
    .Y(_14889_));
 INVx1_ASAP7_75t_R _20214_ (.A(_01707_),
    .Y(_14890_));
 AND3x1_ASAP7_75t_R _20215_ (.A(net318),
    .B(net409),
    .C(_14890_),
    .Y(_14891_));
 OA31x2_ASAP7_75t_R _20216_ (.A1(net315),
    .A2(_14889_),
    .A3(_14891_),
    .B1(net377),
    .Y(_14892_));
 AO32x1_ASAP7_75t_R _20217_ (.A1(_13626_),
    .A2(_14867_),
    .A3(_14877_),
    .B1(_14886_),
    .B2(_14892_),
    .Y(_14893_));
 NAND2x1_ASAP7_75t_R _20218_ (.A(net409),
    .B(_00366_),
    .Y(_14894_));
 OA211x2_ASAP7_75t_R _20219_ (.A1(net409),
    .A2(_14146_),
    .B(_14894_),
    .C(net318),
    .Y(_14895_));
 BUFx2_ASAP7_75t_R output151 (.A(net151),
    .Y(data_addr_o[10]));
 NAND2x1_ASAP7_75t_R _20221_ (.A(net409),
    .B(_00365_),
    .Y(_14897_));
 OA211x2_ASAP7_75t_R _20222_ (.A1(net409),
    .A2(_14143_),
    .B(_14897_),
    .C(net422),
    .Y(_14898_));
 OR3x1_ASAP7_75t_R _20223_ (.A(net385),
    .B(_14895_),
    .C(_14898_),
    .Y(_14899_));
 NAND2x1_ASAP7_75t_R _20224_ (.A(net409),
    .B(_00362_),
    .Y(_14900_));
 OA211x2_ASAP7_75t_R _20225_ (.A1(net409),
    .A2(_14151_),
    .B(_14900_),
    .C(net318),
    .Y(_14901_));
 BUFx2_ASAP7_75t_R output150 (.A(net150),
    .Y(core_sleep_o));
 NAND2x1_ASAP7_75t_R _20227_ (.A(net409),
    .B(_00361_),
    .Y(_14903_));
 OA211x2_ASAP7_75t_R _20228_ (.A1(net409),
    .A2(_14140_),
    .B(_14903_),
    .C(net422),
    .Y(_14904_));
 OR3x1_ASAP7_75t_R _20229_ (.A(net320),
    .B(_14901_),
    .C(_14904_),
    .Y(_14905_));
 AND2x2_ASAP7_75t_R _20230_ (.A(_14899_),
    .B(_14905_),
    .Y(_14906_));
 AND2x2_ASAP7_75t_R _20231_ (.A(_14886_),
    .B(_14892_),
    .Y(_14907_));
 INVx1_ASAP7_75t_R _20232_ (.A(_00377_),
    .Y(_14908_));
 BUFx2_ASAP7_75t_R input149 (.A(net3961),
    .Y(net149));
 NOR2x1_ASAP7_75t_R _20234_ (.A(net408),
    .B(_00379_),
    .Y(_14910_));
 AO21x1_ASAP7_75t_R _20235_ (.A1(net408),
    .A2(_14908_),
    .B(_14910_),
    .Y(_14911_));
 NAND2x1_ASAP7_75t_R _20236_ (.A(net408),
    .B(_00378_),
    .Y(_14912_));
 OA211x2_ASAP7_75t_R _20237_ (.A1(net408),
    .A2(_14127_),
    .B(_14912_),
    .C(net318),
    .Y(_14913_));
 AO21x1_ASAP7_75t_R _20238_ (.A1(net422),
    .A2(_14911_),
    .B(_14913_),
    .Y(_14914_));
 NAND2x1_ASAP7_75t_R _20239_ (.A(net408),
    .B(_00382_),
    .Y(_14915_));
 OA211x2_ASAP7_75t_R _20240_ (.A1(net408),
    .A2(_14135_),
    .B(_14915_),
    .C(net318),
    .Y(_14916_));
 NAND2x1_ASAP7_75t_R _20241_ (.A(net408),
    .B(_00381_),
    .Y(_14917_));
 OA211x2_ASAP7_75t_R _20242_ (.A1(net408),
    .A2(_14132_),
    .B(_14917_),
    .C(net422),
    .Y(_14918_));
 OR3x1_ASAP7_75t_R _20243_ (.A(net385),
    .B(_14916_),
    .C(_14918_),
    .Y(_14919_));
 OA211x2_ASAP7_75t_R _20244_ (.A1(net320),
    .A2(_14914_),
    .B(_14919_),
    .C(_14780_),
    .Y(_14920_));
 AO221x2_ASAP7_75t_R _20245_ (.A1(net380),
    .A2(_14893_),
    .B1(_14906_),
    .B2(_14907_),
    .C(_14920_),
    .Y(_14921_));
 OA21x2_ASAP7_75t_R _20246_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_13808_),
    .B(_13794_),
    .Y(_14922_));
 OAI21x1_ASAP7_75t_R _20247_ (.A1(_13993_),
    .A2(_14921_),
    .B(_14922_),
    .Y(_14923_));
 NAND2x2_ASAP7_75t_R _20248_ (.A(_14854_),
    .B(_14923_),
    .Y(_18335_));
 INVx2_ASAP7_75t_R _20249_ (.A(_18335_),
    .Y(_18336_));
 XNOR2x1_ASAP7_75t_R _20250_ (.B(_14239_),
    .Y(_14924_),
    .A(_13620_));
 INVx1_ASAP7_75t_R _20251_ (.A(_00391_),
    .Y(_14925_));
 NAND2x1_ASAP7_75t_R _20252_ (.A(net392),
    .B(_00389_),
    .Y(_14926_));
 OA211x2_ASAP7_75t_R _20253_ (.A1(net392),
    .A2(_14925_),
    .B(_14926_),
    .C(_13649_),
    .Y(_14927_));
 INVx1_ASAP7_75t_R _20254_ (.A(_00390_),
    .Y(_14928_));
 NAND2x1_ASAP7_75t_R _20255_ (.A(net392),
    .B(_00388_),
    .Y(_14929_));
 OA211x2_ASAP7_75t_R _20256_ (.A1(net392),
    .A2(_14928_),
    .B(_14929_),
    .C(net419),
    .Y(_14930_));
 OR3x1_ASAP7_75t_R _20257_ (.A(_13636_),
    .B(_14927_),
    .C(_14930_),
    .Y(_14931_));
 NAND2x1_ASAP7_75t_R _20258_ (.A(net392),
    .B(_00397_),
    .Y(_14932_));
 OA211x2_ASAP7_75t_R _20259_ (.A1(net392),
    .A2(_14211_),
    .B(_14932_),
    .C(_13649_),
    .Y(_14933_));
 INVx1_ASAP7_75t_R _20260_ (.A(_00398_),
    .Y(_14934_));
 NAND2x1_ASAP7_75t_R _20261_ (.A(net392),
    .B(_00396_),
    .Y(_14935_));
 OA211x2_ASAP7_75t_R _20262_ (.A1(net392),
    .A2(_14934_),
    .B(_14935_),
    .C(net419),
    .Y(_14936_));
 OR3x1_ASAP7_75t_R _20263_ (.A(net381),
    .B(_14933_),
    .C(_14936_),
    .Y(_14937_));
 AO21x1_ASAP7_75t_R _20264_ (.A1(_14931_),
    .A2(_14937_),
    .B(net388),
    .Y(_14938_));
 AND2x2_ASAP7_75t_R _20265_ (.A(net393),
    .B(_01706_),
    .Y(_14939_));
 AO21x1_ASAP7_75t_R _20266_ (.A1(_13675_),
    .A2(_00387_),
    .B(_14939_),
    .Y(_14940_));
 OAI22x1_ASAP7_75t_R _20267_ (.A1(_00386_),
    .A2(net2291),
    .B1(_14940_),
    .B2(net427),
    .Y(_14941_));
 NAND2x2_ASAP7_75t_R _20268_ (.A(net387),
    .B(_13636_),
    .Y(_14942_));
 NAND2x1_ASAP7_75t_R _20269_ (.A(net393),
    .B(_00393_),
    .Y(_14943_));
 BUFx16f_ASAP7_75t_R input148 (.A(net2389),
    .Y(net148));
 OA211x2_ASAP7_75t_R _20271_ (.A1(net393),
    .A2(_14208_),
    .B(_14943_),
    .C(_13649_),
    .Y(_14945_));
 NAND2x1_ASAP7_75t_R _20272_ (.A(net393),
    .B(_00392_),
    .Y(_14946_));
 BUFx2_ASAP7_75t_R input147 (.A(net3206),
    .Y(net147));
 OA211x2_ASAP7_75t_R _20274_ (.A1(net393),
    .A2(_14214_),
    .B(_14946_),
    .C(net427),
    .Y(_14948_));
 OR3x1_ASAP7_75t_R _20275_ (.A(_14942_),
    .B(_14945_),
    .C(_14948_),
    .Y(_14949_));
 OA211x2_ASAP7_75t_R _20276_ (.A1(net315),
    .A2(_14941_),
    .B(_14949_),
    .C(_00286_),
    .Y(_14950_));
 BUFx2_ASAP7_75t_R input146 (.A(net3512),
    .Y(net146));
 INVx1_ASAP7_75t_R _20278_ (.A(_00411_),
    .Y(_14952_));
 BUFx3_ASAP7_75t_R input145 (.A(net3756),
    .Y(net145));
 NAND2x1_ASAP7_75t_R _20280_ (.A(net390),
    .B(_00409_),
    .Y(_14954_));
 OA211x2_ASAP7_75t_R _20281_ (.A1(net390),
    .A2(_14952_),
    .B(_14954_),
    .C(_13649_),
    .Y(_14955_));
 INVx1_ASAP7_75t_R _20282_ (.A(_00410_),
    .Y(_14956_));
 NAND2x1_ASAP7_75t_R _20283_ (.A(net390),
    .B(_00408_),
    .Y(_14957_));
 OA211x2_ASAP7_75t_R _20284_ (.A1(net390),
    .A2(_14956_),
    .B(_14957_),
    .C(net427),
    .Y(_14958_));
 OR3x1_ASAP7_75t_R _20285_ (.A(_13630_),
    .B(_14955_),
    .C(_14958_),
    .Y(_14959_));
 INVx1_ASAP7_75t_R _20286_ (.A(_00415_),
    .Y(_14960_));
 NAND2x1_ASAP7_75t_R _20287_ (.A(net392),
    .B(_00413_),
    .Y(_14961_));
 OA211x2_ASAP7_75t_R _20288_ (.A1(net392),
    .A2(_14960_),
    .B(_14961_),
    .C(_13649_),
    .Y(_14962_));
 INVx1_ASAP7_75t_R _20289_ (.A(_00414_),
    .Y(_14963_));
 NAND2x1_ASAP7_75t_R _20290_ (.A(net392),
    .B(_00412_),
    .Y(_14964_));
 OA211x2_ASAP7_75t_R _20291_ (.A1(net392),
    .A2(_14963_),
    .B(_14964_),
    .C(net419),
    .Y(_14965_));
 OR3x1_ASAP7_75t_R _20292_ (.A(net388),
    .B(_14962_),
    .C(_14965_),
    .Y(_14966_));
 AO21x1_ASAP7_75t_R _20293_ (.A1(_14959_),
    .A2(_14966_),
    .B(net381),
    .Y(_14967_));
 NAND2x1_ASAP7_75t_R _20294_ (.A(net416),
    .B(_00405_),
    .Y(_14968_));
 OA211x2_ASAP7_75t_R _20295_ (.A1(net416),
    .A2(_14200_),
    .B(_14968_),
    .C(net319),
    .Y(_14969_));
 INVx1_ASAP7_75t_R _20296_ (.A(_00406_),
    .Y(_14970_));
 NAND2x1_ASAP7_75t_R _20297_ (.A(net417),
    .B(_00404_),
    .Y(_14971_));
 OA211x2_ASAP7_75t_R _20298_ (.A1(net417),
    .A2(_14970_),
    .B(_14971_),
    .C(net426),
    .Y(_14972_));
 OR3x1_ASAP7_75t_R _20299_ (.A(_14015_),
    .B(_14969_),
    .C(_14972_),
    .Y(_14973_));
 NAND2x1_ASAP7_75t_R _20300_ (.A(net417),
    .B(_00401_),
    .Y(_14974_));
 OA211x2_ASAP7_75t_R _20301_ (.A1(net417),
    .A2(_14194_),
    .B(_14974_),
    .C(net319),
    .Y(_14975_));
 NAND2x1_ASAP7_75t_R _20302_ (.A(net417),
    .B(_00400_),
    .Y(_14976_));
 OA211x2_ASAP7_75t_R _20303_ (.A1(net417),
    .A2(_14197_),
    .B(_14976_),
    .C(net426),
    .Y(_14977_));
 OR3x1_ASAP7_75t_R _20304_ (.A(net315),
    .B(_14975_),
    .C(_14977_),
    .Y(_14978_));
 AND3x1_ASAP7_75t_R _20305_ (.A(_13626_),
    .B(_14973_),
    .C(_14978_),
    .Y(_14979_));
 AO22x2_ASAP7_75t_R _20306_ (.A1(_14938_),
    .A2(_14950_),
    .B1(_14967_),
    .B2(_14979_),
    .Y(_14980_));
 BUFx2_ASAP7_75t_R input144 (.A(net3663),
    .Y(net144));
 AOI22x1_ASAP7_75t_R _20308_ (.A1(_13775_),
    .A2(_00665_),
    .B1(_01449_),
    .B2(_13778_),
    .Y(_14982_));
 OA211x2_ASAP7_75t_R _20309_ (.A1(_00284_),
    .A2(_14980_),
    .B(_14982_),
    .C(_13986_),
    .Y(_14983_));
 BUFx2_ASAP7_75t_R input143 (.A(net3547),
    .Y(net143));
 AOI211x1_ASAP7_75t_R _20311_ (.A1(_13772_),
    .A2(net2230),
    .B(_14983_),
    .C(_13538_),
    .Y(_14985_));
 AO21x1_ASAP7_75t_R _20312_ (.A1(_13538_),
    .A2(_14924_),
    .B(_14985_),
    .Y(_17760_));
 INVx1_ASAP7_75t_R _20313_ (.A(_17760_),
    .Y(_16723_));
 INVx1_ASAP7_75t_R _20314_ (.A(_00170_),
    .Y(\cs_registers_i.pc_id_i[3] ));
 AO21x1_ASAP7_75t_R _20315_ (.A1(_13445_),
    .A2(_13449_),
    .B(_01638_),
    .Y(_14986_));
 OA31x2_ASAP7_75t_R _20316_ (.A1(_00287_),
    .A2(_13784_),
    .A3(_13808_),
    .B1(_14986_),
    .Y(_14987_));
 AO221x2_ASAP7_75t_R _20317_ (.A1(_13570_),
    .A2(_13785_),
    .B1(_13788_),
    .B2(_13792_),
    .C(_13793_),
    .Y(_14988_));
 BUFx2_ASAP7_75t_R input142 (.A(net3491),
    .Y(net142));
 AND2x2_ASAP7_75t_R _20319_ (.A(_00170_),
    .B(_13993_),
    .Y(_14990_));
 AOI221x1_ASAP7_75t_R _20320_ (.A1(_14938_),
    .A2(_14950_),
    .B1(_14967_),
    .B2(_14979_),
    .C(_13993_),
    .Y(_14991_));
 OR3x4_ASAP7_75t_R _20321_ (.A(_14988_),
    .B(_14990_),
    .C(_14991_),
    .Y(_14992_));
 NAND2x2_ASAP7_75t_R _20322_ (.A(_14987_),
    .B(_14992_),
    .Y(_18341_));
 INVx3_ASAP7_75t_R _20323_ (.A(_18341_),
    .Y(_18339_));
 OAI21x1_ASAP7_75t_R _20324_ (.A1(_00665_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_14993_));
 OA21x2_ASAP7_75t_R _20325_ (.A1(_13817_),
    .A2(_18341_),
    .B(_14993_),
    .Y(_17761_));
 INVx1_ASAP7_75t_R _20326_ (.A(_17761_),
    .Y(_16724_));
 INVx1_ASAP7_75t_R _20327_ (.A(_17757_),
    .Y(_16714_));
 OA21x2_ASAP7_75t_R _20328_ (.A1(_00292_),
    .A2(_16714_),
    .B(_00664_),
    .Y(_14994_));
 OA21x2_ASAP7_75t_R _20329_ (.A1(_02262_),
    .A2(_14994_),
    .B(_00667_),
    .Y(_16722_));
 INVx1_ASAP7_75t_R _20330_ (.A(_00437_),
    .Y(_14995_));
 BUFx2_ASAP7_75t_R input141 (.A(net3565),
    .Y(net141));
 NAND2x1_ASAP7_75t_R _20332_ (.A(net405),
    .B(_00435_),
    .Y(_14997_));
 OA211x2_ASAP7_75t_R _20333_ (.A1(net405),
    .A2(_14995_),
    .B(_14997_),
    .C(net318),
    .Y(_14998_));
 NAND2x1_ASAP7_75t_R _20334_ (.A(net405),
    .B(_00434_),
    .Y(_14999_));
 OA211x2_ASAP7_75t_R _20335_ (.A1(net405),
    .A2(_14264_),
    .B(_14999_),
    .C(net420),
    .Y(_15000_));
 OR3x1_ASAP7_75t_R _20336_ (.A(net384),
    .B(_14998_),
    .C(_15000_),
    .Y(_15001_));
 INVx1_ASAP7_75t_R _20337_ (.A(_00433_),
    .Y(_15002_));
 NAND2x1_ASAP7_75t_R _20338_ (.A(net2377),
    .B(_00431_),
    .Y(_15003_));
 OA211x2_ASAP7_75t_R _20339_ (.A1(net2352),
    .A2(_15002_),
    .B(_15003_),
    .C(net318),
    .Y(_15004_));
 BUFx2_ASAP7_75t_R input140 (.A(net3532),
    .Y(net140));
 NAND2x1_ASAP7_75t_R _20341_ (.A(net405),
    .B(_00430_),
    .Y(_15006_));
 OA211x2_ASAP7_75t_R _20342_ (.A1(net405),
    .A2(_14267_),
    .B(_15006_),
    .C(net420),
    .Y(_15007_));
 OR3x1_ASAP7_75t_R _20343_ (.A(net320),
    .B(_15004_),
    .C(_15007_),
    .Y(_15008_));
 INVx1_ASAP7_75t_R _20344_ (.A(_00421_),
    .Y(_15009_));
 BUFx2_ASAP7_75t_R input139 (.A(net3496),
    .Y(net139));
 NAND2x1_ASAP7_75t_R _20346_ (.A(net2377),
    .B(_00419_),
    .Y(_15011_));
 OA211x2_ASAP7_75t_R _20347_ (.A1(net2352),
    .A2(_15009_),
    .B(_15011_),
    .C(net317),
    .Y(_15012_));
 INVx1_ASAP7_75t_R _20348_ (.A(_00420_),
    .Y(_15013_));
 NAND2x1_ASAP7_75t_R _20349_ (.A(net2377),
    .B(_00418_),
    .Y(_15014_));
 OA211x2_ASAP7_75t_R _20350_ (.A1(net2352),
    .A2(_15013_),
    .B(_15014_),
    .C(net420),
    .Y(_15015_));
 OR3x1_ASAP7_75t_R _20351_ (.A(net312),
    .B(_15012_),
    .C(_15015_),
    .Y(_15016_));
 NAND2x1_ASAP7_75t_R _20352_ (.A(net2352),
    .B(_01705_),
    .Y(_15017_));
 OA211x2_ASAP7_75t_R _20353_ (.A1(net2352),
    .A2(_14259_),
    .B(_15017_),
    .C(net317),
    .Y(_15018_));
 AND3x1_ASAP7_75t_R _20354_ (.A(net420),
    .B(net316),
    .C(_14258_),
    .Y(_15019_));
 OA31x2_ASAP7_75t_R _20355_ (.A1(_14005_),
    .A2(_15018_),
    .A3(_15019_),
    .B1(net377),
    .Y(_15020_));
 AO32x1_ASAP7_75t_R _20356_ (.A1(_13626_),
    .A2(_15001_),
    .A3(_15008_),
    .B1(_15016_),
    .B2(_15020_),
    .Y(_15021_));
 BUFx2_ASAP7_75t_R input138 (.A(net3703),
    .Y(net138));
 NAND2x1_ASAP7_75t_R _20358_ (.A(net402),
    .B(_00427_),
    .Y(_15023_));
 OA211x2_ASAP7_75t_R _20359_ (.A1(net2376),
    .A2(_14249_),
    .B(_15023_),
    .C(net317),
    .Y(_15024_));
 NAND2x1_ASAP7_75t_R _20360_ (.A(net402),
    .B(_00426_),
    .Y(_15025_));
 BUFx2_ASAP7_75t_R input137 (.A(net3577),
    .Y(net137));
 OA211x2_ASAP7_75t_R _20362_ (.A1(net2376),
    .A2(_14241_),
    .B(_15025_),
    .C(net420),
    .Y(_15027_));
 OR3x1_ASAP7_75t_R _20363_ (.A(net384),
    .B(_15024_),
    .C(_15027_),
    .Y(_15028_));
 INVx1_ASAP7_75t_R _20364_ (.A(_00425_),
    .Y(_15029_));
 NAND2x1_ASAP7_75t_R _20365_ (.A(net403),
    .B(_00423_),
    .Y(_15030_));
 OA211x2_ASAP7_75t_R _20366_ (.A1(net403),
    .A2(_15029_),
    .B(_15030_),
    .C(net317),
    .Y(_15031_));
 INVx1_ASAP7_75t_R _20367_ (.A(_00424_),
    .Y(_15032_));
 NAND2x1_ASAP7_75t_R _20368_ (.A(net403),
    .B(_00422_),
    .Y(_15033_));
 OA211x2_ASAP7_75t_R _20369_ (.A1(net403),
    .A2(_15032_),
    .B(_15033_),
    .C(net420),
    .Y(_15034_));
 OR3x1_ASAP7_75t_R _20370_ (.A(net320),
    .B(_15031_),
    .C(_15034_),
    .Y(_15035_));
 AND2x2_ASAP7_75t_R _20371_ (.A(_15028_),
    .B(_15035_),
    .Y(_15036_));
 AND2x2_ASAP7_75t_R _20372_ (.A(_15016_),
    .B(_15020_),
    .Y(_15037_));
 INVx1_ASAP7_75t_R _20373_ (.A(_00441_),
    .Y(_15038_));
 NAND2x1_ASAP7_75t_R _20374_ (.A(net400),
    .B(_00439_),
    .Y(_15039_));
 OA211x2_ASAP7_75t_R _20375_ (.A1(net400),
    .A2(_15038_),
    .B(_15039_),
    .C(net318),
    .Y(_15040_));
 NAND2x1_ASAP7_75t_R _20376_ (.A(net400),
    .B(_00438_),
    .Y(_15041_));
 OA211x2_ASAP7_75t_R _20377_ (.A1(net400),
    .A2(_14280_),
    .B(_15041_),
    .C(net421),
    .Y(_15042_));
 OR3x1_ASAP7_75t_R _20378_ (.A(net320),
    .B(_15040_),
    .C(_15042_),
    .Y(_15043_));
 NAND2x1_ASAP7_75t_R _20379_ (.A(net2352),
    .B(_00443_),
    .Y(_15044_));
 OA211x2_ASAP7_75t_R _20380_ (.A1(net2352),
    .A2(_14286_),
    .B(_15044_),
    .C(net318),
    .Y(_15045_));
 NAND2x1_ASAP7_75t_R _20381_ (.A(net2352),
    .B(_00442_),
    .Y(_15046_));
 OA211x2_ASAP7_75t_R _20382_ (.A1(net2352),
    .A2(_14283_),
    .B(_15046_),
    .C(net420),
    .Y(_15047_));
 OR3x1_ASAP7_75t_R _20383_ (.A(net384),
    .B(_15045_),
    .C(_15047_),
    .Y(_15048_));
 AND3x1_ASAP7_75t_R _20384_ (.A(_14780_),
    .B(_15043_),
    .C(_15048_),
    .Y(_15049_));
 AO221x2_ASAP7_75t_R _20385_ (.A1(net380),
    .A2(_15021_),
    .B1(_15036_),
    .B2(_15037_),
    .C(_15049_),
    .Y(_15050_));
 INVx1_ASAP7_75t_R _20386_ (.A(_00174_),
    .Y(_15051_));
 AND3x2_ASAP7_75t_R _20387_ (.A(_15051_),
    .B(_13993_),
    .C(_13794_),
    .Y(_15052_));
 INVx1_ASAP7_75t_R _20388_ (.A(_01637_),
    .Y(_15053_));
 AO32x1_ASAP7_75t_R _20389_ (.A1(_13626_),
    .A2(_13802_),
    .A3(_13993_),
    .B1(_15053_),
    .B2(_13450_),
    .Y(_15054_));
 AOI211x1_ASAP7_75t_R _20390_ (.A1(_13810_),
    .A2(net2322),
    .B(_15052_),
    .C(_15054_),
    .Y(_18344_));
 NAND2x1_ASAP7_75t_R _20391_ (.A(net403),
    .B(_00460_),
    .Y(_15055_));
 OA211x2_ASAP7_75t_R _20392_ (.A1(net403),
    .A2(_14312_),
    .B(_15055_),
    .C(net384),
    .Y(_15056_));
 NAND2x1_ASAP7_75t_R _20393_ (.A(net404),
    .B(_00464_),
    .Y(_15057_));
 OA211x2_ASAP7_75t_R _20394_ (.A1(net404),
    .A2(_14309_),
    .B(_15057_),
    .C(net320),
    .Y(_15058_));
 OR3x1_ASAP7_75t_R _20395_ (.A(net317),
    .B(_15056_),
    .C(_15058_),
    .Y(_15059_));
 NAND2x1_ASAP7_75t_R _20396_ (.A(net404),
    .B(_00461_),
    .Y(_15060_));
 OA211x2_ASAP7_75t_R _20397_ (.A1(net404),
    .A2(_14301_),
    .B(_15060_),
    .C(net384),
    .Y(_15061_));
 NAND2x1_ASAP7_75t_R _20398_ (.A(net404),
    .B(_00465_),
    .Y(_15062_));
 OA211x2_ASAP7_75t_R _20399_ (.A1(net404),
    .A2(_14305_),
    .B(_15062_),
    .C(net320),
    .Y(_15063_));
 OR3x1_ASAP7_75t_R _20400_ (.A(net420),
    .B(_15061_),
    .C(_15063_),
    .Y(_15064_));
 INVx1_ASAP7_75t_R _20401_ (.A(_00450_),
    .Y(_15065_));
 BUFx2_ASAP7_75t_R input136 (.A(net3664),
    .Y(net136));
 NAND2x1_ASAP7_75t_R _20403_ (.A(net404),
    .B(_00448_),
    .Y(_15067_));
 OA211x2_ASAP7_75t_R _20404_ (.A1(net404),
    .A2(_15065_),
    .B(_15067_),
    .C(net420),
    .Y(_15068_));
 INVx1_ASAP7_75t_R _20405_ (.A(_00451_),
    .Y(_15069_));
 NAND2x1_ASAP7_75t_R _20406_ (.A(net404),
    .B(_00449_),
    .Y(_15070_));
 OA211x2_ASAP7_75t_R _20407_ (.A1(net404),
    .A2(_15069_),
    .B(_15070_),
    .C(net317),
    .Y(_15071_));
 OR3x1_ASAP7_75t_R _20408_ (.A(net312),
    .B(_15068_),
    .C(_15071_),
    .Y(_15072_));
 NAND2x1_ASAP7_75t_R _20409_ (.A(net405),
    .B(_01704_),
    .Y(_15073_));
 OA211x2_ASAP7_75t_R _20410_ (.A1(net405),
    .A2(_14350_),
    .B(_15073_),
    .C(net318),
    .Y(_15074_));
 AND3x1_ASAP7_75t_R _20411_ (.A(net420),
    .B(net316),
    .C(_14349_),
    .Y(_15075_));
 OA31x2_ASAP7_75t_R _20412_ (.A1(_14005_),
    .A2(_15074_),
    .A3(_15075_),
    .B1(net377),
    .Y(_15076_));
 AO32x1_ASAP7_75t_R _20413_ (.A1(_13626_),
    .A2(_15059_),
    .A3(_15064_),
    .B1(_15072_),
    .B2(_15076_),
    .Y(_15077_));
 BUFx2_ASAP7_75t_R input135 (.A(net3485),
    .Y(net135));
 NAND2x1_ASAP7_75t_R _20415_ (.A(net402),
    .B(_00457_),
    .Y(_15079_));
 OA211x2_ASAP7_75t_R _20416_ (.A1(net2376),
    .A2(_14337_),
    .B(_15079_),
    .C(net317),
    .Y(_15080_));
 NAND2x1_ASAP7_75t_R _20417_ (.A(net402),
    .B(_00456_),
    .Y(_15081_));
 OA211x2_ASAP7_75t_R _20418_ (.A1(net2376),
    .A2(_14330_),
    .B(_15081_),
    .C(net420),
    .Y(_15082_));
 OR3x1_ASAP7_75t_R _20419_ (.A(net384),
    .B(_15080_),
    .C(_15082_),
    .Y(_15083_));
 BUFx2_ASAP7_75t_R input134 (.A(net3386),
    .Y(net134));
 NAND2x1_ASAP7_75t_R _20421_ (.A(net402),
    .B(_00453_),
    .Y(_15085_));
 OA211x2_ASAP7_75t_R _20422_ (.A1(net2376),
    .A2(_14340_),
    .B(_15085_),
    .C(net317),
    .Y(_15086_));
 NAND2x1_ASAP7_75t_R _20423_ (.A(net402),
    .B(_00452_),
    .Y(_15087_));
 OA211x2_ASAP7_75t_R _20424_ (.A1(net2376),
    .A2(_14333_),
    .B(_15087_),
    .C(net420),
    .Y(_15088_));
 OR3x1_ASAP7_75t_R _20425_ (.A(net320),
    .B(_15086_),
    .C(_15088_),
    .Y(_15089_));
 AND2x2_ASAP7_75t_R _20426_ (.A(_15083_),
    .B(_15089_),
    .Y(_15090_));
 AND2x2_ASAP7_75t_R _20427_ (.A(_15072_),
    .B(_15076_),
    .Y(_15091_));
 NAND2x1_ASAP7_75t_R _20428_ (.A(net403),
    .B(_00473_),
    .Y(_15092_));
 OA211x2_ASAP7_75t_R _20429_ (.A1(net2376),
    .A2(_14319_),
    .B(_15092_),
    .C(net317),
    .Y(_15093_));
 NAND2x1_ASAP7_75t_R _20430_ (.A(net402),
    .B(_00472_),
    .Y(_15094_));
 OA211x2_ASAP7_75t_R _20431_ (.A1(net2376),
    .A2(_14325_),
    .B(_15094_),
    .C(net420),
    .Y(_15095_));
 OR3x1_ASAP7_75t_R _20432_ (.A(net384),
    .B(_15093_),
    .C(_15095_),
    .Y(_15096_));
 NAND2x1_ASAP7_75t_R _20433_ (.A(net402),
    .B(_00469_),
    .Y(_15097_));
 OA211x2_ASAP7_75t_R _20434_ (.A1(net2376),
    .A2(_14316_),
    .B(_15097_),
    .C(net318),
    .Y(_15098_));
 NAND2x1_ASAP7_75t_R _20435_ (.A(net402),
    .B(_00468_),
    .Y(_15099_));
 OA211x2_ASAP7_75t_R _20436_ (.A1(net2376),
    .A2(_14322_),
    .B(_15099_),
    .C(net420),
    .Y(_15100_));
 OR3x1_ASAP7_75t_R _20437_ (.A(net320),
    .B(_15098_),
    .C(_15100_),
    .Y(_15101_));
 AND3x1_ASAP7_75t_R _20438_ (.A(_14780_),
    .B(_15096_),
    .C(_15101_),
    .Y(_15102_));
 AO221x2_ASAP7_75t_R _20439_ (.A1(net380),
    .A2(_15077_),
    .B1(_15090_),
    .B2(_15091_),
    .C(_15102_),
    .Y(_15103_));
 BUFx2_ASAP7_75t_R input133 (.A(net3549),
    .Y(net133));
 INVx1_ASAP7_75t_R _20441_ (.A(_00670_),
    .Y(_15105_));
 INVx1_ASAP7_75t_R _20442_ (.A(_01447_),
    .Y(_15106_));
 BUFx2_ASAP7_75t_R input132 (.A(net3538),
    .Y(net132));
 OA222x2_ASAP7_75t_R _20444_ (.A1(_00285_),
    .A2(_15105_),
    .B1(_15106_),
    .B2(_13815_),
    .C1(_13986_),
    .C2(_14355_),
    .Y(_15108_));
 OA21x2_ASAP7_75t_R _20445_ (.A1(_00284_),
    .A2(_15103_),
    .B(_15108_),
    .Y(_15109_));
 XNOR2x1_ASAP7_75t_R _20446_ (.B(_14359_),
    .Y(_15110_),
    .A(_13620_));
 AND2x2_ASAP7_75t_R _20447_ (.A(net309),
    .B(_15110_),
    .Y(_15111_));
 AOI21x1_ASAP7_75t_R _20448_ (.A1(_13817_),
    .A2(_15109_),
    .B(_15111_),
    .Y(_17764_));
 INVx1_ASAP7_75t_R _20449_ (.A(_17764_),
    .Y(_16725_));
 INVx2_ASAP7_75t_R _20450_ (.A(_00177_),
    .Y(\cs_registers_i.pc_id_i[5] ));
 NAND2x2_ASAP7_75t_R _20451_ (.A(_13808_),
    .B(_13794_),
    .Y(_15112_));
 NOR2x1_ASAP7_75t_R _20452_ (.A(_01636_),
    .B(_13807_),
    .Y(_15113_));
 OA21x2_ASAP7_75t_R _20453_ (.A1(\cs_registers_i.pc_id_i[5] ),
    .A2(_13808_),
    .B(_13794_),
    .Y(_15114_));
 OA22x2_ASAP7_75t_R _20454_ (.A1(_15112_),
    .A2(_15103_),
    .B1(_15113_),
    .B2(_15114_),
    .Y(_15115_));
 BUFx2_ASAP7_75t_R input131 (.A(net3406),
    .Y(net131));
 INVx3_ASAP7_75t_R _20456_ (.A(_15115_),
    .Y(_18351_));
 OR3x1_ASAP7_75t_R _20457_ (.A(_00670_),
    .B(net309),
    .C(_13815_),
    .Y(_15116_));
 OAI21x1_ASAP7_75t_R _20458_ (.A1(_13817_),
    .A2(_18351_),
    .B(_15116_),
    .Y(_17765_));
 INVx1_ASAP7_75t_R _20459_ (.A(_17765_),
    .Y(_16726_));
 OR2x2_ASAP7_75t_R _20460_ (.A(_00666_),
    .B(_02264_),
    .Y(_15117_));
 OA21x2_ASAP7_75t_R _20461_ (.A1(_00667_),
    .A2(_00666_),
    .B(_00669_),
    .Y(_15118_));
 OA21x2_ASAP7_75t_R _20462_ (.A1(_02264_),
    .A2(_15118_),
    .B(_02263_),
    .Y(_15119_));
 OA31x2_ASAP7_75t_R _20463_ (.A1(_02262_),
    .A2(_14994_),
    .A3(_15117_),
    .B1(_15119_),
    .Y(_16727_));
 NAND2x1_ASAP7_75t_R _20464_ (.A(net408),
    .B(_00495_),
    .Y(_15120_));
 OA211x2_ASAP7_75t_R _20465_ (.A1(net408),
    .A2(_14398_),
    .B(_15120_),
    .C(net318),
    .Y(_15121_));
 NAND2x1_ASAP7_75t_R _20466_ (.A(net2377),
    .B(_00494_),
    .Y(_15122_));
 OA211x2_ASAP7_75t_R _20467_ (.A1(net406),
    .A2(_14395_),
    .B(_15122_),
    .C(net422),
    .Y(_15123_));
 OR3x1_ASAP7_75t_R _20468_ (.A(net312),
    .B(_15121_),
    .C(_15123_),
    .Y(_15124_));
 INVx1_ASAP7_75t_R _20469_ (.A(_00493_),
    .Y(_15125_));
 NAND2x1_ASAP7_75t_R _20470_ (.A(net2377),
    .B(_00491_),
    .Y(_15126_));
 OA211x2_ASAP7_75t_R _20471_ (.A1(net406),
    .A2(_15125_),
    .B(_15126_),
    .C(net318),
    .Y(_15127_));
 INVx1_ASAP7_75t_R _20472_ (.A(_00492_),
    .Y(_15128_));
 NAND2x1_ASAP7_75t_R _20473_ (.A(net2377),
    .B(_00490_),
    .Y(_15129_));
 OA211x2_ASAP7_75t_R _20474_ (.A1(net406),
    .A2(_15128_),
    .B(_15129_),
    .C(net422),
    .Y(_15130_));
 OR3x1_ASAP7_75t_R _20475_ (.A(_14005_),
    .B(_15127_),
    .C(_15130_),
    .Y(_15131_));
 AND3x1_ASAP7_75t_R _20476_ (.A(_13626_),
    .B(_15124_),
    .C(_15131_),
    .Y(_15132_));
 OR2x2_ASAP7_75t_R _20477_ (.A(net408),
    .B(_00504_),
    .Y(_15133_));
 OAI21x1_ASAP7_75t_R _20478_ (.A1(net316),
    .A2(_00502_),
    .B(_15133_),
    .Y(_15134_));
 INVx1_ASAP7_75t_R _20479_ (.A(_00505_),
    .Y(_15135_));
 NAND2x1_ASAP7_75t_R _20480_ (.A(net408),
    .B(_00503_),
    .Y(_15136_));
 OA211x2_ASAP7_75t_R _20481_ (.A1(net408),
    .A2(_15135_),
    .B(_15136_),
    .C(net318),
    .Y(_15137_));
 AO21x1_ASAP7_75t_R _20482_ (.A1(net422),
    .A2(_15134_),
    .B(_15137_),
    .Y(_15138_));
 NAND2x1_ASAP7_75t_R _20483_ (.A(net408),
    .B(_00499_),
    .Y(_15139_));
 OA211x2_ASAP7_75t_R _20484_ (.A1(net408),
    .A2(_14412_),
    .B(_15139_),
    .C(net318),
    .Y(_15140_));
 NAND2x1_ASAP7_75t_R _20485_ (.A(net408),
    .B(_00498_),
    .Y(_15141_));
 OA211x2_ASAP7_75t_R _20486_ (.A1(net408),
    .A2(_14415_),
    .B(_15141_),
    .C(net422),
    .Y(_15142_));
 OR3x1_ASAP7_75t_R _20487_ (.A(net320),
    .B(_15140_),
    .C(_15142_),
    .Y(_15143_));
 OA21x2_ASAP7_75t_R _20488_ (.A1(net384),
    .A2(_15138_),
    .B(_15143_),
    .Y(_15144_));
 NAND2x1_ASAP7_75t_R _20489_ (.A(net408),
    .B(_00478_),
    .Y(_15145_));
 OA211x2_ASAP7_75t_R _20490_ (.A1(net408),
    .A2(_14380_),
    .B(_15145_),
    .C(net422),
    .Y(_15146_));
 NAND2x1_ASAP7_75t_R _20491_ (.A(net408),
    .B(_00479_),
    .Y(_15147_));
 OA211x2_ASAP7_75t_R _20492_ (.A1(net408),
    .A2(_14384_),
    .B(_15147_),
    .C(net318),
    .Y(_15148_));
 OR3x1_ASAP7_75t_R _20493_ (.A(net312),
    .B(_15146_),
    .C(_15148_),
    .Y(_15149_));
 NAND2x1_ASAP7_75t_R _20494_ (.A(net405),
    .B(_01703_),
    .Y(_15150_));
 OA211x2_ASAP7_75t_R _20495_ (.A1(net405),
    .A2(_14390_),
    .B(_15150_),
    .C(net318),
    .Y(_15151_));
 AND3x1_ASAP7_75t_R _20496_ (.A(net422),
    .B(net316),
    .C(_14388_),
    .Y(_15152_));
 OA31x2_ASAP7_75t_R _20497_ (.A1(_14005_),
    .A2(_15151_),
    .A3(_15152_),
    .B1(net377),
    .Y(_15153_));
 AO32x1_ASAP7_75t_R _20498_ (.A1(_13626_),
    .A2(_15124_),
    .A3(_15131_),
    .B1(_15149_),
    .B2(_15153_),
    .Y(_15154_));
 NAND2x1_ASAP7_75t_R _20499_ (.A(net2369),
    .B(_00487_),
    .Y(_15155_));
 OA211x2_ASAP7_75t_R _20500_ (.A1(net2369),
    .A2(_14373_),
    .B(_15155_),
    .C(net318),
    .Y(_15156_));
 NAND2x1_ASAP7_75t_R _20501_ (.A(net2369),
    .B(_00486_),
    .Y(_15157_));
 OA211x2_ASAP7_75t_R _20502_ (.A1(net2369),
    .A2(_14366_),
    .B(_15157_),
    .C(net422),
    .Y(_15158_));
 OR3x1_ASAP7_75t_R _20503_ (.A(net384),
    .B(_15156_),
    .C(_15158_),
    .Y(_15159_));
 INVx1_ASAP7_75t_R _20504_ (.A(_00485_),
    .Y(_15160_));
 NAND2x1_ASAP7_75t_R _20505_ (.A(net2369),
    .B(_00483_),
    .Y(_15161_));
 OA211x2_ASAP7_75t_R _20506_ (.A1(net2369),
    .A2(_15160_),
    .B(_15161_),
    .C(net318),
    .Y(_15162_));
 NAND2x1_ASAP7_75t_R _20507_ (.A(net2369),
    .B(_00482_),
    .Y(_15163_));
 OA211x2_ASAP7_75t_R _20508_ (.A1(net2352),
    .A2(_14369_),
    .B(_15163_),
    .C(net422),
    .Y(_15164_));
 OR3x1_ASAP7_75t_R _20509_ (.A(net320),
    .B(_15162_),
    .C(_15164_),
    .Y(_15165_));
 AND4x1_ASAP7_75t_R _20510_ (.A(_15149_),
    .B(_15153_),
    .C(_15159_),
    .D(_15165_),
    .Y(_15166_));
 AO221x2_ASAP7_75t_R _20511_ (.A1(_15132_),
    .A2(_15144_),
    .B1(_15154_),
    .B2(net380),
    .C(_15166_),
    .Y(_15167_));
 BUFx2_ASAP7_75t_R input130 (.A(net3298),
    .Y(net130));
 INVx2_ASAP7_75t_R _20513_ (.A(_00180_),
    .Y(_15169_));
 INVx1_ASAP7_75t_R _20514_ (.A(_01635_),
    .Y(_15170_));
 AO32x2_ASAP7_75t_R _20515_ (.A1(_15169_),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_15170_),
    .B2(_13450_),
    .Y(_15171_));
 AO21x2_ASAP7_75t_R _20516_ (.A1(_13810_),
    .A2(_15167_),
    .B(_15171_),
    .Y(_15172_));
 BUFx2_ASAP7_75t_R input129 (.A(net3625),
    .Y(net129));
 INVx1_ASAP7_75t_R _20518_ (.A(_15172_),
    .Y(_18356_));
 INVx2_ASAP7_75t_R _20519_ (.A(_00182_),
    .Y(\cs_registers_i.pc_id_i[7] ));
 BUFx3_ASAP7_75t_R input128 (.A(net2972),
    .Y(net128));
 INVx1_ASAP7_75t_R _20521_ (.A(_00515_),
    .Y(_15174_));
 NAND2x1_ASAP7_75t_R _20522_ (.A(net2379),
    .B(_00513_),
    .Y(_15175_));
 BUFx2_ASAP7_75t_R input127 (.A(net2793),
    .Y(net127));
 OA211x2_ASAP7_75t_R _20524_ (.A1(net2379),
    .A2(_15174_),
    .B(_15175_),
    .C(net318),
    .Y(_15177_));
 NAND2x1_ASAP7_75t_R _20525_ (.A(net398),
    .B(_00512_),
    .Y(_15178_));
 OA211x2_ASAP7_75t_R _20526_ (.A1(net398),
    .A2(_14428_),
    .B(_15178_),
    .C(net425),
    .Y(_15179_));
 NAND2x1_ASAP7_75t_R _20527_ (.A(net2379),
    .B(_01702_),
    .Y(_15180_));
 OA211x2_ASAP7_75t_R _20528_ (.A1(net2379),
    .A2(_14448_),
    .B(_15180_),
    .C(net318),
    .Y(_15181_));
 AND3x1_ASAP7_75t_R _20529_ (.A(net425),
    .B(net316),
    .C(_14446_),
    .Y(_15182_));
 OA33x2_ASAP7_75t_R _20530_ (.A1(_14942_),
    .A2(_15177_),
    .A3(_15179_),
    .B1(_15181_),
    .B2(_15182_),
    .B3(net315),
    .Y(_15183_));
 NAND2x1_ASAP7_75t_R _20531_ (.A(net409),
    .B(_00509_),
    .Y(_15184_));
 OA211x2_ASAP7_75t_R _20532_ (.A1(net409),
    .A2(_14442_),
    .B(_15184_),
    .C(net318),
    .Y(_15185_));
 BUFx2_ASAP7_75t_R input126 (.A(net2982),
    .Y(net126));
 NAND2x1_ASAP7_75t_R _20534_ (.A(net2379),
    .B(_00508_),
    .Y(_15187_));
 OA211x2_ASAP7_75t_R _20535_ (.A1(net411),
    .A2(_14439_),
    .B(_15187_),
    .C(net425),
    .Y(_15188_));
 OR3x1_ASAP7_75t_R _20536_ (.A(_13636_),
    .B(_15185_),
    .C(_15188_),
    .Y(_15189_));
 NAND2x1_ASAP7_75t_R _20537_ (.A(net2379),
    .B(_00517_),
    .Y(_15190_));
 OA211x2_ASAP7_75t_R _20538_ (.A1(net411),
    .A2(_14432_),
    .B(_15190_),
    .C(net318),
    .Y(_15191_));
 NAND2x1_ASAP7_75t_R _20539_ (.A(net2379),
    .B(_00516_),
    .Y(_15192_));
 OA211x2_ASAP7_75t_R _20540_ (.A1(net411),
    .A2(_14425_),
    .B(_15192_),
    .C(net425),
    .Y(_15193_));
 OR3x1_ASAP7_75t_R _20541_ (.A(net380),
    .B(_15191_),
    .C(_15193_),
    .Y(_15194_));
 AO21x1_ASAP7_75t_R _20542_ (.A1(_15189_),
    .A2(_15194_),
    .B(net385),
    .Y(_15195_));
 AO21x1_ASAP7_75t_R _20543_ (.A1(_15183_),
    .A2(_15195_),
    .B(_13626_),
    .Y(_15196_));
 INVx1_ASAP7_75t_R _20544_ (.A(_00529_),
    .Y(_15197_));
 NAND2x1_ASAP7_75t_R _20545_ (.A(net425),
    .B(_00528_),
    .Y(_15198_));
 OA211x2_ASAP7_75t_R _20546_ (.A1(net425),
    .A2(_15197_),
    .B(_15198_),
    .C(net409),
    .Y(_15199_));
 AND2x2_ASAP7_75t_R _20547_ (.A(net425),
    .B(_00530_),
    .Y(_15200_));
 AO21x1_ASAP7_75t_R _20548_ (.A1(net318),
    .A2(_00531_),
    .B(_15200_),
    .Y(_15201_));
 OAI21x1_ASAP7_75t_R _20549_ (.A1(net409),
    .A2(_15201_),
    .B(net385),
    .Y(_15202_));
 NAND2x1_ASAP7_75t_R _20550_ (.A(net409),
    .B(_00533_),
    .Y(_15203_));
 OA211x2_ASAP7_75t_R _20551_ (.A1(net409),
    .A2(_14471_),
    .B(_15203_),
    .C(net318),
    .Y(_15204_));
 NAND2x1_ASAP7_75t_R _20552_ (.A(net409),
    .B(_00532_),
    .Y(_15205_));
 OA211x2_ASAP7_75t_R _20553_ (.A1(net409),
    .A2(_14474_),
    .B(_15205_),
    .C(net425),
    .Y(_15206_));
 OR3x1_ASAP7_75t_R _20554_ (.A(net385),
    .B(_15204_),
    .C(_15206_),
    .Y(_15207_));
 OA211x2_ASAP7_75t_R _20555_ (.A1(_15199_),
    .A2(_15202_),
    .B(_15207_),
    .C(_13636_),
    .Y(_15208_));
 NAND2x1_ASAP7_75t_R _20556_ (.A(net2379),
    .B(_00524_),
    .Y(_15209_));
 OA211x2_ASAP7_75t_R _20557_ (.A1(net411),
    .A2(_14456_),
    .B(_15209_),
    .C(net320),
    .Y(_15210_));
 INVx1_ASAP7_75t_R _20558_ (.A(_00522_),
    .Y(_15211_));
 NAND2x1_ASAP7_75t_R _20559_ (.A(net2379),
    .B(_00520_),
    .Y(_15212_));
 OA211x2_ASAP7_75t_R _20560_ (.A1(net411),
    .A2(_15211_),
    .B(_15212_),
    .C(net385),
    .Y(_15213_));
 OR3x1_ASAP7_75t_R _20561_ (.A(net318),
    .B(_15210_),
    .C(_15213_),
    .Y(_15214_));
 INVx1_ASAP7_75t_R _20562_ (.A(_00523_),
    .Y(_15215_));
 NAND2x1_ASAP7_75t_R _20563_ (.A(net2379),
    .B(_00521_),
    .Y(_15216_));
 OA211x2_ASAP7_75t_R _20564_ (.A1(net411),
    .A2(_15215_),
    .B(_15216_),
    .C(net385),
    .Y(_15217_));
 NAND2x1_ASAP7_75t_R _20565_ (.A(net2379),
    .B(_00525_),
    .Y(_15218_));
 OA211x2_ASAP7_75t_R _20566_ (.A1(net411),
    .A2(_14453_),
    .B(_15218_),
    .C(net320),
    .Y(_15219_));
 OR3x1_ASAP7_75t_R _20567_ (.A(net425),
    .B(_15217_),
    .C(_15219_),
    .Y(_15220_));
 AND3x1_ASAP7_75t_R _20568_ (.A(net379),
    .B(_15214_),
    .C(_15220_),
    .Y(_15221_));
 OR3x2_ASAP7_75t_R _20569_ (.A(net377),
    .B(_15208_),
    .C(_15221_),
    .Y(_15222_));
 AND3x2_ASAP7_75t_R _20570_ (.A(_13810_),
    .B(_15196_),
    .C(_15222_),
    .Y(_15223_));
 INVx1_ASAP7_75t_R _20571_ (.A(_01634_),
    .Y(_15224_));
 AO32x2_ASAP7_75t_R _20572_ (.A1(\cs_registers_i.pc_id_i[7] ),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_15224_),
    .B2(_13450_),
    .Y(_15225_));
 OR2x2_ASAP7_75t_R _20573_ (.A(_15223_),
    .B(_15225_),
    .Y(_15226_));
 BUFx2_ASAP7_75t_R input125 (.A(net2866),
    .Y(net125));
 INVx2_ASAP7_75t_R _20575_ (.A(_15226_),
    .Y(_18361_));
 OA21x2_ASAP7_75t_R _20576_ (.A1(_00673_),
    .A2(_02266_),
    .B(_02265_),
    .Y(_15227_));
 OR3x1_ASAP7_75t_R _20577_ (.A(_00671_),
    .B(_02266_),
    .C(_16727_),
    .Y(_15228_));
 NAND2x1_ASAP7_75t_R _20578_ (.A(_15227_),
    .B(_15228_),
    .Y(_16730_));
 INVx1_ASAP7_75t_R _20579_ (.A(_01633_),
    .Y(_15229_));
 AND2x2_ASAP7_75t_R _20580_ (.A(_15229_),
    .B(_13450_),
    .Y(_15230_));
 AOI21x1_ASAP7_75t_R _20581_ (.A1(_00186_),
    .A2(_13993_),
    .B(_14988_),
    .Y(_15231_));
 NAND2x1_ASAP7_75t_R _20582_ (.A(net397),
    .B(_00550_),
    .Y(_15232_));
 OA211x2_ASAP7_75t_R _20583_ (.A1(net397),
    .A2(_14527_),
    .B(_15232_),
    .C(net386),
    .Y(_15233_));
 NAND2x1_ASAP7_75t_R _20584_ (.A(net397),
    .B(_00554_),
    .Y(_15234_));
 OA211x2_ASAP7_75t_R _20585_ (.A1(net397),
    .A2(_14524_),
    .B(_15234_),
    .C(net320),
    .Y(_15235_));
 OR3x1_ASAP7_75t_R _20586_ (.A(net318),
    .B(_15233_),
    .C(_15235_),
    .Y(_15236_));
 NAND2x1_ASAP7_75t_R _20587_ (.A(net397),
    .B(_00551_),
    .Y(_15237_));
 OA211x2_ASAP7_75t_R _20588_ (.A1(net397),
    .A2(_14534_),
    .B(_15237_),
    .C(net386),
    .Y(_15238_));
 NAND2x1_ASAP7_75t_R _20589_ (.A(net397),
    .B(_00555_),
    .Y(_15239_));
 OA211x2_ASAP7_75t_R _20590_ (.A1(net397),
    .A2(_14531_),
    .B(_15239_),
    .C(net320),
    .Y(_15240_));
 OR3x1_ASAP7_75t_R _20591_ (.A(net424),
    .B(_15238_),
    .C(_15240_),
    .Y(_15241_));
 INVx1_ASAP7_75t_R _20592_ (.A(_00541_),
    .Y(_15242_));
 NAND2x1_ASAP7_75t_R _20593_ (.A(net397),
    .B(_00539_),
    .Y(_15243_));
 OA211x2_ASAP7_75t_R _20594_ (.A1(net397),
    .A2(_15242_),
    .B(_15243_),
    .C(net318),
    .Y(_15244_));
 INVx1_ASAP7_75t_R _20595_ (.A(_00540_),
    .Y(_15245_));
 NAND2x1_ASAP7_75t_R _20596_ (.A(net411),
    .B(_00538_),
    .Y(_15246_));
 OA211x2_ASAP7_75t_R _20597_ (.A1(net411),
    .A2(_15245_),
    .B(_15246_),
    .C(net424),
    .Y(_15247_));
 OR3x1_ASAP7_75t_R _20598_ (.A(_14015_),
    .B(_15244_),
    .C(_15247_),
    .Y(_15248_));
 NAND2x1_ASAP7_75t_R _20599_ (.A(net397),
    .B(_01701_),
    .Y(_15249_));
 OA211x2_ASAP7_75t_R _20600_ (.A1(net397),
    .A2(_14505_),
    .B(_15249_),
    .C(net318),
    .Y(_15250_));
 AND3x1_ASAP7_75t_R _20601_ (.A(net424),
    .B(net316),
    .C(_14504_),
    .Y(_15251_));
 OA31x2_ASAP7_75t_R _20602_ (.A1(net315),
    .A2(_15250_),
    .A3(_15251_),
    .B1(net378),
    .Y(_15252_));
 AO32x1_ASAP7_75t_R _20603_ (.A1(_13626_),
    .A2(_15236_),
    .A3(_15241_),
    .B1(_15248_),
    .B2(_15252_),
    .Y(_15253_));
 NAND2x1_ASAP7_75t_R _20604_ (.A(net397),
    .B(_00547_),
    .Y(_15254_));
 OA211x2_ASAP7_75t_R _20605_ (.A1(net397),
    .A2(_14482_),
    .B(_15254_),
    .C(net318),
    .Y(_15255_));
 NAND2x1_ASAP7_75t_R _20606_ (.A(net398),
    .B(_00546_),
    .Y(_15256_));
 OA211x2_ASAP7_75t_R _20607_ (.A1(net398),
    .A2(_14485_),
    .B(_15256_),
    .C(net424),
    .Y(_15257_));
 OR3x1_ASAP7_75t_R _20608_ (.A(net386),
    .B(_15255_),
    .C(_15257_),
    .Y(_15258_));
 INVx1_ASAP7_75t_R _20609_ (.A(_00545_),
    .Y(_15259_));
 NAND2x1_ASAP7_75t_R _20610_ (.A(net397),
    .B(_00543_),
    .Y(_15260_));
 OA211x2_ASAP7_75t_R _20611_ (.A1(net397),
    .A2(_15259_),
    .B(_15260_),
    .C(net318),
    .Y(_15261_));
 NAND2x1_ASAP7_75t_R _20612_ (.A(net398),
    .B(_00542_),
    .Y(_15262_));
 OA211x2_ASAP7_75t_R _20613_ (.A1(net398),
    .A2(_14490_),
    .B(_15262_),
    .C(net424),
    .Y(_15263_));
 OR3x1_ASAP7_75t_R _20614_ (.A(net320),
    .B(_15261_),
    .C(_15263_),
    .Y(_15264_));
 AND2x2_ASAP7_75t_R _20615_ (.A(_15258_),
    .B(_15264_),
    .Y(_15265_));
 AND2x2_ASAP7_75t_R _20616_ (.A(_15248_),
    .B(_15252_),
    .Y(_15266_));
 NAND2x1_ASAP7_75t_R _20617_ (.A(net397),
    .B(_00563_),
    .Y(_15267_));
 OA211x2_ASAP7_75t_R _20618_ (.A1(net397),
    .A2(_14517_),
    .B(_15267_),
    .C(net318),
    .Y(_15268_));
 BUFx2_ASAP7_75t_R input124 (.A(net3073),
    .Y(net124));
 NAND2x1_ASAP7_75t_R _20620_ (.A(net397),
    .B(_00562_),
    .Y(_15270_));
 OA211x2_ASAP7_75t_R _20621_ (.A1(net397),
    .A2(_14510_),
    .B(_15270_),
    .C(net424),
    .Y(_15271_));
 OR3x1_ASAP7_75t_R _20622_ (.A(net386),
    .B(_15268_),
    .C(_15271_),
    .Y(_15272_));
 NAND2x1_ASAP7_75t_R _20623_ (.A(net397),
    .B(_00559_),
    .Y(_15273_));
 OA211x2_ASAP7_75t_R _20624_ (.A1(net397),
    .A2(_14520_),
    .B(_15273_),
    .C(net318),
    .Y(_15274_));
 NAND2x1_ASAP7_75t_R _20625_ (.A(net397),
    .B(_00558_),
    .Y(_15275_));
 OA211x2_ASAP7_75t_R _20626_ (.A1(net397),
    .A2(_14513_),
    .B(_15275_),
    .C(net424),
    .Y(_15276_));
 OR3x1_ASAP7_75t_R _20627_ (.A(net320),
    .B(_15274_),
    .C(_15276_),
    .Y(_15277_));
 AND3x1_ASAP7_75t_R _20628_ (.A(_14780_),
    .B(_15272_),
    .C(_15277_),
    .Y(_15278_));
 AO221x2_ASAP7_75t_R _20629_ (.A1(net379),
    .A2(_15253_),
    .B1(_15265_),
    .B2(_15266_),
    .C(_15278_),
    .Y(_15279_));
 OA22x2_ASAP7_75t_R _20630_ (.A1(_15230_),
    .A2(_15231_),
    .B1(_15279_),
    .B2(_15112_),
    .Y(_15280_));
 BUFx2_ASAP7_75t_R input123 (.A(net2882),
    .Y(net123));
 INVx3_ASAP7_75t_R _20632_ (.A(_15280_),
    .Y(_18366_));
 XNOR2x1_ASAP7_75t_R _20633_ (.B(_14599_),
    .Y(_15281_),
    .A(_13620_));
 INVx3_ASAP7_75t_R _20634_ (.A(_00680_),
    .Y(_15282_));
 INVx1_ASAP7_75t_R _20635_ (.A(_01443_),
    .Y(_15283_));
 NAND2x1_ASAP7_75t_R _20636_ (.A(net416),
    .B(_00581_),
    .Y(_15284_));
 OA211x2_ASAP7_75t_R _20637_ (.A1(net416),
    .A2(_14582_),
    .B(_15284_),
    .C(net319),
    .Y(_15285_));
 NAND2x1_ASAP7_75t_R _20638_ (.A(net416),
    .B(_00580_),
    .Y(_15286_));
 OA211x2_ASAP7_75t_R _20639_ (.A1(net416),
    .A2(_14576_),
    .B(_15286_),
    .C(net425),
    .Y(_15287_));
 OR3x1_ASAP7_75t_R _20640_ (.A(net315),
    .B(_15285_),
    .C(_15287_),
    .Y(_15288_));
 NAND2x1_ASAP7_75t_R _20641_ (.A(net416),
    .B(_00584_),
    .Y(_15289_));
 OA211x2_ASAP7_75t_R _20642_ (.A1(net416),
    .A2(_14579_),
    .B(_15289_),
    .C(net426),
    .Y(_15290_));
 NAND2x1_ASAP7_75t_R _20643_ (.A(net416),
    .B(_00585_),
    .Y(_15291_));
 OA211x2_ASAP7_75t_R _20644_ (.A1(net416),
    .A2(_14573_),
    .B(_15291_),
    .C(net319),
    .Y(_15292_));
 OR3x1_ASAP7_75t_R _20645_ (.A(_14015_),
    .B(_15290_),
    .C(_15292_),
    .Y(_15293_));
 AND2x2_ASAP7_75t_R _20646_ (.A(net416),
    .B(_01700_),
    .Y(_15294_));
 AOI21x1_ASAP7_75t_R _20647_ (.A1(_13675_),
    .A2(_00567_),
    .B(_15294_),
    .Y(_15295_));
 AO221x1_ASAP7_75t_R _20648_ (.A1(_14568_),
    .A2(_13687_),
    .B1(_15295_),
    .B2(net319),
    .C(net315),
    .Y(_15296_));
 INVx1_ASAP7_75t_R _20649_ (.A(_00570_),
    .Y(_15297_));
 NAND2x1_ASAP7_75t_R _20650_ (.A(net414),
    .B(_00568_),
    .Y(_15298_));
 OA211x2_ASAP7_75t_R _20651_ (.A1(net414),
    .A2(_15297_),
    .B(_15298_),
    .C(net425),
    .Y(_15299_));
 INVx1_ASAP7_75t_R _20652_ (.A(_00571_),
    .Y(_15300_));
 NAND2x1_ASAP7_75t_R _20653_ (.A(net414),
    .B(_00569_),
    .Y(_15301_));
 OA211x2_ASAP7_75t_R _20654_ (.A1(net414),
    .A2(_15300_),
    .B(_15301_),
    .C(net319),
    .Y(_15302_));
 OA31x2_ASAP7_75t_R _20655_ (.A1(_14015_),
    .A2(_15299_),
    .A3(_15302_),
    .B1(net378),
    .Y(_15303_));
 AO32x1_ASAP7_75t_R _20656_ (.A1(_13626_),
    .A2(_15288_),
    .A3(_15293_),
    .B1(_15296_),
    .B2(_15303_),
    .Y(_15304_));
 NAND2x1_ASAP7_75t_R _20657_ (.A(net418),
    .B(_00577_),
    .Y(_15305_));
 OA211x2_ASAP7_75t_R _20658_ (.A1(net418),
    .A2(_14555_),
    .B(_15305_),
    .C(_13649_),
    .Y(_15306_));
 NAND2x1_ASAP7_75t_R _20659_ (.A(net418),
    .B(_00576_),
    .Y(_15307_));
 OA211x2_ASAP7_75t_R _20660_ (.A1(net418),
    .A2(_14549_),
    .B(_15307_),
    .C(net419),
    .Y(_15308_));
 OR3x2_ASAP7_75t_R _20661_ (.A(net388),
    .B(_15306_),
    .C(_15308_),
    .Y(_15309_));
 INVx1_ASAP7_75t_R _20662_ (.A(_00575_),
    .Y(_15310_));
 NAND2x1_ASAP7_75t_R _20663_ (.A(net418),
    .B(_00573_),
    .Y(_15311_));
 OA211x2_ASAP7_75t_R _20664_ (.A1(net418),
    .A2(_15310_),
    .B(_15311_),
    .C(_13649_),
    .Y(_15312_));
 NAND2x1_ASAP7_75t_R _20665_ (.A(net393),
    .B(_00572_),
    .Y(_15313_));
 OA211x2_ASAP7_75t_R _20666_ (.A1(net418),
    .A2(_14552_),
    .B(_15313_),
    .C(net427),
    .Y(_15314_));
 OR3x1_ASAP7_75t_R _20667_ (.A(_13630_),
    .B(_15312_),
    .C(_15314_),
    .Y(_15315_));
 AND4x1_ASAP7_75t_R _20668_ (.A(_15296_),
    .B(_15303_),
    .C(_15309_),
    .D(_15315_),
    .Y(_15316_));
 INVx1_ASAP7_75t_R _20669_ (.A(_00591_),
    .Y(_15317_));
 NAND2x1_ASAP7_75t_R _20670_ (.A(net398),
    .B(_00589_),
    .Y(_15318_));
 OA211x2_ASAP7_75t_R _20671_ (.A1(net398),
    .A2(_15317_),
    .B(_15318_),
    .C(net319),
    .Y(_15319_));
 NAND2x1_ASAP7_75t_R _20672_ (.A(net398),
    .B(_00588_),
    .Y(_15320_));
 OA211x2_ASAP7_75t_R _20673_ (.A1(net398),
    .A2(_14588_),
    .B(_15320_),
    .C(net425),
    .Y(_15321_));
 OR3x1_ASAP7_75t_R _20674_ (.A(net321),
    .B(_15319_),
    .C(_15321_),
    .Y(_15322_));
 INVx1_ASAP7_75t_R _20675_ (.A(_00595_),
    .Y(_15323_));
 NAND2x1_ASAP7_75t_R _20676_ (.A(net414),
    .B(_00593_),
    .Y(_15324_));
 OA211x2_ASAP7_75t_R _20677_ (.A1(net414),
    .A2(_15323_),
    .B(_15324_),
    .C(net319),
    .Y(_15325_));
 INVx1_ASAP7_75t_R _20678_ (.A(_00594_),
    .Y(_15326_));
 NAND2x1_ASAP7_75t_R _20679_ (.A(net398),
    .B(_00592_),
    .Y(_15327_));
 OA211x2_ASAP7_75t_R _20680_ (.A1(net410),
    .A2(_15326_),
    .B(_15327_),
    .C(net425),
    .Y(_15328_));
 OR3x1_ASAP7_75t_R _20681_ (.A(net386),
    .B(_15325_),
    .C(_15328_),
    .Y(_15329_));
 AND5x1_ASAP7_75t_R _20682_ (.A(_13626_),
    .B(_15288_),
    .C(_15293_),
    .D(_15322_),
    .E(_15329_),
    .Y(_15330_));
 AO211x2_ASAP7_75t_R _20683_ (.A1(net380),
    .A2(_15304_),
    .B(_15316_),
    .C(_15330_),
    .Y(_15331_));
 OA222x2_ASAP7_75t_R _20684_ (.A1(_00285_),
    .A2(_15282_),
    .B1(_15283_),
    .B2(_13815_),
    .C1(_15331_),
    .C2(_00284_),
    .Y(_15332_));
 AND2x2_ASAP7_75t_R _20685_ (.A(_13772_),
    .B(_14597_),
    .Y(_15333_));
 AOI211x1_ASAP7_75t_R _20686_ (.A1(_13986_),
    .A2(_15332_),
    .B(_15333_),
    .C(net309),
    .Y(_15334_));
 AO21x1_ASAP7_75t_R _20687_ (.A1(net309),
    .A2(_15281_),
    .B(_15334_),
    .Y(_17770_));
 INVx1_ASAP7_75t_R _20688_ (.A(_17770_),
    .Y(_16731_));
 INVx2_ASAP7_75t_R _20689_ (.A(_00189_),
    .Y(\cs_registers_i.pc_id_i[9] ));
 NOR2x1_ASAP7_75t_R _20690_ (.A(_01632_),
    .B(_13807_),
    .Y(_15335_));
 OA21x2_ASAP7_75t_R _20691_ (.A1(\cs_registers_i.pc_id_i[9] ),
    .A2(_13808_),
    .B(_13794_),
    .Y(_15336_));
 OA22x2_ASAP7_75t_R _20692_ (.A1(_15112_),
    .A2(_15331_),
    .B1(_15335_),
    .B2(_15336_),
    .Y(_15337_));
 BUFx2_ASAP7_75t_R input122 (.A(net3118),
    .Y(net122));
 INVx3_ASAP7_75t_R _20694_ (.A(_15337_),
    .Y(_18371_));
 BUFx2_ASAP7_75t_R input121 (.A(net2957),
    .Y(net121));
 AND3x1_ASAP7_75t_R _20696_ (.A(_15282_),
    .B(_13817_),
    .C(_13778_),
    .Y(_15339_));
 AO21x1_ASAP7_75t_R _20697_ (.A1(net309),
    .A2(_15337_),
    .B(_15339_),
    .Y(_17771_));
 INVx1_ASAP7_75t_R _20698_ (.A(_17771_),
    .Y(_16732_));
 OA21x2_ASAP7_75t_R _20699_ (.A1(_00678_),
    .A2(_02268_),
    .B(_02267_),
    .Y(_15340_));
 AO21x1_ASAP7_75t_R _20700_ (.A1(_00673_),
    .A2(_00671_),
    .B(_02266_),
    .Y(_15341_));
 OR2x2_ASAP7_75t_R _20701_ (.A(_00675_),
    .B(_02268_),
    .Y(_15342_));
 AO21x1_ASAP7_75t_R _20702_ (.A1(_02265_),
    .A2(_15341_),
    .B(_15342_),
    .Y(_15343_));
 AO21x1_ASAP7_75t_R _20703_ (.A1(_16727_),
    .A2(_15227_),
    .B(_15343_),
    .Y(_15344_));
 AND2x2_ASAP7_75t_R _20704_ (.A(_15340_),
    .B(_15344_),
    .Y(_16733_));
 INVx1_ASAP7_75t_R _20705_ (.A(_00612_),
    .Y(_15345_));
 NAND2x1_ASAP7_75t_R _20706_ (.A(net405),
    .B(_00610_),
    .Y(_15346_));
 OA211x2_ASAP7_75t_R _20707_ (.A1(net405),
    .A2(_15345_),
    .B(_15346_),
    .C(net384),
    .Y(_15347_));
 NAND2x1_ASAP7_75t_R _20708_ (.A(net405),
    .B(_00614_),
    .Y(_15348_));
 OA211x2_ASAP7_75t_R _20709_ (.A1(net405),
    .A2(_14629_),
    .B(_15348_),
    .C(net320),
    .Y(_15349_));
 OR3x1_ASAP7_75t_R _20710_ (.A(net318),
    .B(_15347_),
    .C(_15349_),
    .Y(_15350_));
 INVx1_ASAP7_75t_R _20711_ (.A(_00613_),
    .Y(_15351_));
 NAND2x1_ASAP7_75t_R _20712_ (.A(net405),
    .B(_00611_),
    .Y(_15352_));
 OA211x2_ASAP7_75t_R _20713_ (.A1(net405),
    .A2(_15351_),
    .B(_15352_),
    .C(net384),
    .Y(_15353_));
 NAND2x1_ASAP7_75t_R _20714_ (.A(net405),
    .B(_00615_),
    .Y(_15354_));
 OA211x2_ASAP7_75t_R _20715_ (.A1(net405),
    .A2(_14626_),
    .B(_15354_),
    .C(net320),
    .Y(_15355_));
 OR3x1_ASAP7_75t_R _20716_ (.A(net420),
    .B(_15353_),
    .C(_15355_),
    .Y(_15356_));
 NAND2x1_ASAP7_75t_R _20717_ (.A(net405),
    .B(_00599_),
    .Y(_15357_));
 OA211x2_ASAP7_75t_R _20718_ (.A1(net405),
    .A2(_14618_),
    .B(_15357_),
    .C(net318),
    .Y(_15358_));
 NAND2x1_ASAP7_75t_R _20719_ (.A(net405),
    .B(_00598_),
    .Y(_15359_));
 OA211x2_ASAP7_75t_R _20720_ (.A1(net405),
    .A2(_14621_),
    .B(_15359_),
    .C(net420),
    .Y(_15360_));
 OR3x1_ASAP7_75t_R _20721_ (.A(net312),
    .B(_15358_),
    .C(_15360_),
    .Y(_15361_));
 INVx1_ASAP7_75t_R _20722_ (.A(_00597_),
    .Y(_15362_));
 NAND2x1_ASAP7_75t_R _20723_ (.A(net405),
    .B(_01699_),
    .Y(_15363_));
 OA211x2_ASAP7_75t_R _20724_ (.A1(net405),
    .A2(_15362_),
    .B(_15363_),
    .C(net318),
    .Y(_15364_));
 NOR2x1_ASAP7_75t_R _20725_ (.A(net405),
    .B(_00596_),
    .Y(_15365_));
 AO21x1_ASAP7_75t_R _20726_ (.A1(net420),
    .A2(_15365_),
    .B(_14005_),
    .Y(_15366_));
 OA21x2_ASAP7_75t_R _20727_ (.A1(_15364_),
    .A2(_15366_),
    .B(net377),
    .Y(_15367_));
 AO32x1_ASAP7_75t_R _20728_ (.A1(_13626_),
    .A2(_15350_),
    .A3(_15356_),
    .B1(_15361_),
    .B2(_15367_),
    .Y(_15368_));
 NAND2x1_ASAP7_75t_R _20729_ (.A(net402),
    .B(_00607_),
    .Y(_15369_));
 OA211x2_ASAP7_75t_R _20730_ (.A1(net2376),
    .A2(_14608_),
    .B(_15369_),
    .C(net317),
    .Y(_15370_));
 NAND2x1_ASAP7_75t_R _20731_ (.A(net402),
    .B(_00606_),
    .Y(_15371_));
 OA211x2_ASAP7_75t_R _20732_ (.A1(net2376),
    .A2(_14600_),
    .B(_15371_),
    .C(net420),
    .Y(_15372_));
 OR3x1_ASAP7_75t_R _20733_ (.A(net384),
    .B(_15370_),
    .C(_15372_),
    .Y(_15373_));
 INVx1_ASAP7_75t_R _20734_ (.A(_00605_),
    .Y(_15374_));
 NAND2x1_ASAP7_75t_R _20735_ (.A(net402),
    .B(_00603_),
    .Y(_15375_));
 OA211x2_ASAP7_75t_R _20736_ (.A1(net2376),
    .A2(_15374_),
    .B(_15375_),
    .C(net317),
    .Y(_15376_));
 INVx1_ASAP7_75t_R _20737_ (.A(_00604_),
    .Y(_15377_));
 NAND2x1_ASAP7_75t_R _20738_ (.A(net402),
    .B(_00602_),
    .Y(_15378_));
 OA211x2_ASAP7_75t_R _20739_ (.A1(net2376),
    .A2(_15377_),
    .B(_15378_),
    .C(net420),
    .Y(_15379_));
 OR3x1_ASAP7_75t_R _20740_ (.A(net320),
    .B(_15376_),
    .C(_15379_),
    .Y(_15380_));
 AND2x2_ASAP7_75t_R _20741_ (.A(_15373_),
    .B(_15380_),
    .Y(_15381_));
 AND2x2_ASAP7_75t_R _20742_ (.A(_15361_),
    .B(_15367_),
    .Y(_15382_));
 INVx1_ASAP7_75t_R _20743_ (.A(_00618_),
    .Y(_15383_));
 NOR2x1_ASAP7_75t_R _20744_ (.A(net384),
    .B(_00622_),
    .Y(_15384_));
 AO21x1_ASAP7_75t_R _20745_ (.A1(net384),
    .A2(_15383_),
    .B(_15384_),
    .Y(_15385_));
 NAND2x1_ASAP7_75t_R _20746_ (.A(net384),
    .B(_00620_),
    .Y(_15386_));
 OA211x2_ASAP7_75t_R _20747_ (.A1(net384),
    .A2(_14638_),
    .B(_15386_),
    .C(net316),
    .Y(_15387_));
 AO21x1_ASAP7_75t_R _20748_ (.A1(net405),
    .A2(_15385_),
    .B(_15387_),
    .Y(_15388_));
 INVx1_ASAP7_75t_R _20749_ (.A(_00621_),
    .Y(_15389_));
 NAND2x1_ASAP7_75t_R _20750_ (.A(net402),
    .B(_00619_),
    .Y(_15390_));
 OA211x2_ASAP7_75t_R _20751_ (.A1(net2376),
    .A2(_15389_),
    .B(_15390_),
    .C(net384),
    .Y(_15391_));
 NAND2x1_ASAP7_75t_R _20752_ (.A(net405),
    .B(_00623_),
    .Y(_15392_));
 OA211x2_ASAP7_75t_R _20753_ (.A1(net405),
    .A2(_14641_),
    .B(_15392_),
    .C(net320),
    .Y(_15393_));
 OR3x1_ASAP7_75t_R _20754_ (.A(net420),
    .B(_15391_),
    .C(_15393_),
    .Y(_15394_));
 OA211x2_ASAP7_75t_R _20755_ (.A1(net318),
    .A2(_15388_),
    .B(_15394_),
    .C(_14780_),
    .Y(_15395_));
 AO221x2_ASAP7_75t_R _20756_ (.A1(net380),
    .A2(_15368_),
    .B1(_15381_),
    .B2(_15382_),
    .C(_15395_),
    .Y(_15396_));
 BUFx2_ASAP7_75t_R input120 (.A(net2858),
    .Y(net120));
 INVx2_ASAP7_75t_R _20758_ (.A(_00193_),
    .Y(_15398_));
 INVx1_ASAP7_75t_R _20759_ (.A(_01631_),
    .Y(_15399_));
 AO32x2_ASAP7_75t_R _20760_ (.A1(_15398_),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_15399_),
    .B2(_13450_),
    .Y(_15400_));
 AO21x2_ASAP7_75t_R _20761_ (.A1(_13810_),
    .A2(net2310),
    .B(_15400_),
    .Y(_15401_));
 BUFx2_ASAP7_75t_R input119 (.A(net2810),
    .Y(net119));
 INVx2_ASAP7_75t_R _20763_ (.A(_15401_),
    .Y(_18376_));
 XNOR2x1_ASAP7_75t_R _20764_ (.B(_18380_),
    .Y(_15402_),
    .A(_13620_));
 BUFx2_ASAP7_75t_R input118 (.A(net2842),
    .Y(net118));
 INVx1_ASAP7_75t_R _20766_ (.A(_00684_),
    .Y(_15404_));
 INVx1_ASAP7_75t_R _20767_ (.A(_01441_),
    .Y(_15405_));
 OA222x2_ASAP7_75t_R _20768_ (.A1(_00285_),
    .A2(_15404_),
    .B1(_15405_),
    .B2(_13815_),
    .C1(_14783_),
    .C2(_00284_),
    .Y(_15406_));
 NAND2x1_ASAP7_75t_R _20769_ (.A(_13986_),
    .B(_15406_),
    .Y(_15407_));
 OA211x2_ASAP7_75t_R _20770_ (.A1(_13986_),
    .A2(_14703_),
    .B(_15407_),
    .C(_13817_),
    .Y(_15408_));
 AO21x1_ASAP7_75t_R _20771_ (.A1(net309),
    .A2(_15402_),
    .B(_15408_),
    .Y(_17775_));
 INVx1_ASAP7_75t_R _20772_ (.A(_17775_),
    .Y(_16736_));
 OA21x2_ASAP7_75t_R _20773_ (.A1(_00684_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_15409_));
 AOI21x1_ASAP7_75t_R _20774_ (.A1(net309),
    .A2(_18379_),
    .B(_15409_),
    .Y(_17774_));
 INVx1_ASAP7_75t_R _20775_ (.A(_17774_),
    .Y(_16734_));
 OA21x2_ASAP7_75t_R _20776_ (.A1(_00681_),
    .A2(_16733_),
    .B(_00683_),
    .Y(_15410_));
 OA21x2_ASAP7_75t_R _20777_ (.A1(_02270_),
    .A2(_15410_),
    .B(_02269_),
    .Y(_16735_));
 BUFx2_ASAP7_75t_R input117 (.A(net2906),
    .Y(net117));
 BUFx2_ASAP7_75t_R input116 (.A(net2777),
    .Y(net116));
 BUFx2_ASAP7_75t_R input115 (.A(net2850),
    .Y(net115));
 BUFx2_ASAP7_75t_R input114 (.A(net2941),
    .Y(net114));
 BUFx2_ASAP7_75t_R input113 (.A(net2914),
    .Y(net113));
 BUFx2_ASAP7_75t_R input112 (.A(net3110),
    .Y(net112));
 BUFx2_ASAP7_75t_R input111 (.A(net2927),
    .Y(net111));
 BUFx2_ASAP7_75t_R input110 (.A(net3081),
    .Y(net110));
 BUFx2_ASAP7_75t_R input109 (.A(net2874),
    .Y(net109));
 BUFx2_ASAP7_75t_R input108 (.A(net3094),
    .Y(net108));
 AND2x2_ASAP7_75t_R _20788_ (.A(net2371),
    .B(_01697_),
    .Y(_15421_));
 AO21x1_ASAP7_75t_R _20789_ (.A1(net2260),
    .A2(_00326_),
    .B(_15421_),
    .Y(_15422_));
 BUFx2_ASAP7_75t_R input107 (.A(net3018),
    .Y(net107));
 BUFx2_ASAP7_75t_R input106 (.A(net3006),
    .Y(net106));
 BUFx2_ASAP7_75t_R input105 (.A(net2890),
    .Y(net105));
 OAI22x1_ASAP7_75t_R _20793_ (.A1(_00325_),
    .A2(_14184_),
    .B1(_15422_),
    .B2(net371),
    .Y(_15426_));
 BUFx3_ASAP7_75t_R input104 (.A(net2898),
    .Y(net104));
 BUFx2_ASAP7_75t_R input103 (.A(net2990),
    .Y(net103));
 BUFx2_ASAP7_75t_R input102 (.A(net2764),
    .Y(net102));
 BUFx2_ASAP7_75t_R input101 (.A(net2826),
    .Y(net101));
 NAND2x1_ASAP7_75t_R _20798_ (.A(net356),
    .B(_00332_),
    .Y(_15431_));
 BUFx2_ASAP7_75t_R input100 (.A(net2818),
    .Y(net100));
 BUFx2_ASAP7_75t_R input99 (.A(net2785),
    .Y(net99));
 OA211x2_ASAP7_75t_R _20801_ (.A1(net356),
    .A2(_14059_),
    .B(_15431_),
    .C(net324),
    .Y(_15434_));
 BUFx2_ASAP7_75t_R input98 (.A(net2834),
    .Y(net98));
 NAND2x1_ASAP7_75t_R _20803_ (.A(net356),
    .B(_00331_),
    .Y(_15436_));
 BUFx2_ASAP7_75t_R input97 (.A(net2949),
    .Y(net97));
 OA211x2_ASAP7_75t_R _20805_ (.A1(net356),
    .A2(_14052_),
    .B(_15436_),
    .C(net372),
    .Y(_15438_));
 OR3x1_ASAP7_75t_R _20806_ (.A(net330),
    .B(_15434_),
    .C(_15438_),
    .Y(_15439_));
 OA21x2_ASAP7_75t_R _20807_ (.A1(_13373_),
    .A2(_15426_),
    .B(_15439_),
    .Y(_15440_));
 BUFx2_ASAP7_75t_R input96 (.A(net2998),
    .Y(net96));
 BUFx2_ASAP7_75t_R input95 (.A(net3294),
    .Y(net95));
 BUFx2_ASAP7_75t_R input94 (.A(net2965),
    .Y(net94));
 NAND2x1_ASAP7_75t_R _20811_ (.A(net357),
    .B(_00328_),
    .Y(_15444_));
 OA211x2_ASAP7_75t_R _20812_ (.A1(net357),
    .A2(_14022_),
    .B(_15444_),
    .C(net324),
    .Y(_15445_));
 BUFx2_ASAP7_75t_R input93 (.A(net3713),
    .Y(net93));
 NAND2x1_ASAP7_75t_R _20814_ (.A(net357),
    .B(_00327_),
    .Y(_15447_));
 BUFx2_ASAP7_75t_R input92 (.A(net3722),
    .Y(net92));
 OA211x2_ASAP7_75t_R _20816_ (.A1(net357),
    .A2(_14019_),
    .B(_15447_),
    .C(net371),
    .Y(_15449_));
 OR3x1_ASAP7_75t_R _20817_ (.A(_13373_),
    .B(_15445_),
    .C(_15449_),
    .Y(_15450_));
 NAND2x1_ASAP7_75t_R _20818_ (.A(net356),
    .B(_00336_),
    .Y(_15451_));
 BUFx2_ASAP7_75t_R input91 (.A(net3652),
    .Y(net91));
 OA211x2_ASAP7_75t_R _20820_ (.A1(net356),
    .A2(_14069_),
    .B(_15451_),
    .C(net324),
    .Y(_15453_));
 NAND2x1_ASAP7_75t_R _20821_ (.A(net356),
    .B(_00335_),
    .Y(_15454_));
 OA211x2_ASAP7_75t_R _20822_ (.A1(net356),
    .A2(_14066_),
    .B(_15454_),
    .C(net372),
    .Y(_15455_));
 OR3x1_ASAP7_75t_R _20823_ (.A(net330),
    .B(_15453_),
    .C(_15455_),
    .Y(_15456_));
 AND3x1_ASAP7_75t_R _20824_ (.A(_13350_),
    .B(_15450_),
    .C(_15456_),
    .Y(_15457_));
 AO21x1_ASAP7_75t_R _20825_ (.A1(net334),
    .A2(_15440_),
    .B(_15457_),
    .Y(_15458_));
 BUFx2_ASAP7_75t_R input90 (.A(net3743),
    .Y(net90));
 BUFx2_ASAP7_75t_R input89 (.A(net3635),
    .Y(net89));
 NAND2x1_ASAP7_75t_R _20828_ (.A(net2281),
    .B(_00340_),
    .Y(_15461_));
 OA211x2_ASAP7_75t_R _20829_ (.A1(net2372),
    .A2(_14043_),
    .B(_15461_),
    .C(net324),
    .Y(_15462_));
 NAND2x1_ASAP7_75t_R _20830_ (.A(net2281),
    .B(_00339_),
    .Y(_15463_));
 OA211x2_ASAP7_75t_R _20831_ (.A1(net2372),
    .A2(_14033_),
    .B(_15463_),
    .C(net371),
    .Y(_15464_));
 OR3x1_ASAP7_75t_R _20832_ (.A(_13350_),
    .B(_15462_),
    .C(_15464_),
    .Y(_15465_));
 NAND2x1_ASAP7_75t_R _20833_ (.A(net357),
    .B(_00344_),
    .Y(_15466_));
 OA211x2_ASAP7_75t_R _20834_ (.A1(net357),
    .A2(_14040_),
    .B(_15466_),
    .C(net324),
    .Y(_15467_));
 BUFx2_ASAP7_75t_R input88 (.A(net3382),
    .Y(net88));
 BUFx2_ASAP7_75t_R input87 (.A(net3560),
    .Y(net87));
 NAND2x1_ASAP7_75t_R _20837_ (.A(net357),
    .B(_00343_),
    .Y(_15470_));
 OA211x2_ASAP7_75t_R _20838_ (.A1(net357),
    .A2(_14027_),
    .B(_15470_),
    .C(net371),
    .Y(_15471_));
 OR3x1_ASAP7_75t_R _20839_ (.A(net334),
    .B(_15467_),
    .C(_15471_),
    .Y(_15472_));
 AND3x1_ASAP7_75t_R _20840_ (.A(net330),
    .B(_15465_),
    .C(_15472_),
    .Y(_15473_));
 BUFx2_ASAP7_75t_R input86 (.A(net3574),
    .Y(net86));
 NAND2x1_ASAP7_75t_R _20842_ (.A(net356),
    .B(_00352_),
    .Y(_15475_));
 OA211x2_ASAP7_75t_R _20843_ (.A1(net356),
    .A2(_14078_),
    .B(_15475_),
    .C(net324),
    .Y(_15476_));
 NAND2x1_ASAP7_75t_R _20844_ (.A(net356),
    .B(_00351_),
    .Y(_15477_));
 OA211x2_ASAP7_75t_R _20845_ (.A1(net356),
    .A2(_14090_),
    .B(_15477_),
    .C(net372),
    .Y(_15478_));
 OR3x1_ASAP7_75t_R _20846_ (.A(net334),
    .B(_15476_),
    .C(_15478_),
    .Y(_15479_));
 NAND2x1_ASAP7_75t_R _20847_ (.A(net356),
    .B(_00348_),
    .Y(_15480_));
 OA211x2_ASAP7_75t_R _20848_ (.A1(net356),
    .A2(_14082_),
    .B(_15480_),
    .C(net324),
    .Y(_15481_));
 NAND2x1_ASAP7_75t_R _20849_ (.A(net356),
    .B(_00347_),
    .Y(_15482_));
 OA211x2_ASAP7_75t_R _20850_ (.A1(net356),
    .A2(_14093_),
    .B(_15482_),
    .C(net372),
    .Y(_15483_));
 OR3x1_ASAP7_75t_R _20851_ (.A(_13350_),
    .B(_15481_),
    .C(_15483_),
    .Y(_15484_));
 AND3x1_ASAP7_75t_R _20852_ (.A(_13373_),
    .B(_15479_),
    .C(_15484_),
    .Y(_15485_));
 OR3x1_ASAP7_75t_R _20853_ (.A(net327),
    .B(_15473_),
    .C(_15485_),
    .Y(_15486_));
 OA21x2_ASAP7_75t_R _20854_ (.A1(_13355_),
    .A2(_15458_),
    .B(_15486_),
    .Y(_15487_));
 INVx2_ASAP7_75t_R _20855_ (.A(_15487_),
    .Y(_15488_));
 OR3x4_ASAP7_75t_R _20856_ (.A(_13507_),
    .B(_13510_),
    .C(_13481_),
    .Y(_15489_));
 OA21x2_ASAP7_75t_R _20857_ (.A1(_13520_),
    .A2(_13888_),
    .B(_15489_),
    .Y(_15490_));
 BUFx2_ASAP7_75t_R input85 (.A(net3694),
    .Y(net85));
 OA21x2_ASAP7_75t_R _20859_ (.A1(_00280_),
    .A2(_13506_),
    .B(_13521_),
    .Y(_15492_));
 BUFx2_ASAP7_75t_R input84 (.A(net3535),
    .Y(net84));
 OA21x2_ASAP7_75t_R _20861_ (.A1(_00281_),
    .A2(_15490_),
    .B(_15492_),
    .Y(_15494_));
 AO21x1_ASAP7_75t_R _20862_ (.A1(_13474_),
    .A2(_15488_),
    .B(_15494_),
    .Y(_18386_));
 INVx1_ASAP7_75t_R _20863_ (.A(_18386_),
    .Y(_18384_));
 BUFx2_ASAP7_75t_R input83 (.A(net3606),
    .Y(net83));
 BUFx2_ASAP7_75t_R input82 (.A(net3739),
    .Y(net82));
 BUFx2_ASAP7_75t_R input81 (.A(net3617),
    .Y(net81));
 BUFx2_ASAP7_75t_R input80 (.A(net3749),
    .Y(net80));
 BUFx2_ASAP7_75t_R input79 (.A(net3642),
    .Y(net79));
 BUFx2_ASAP7_75t_R input78 (.A(net3588),
    .Y(net78));
 BUFx2_ASAP7_75t_R input77 (.A(net3597),
    .Y(net77));
 BUFx2_ASAP7_75t_R input76 (.A(net3687),
    .Y(net76));
 BUFx2_ASAP7_75t_R input75 (.A(net3674),
    .Y(net75));
 BUFx2_ASAP7_75t_R input74 (.A(net3679),
    .Y(net74));
 INVx1_ASAP7_75t_R _20874_ (.A(_00698_),
    .Y(_15505_));
 BUFx2_ASAP7_75t_R input73 (.A(net3650),
    .Y(net73));
 NOR2x1_ASAP7_75t_R _20876_ (.A(net339),
    .B(_00700_),
    .Y(_15507_));
 AO21x1_ASAP7_75t_R _20877_ (.A1(net339),
    .A2(_15505_),
    .B(_15507_),
    .Y(_15508_));
 BUFx2_ASAP7_75t_R input72 (.A(net3718),
    .Y(net72));
 INVx1_ASAP7_75t_R _20879_ (.A(_00701_),
    .Y(_15510_));
 BUFx2_ASAP7_75t_R input71 (.A(net3568),
    .Y(net71));
 NAND2x1_ASAP7_75t_R _20881_ (.A(net339),
    .B(_00699_),
    .Y(_15512_));
 BUFx2_ASAP7_75t_R input70 (.A(net3657),
    .Y(net70));
 OA211x2_ASAP7_75t_R _20883_ (.A1(net339),
    .A2(_15510_),
    .B(_15512_),
    .C(net325),
    .Y(_15514_));
 AO21x1_ASAP7_75t_R _20884_ (.A1(net370),
    .A2(_15508_),
    .B(_15514_),
    .Y(_15515_));
 BUFx2_ASAP7_75t_R input69 (.A(net3620),
    .Y(net69));
 BUFx2_ASAP7_75t_R input68 (.A(net3767),
    .Y(net68));
 INVx1_ASAP7_75t_R _20887_ (.A(_00693_),
    .Y(_15518_));
 BUFx2_ASAP7_75t_R input67 (.A(net3584),
    .Y(net67));
 NAND2x1_ASAP7_75t_R _20889_ (.A(net339),
    .B(_00691_),
    .Y(_15520_));
 BUFx2_ASAP7_75t_R input66 (.A(net3731),
    .Y(net66));
 OA211x2_ASAP7_75t_R _20891_ (.A1(net339),
    .A2(_15518_),
    .B(_15520_),
    .C(net325),
    .Y(_15522_));
 INVx1_ASAP7_75t_R _20892_ (.A(_00692_),
    .Y(_15523_));
 NAND2x1_ASAP7_75t_R _20893_ (.A(net339),
    .B(_00690_),
    .Y(_15524_));
 BUFx2_ASAP7_75t_R input65 (.A(net3670),
    .Y(net65));
 OA211x2_ASAP7_75t_R _20895_ (.A1(net339),
    .A2(_15523_),
    .B(_15524_),
    .C(net370),
    .Y(_15526_));
 OR3x1_ASAP7_75t_R _20896_ (.A(_13373_),
    .B(_15522_),
    .C(_15526_),
    .Y(_15527_));
 OA21x2_ASAP7_75t_R _20897_ (.A1(net331),
    .A2(_15515_),
    .B(_15527_),
    .Y(_15528_));
 BUFx2_ASAP7_75t_R input64 (.A(net3700),
    .Y(net64));
 BUFx2_ASAP7_75t_R input63 (.A(net3733),
    .Y(net63));
 BUFx2_ASAP7_75t_R input62 (.A(net3627),
    .Y(net62));
 BUFx2_ASAP7_75t_R input61 (.A(net3946),
    .Y(net61));
 AND2x2_ASAP7_75t_R _20902_ (.A(net346),
    .B(_01696_),
    .Y(_15533_));
 AO21x1_ASAP7_75t_R _20903_ (.A1(_13359_),
    .A2(_00689_),
    .B(_15533_),
    .Y(_15534_));
 OAI22x1_ASAP7_75t_R _20904_ (.A1(_00688_),
    .A2(net311),
    .B1(_15534_),
    .B2(net369),
    .Y(_15535_));
 BUFx2_ASAP7_75t_R input60 (.A(net3182),
    .Y(net60));
 INVx1_ASAP7_75t_R _20906_ (.A(_00697_),
    .Y(_15537_));
 NAND2x1_ASAP7_75t_R _20907_ (.A(net339),
    .B(_00695_),
    .Y(_15538_));
 BUFx4f_ASAP7_75t_R input59 (.A(net3138),
    .Y(net59));
 OA211x2_ASAP7_75t_R _20909_ (.A1(net339),
    .A2(_15537_),
    .B(_15538_),
    .C(net323),
    .Y(_15540_));
 INVx1_ASAP7_75t_R _20910_ (.A(_00696_),
    .Y(_15541_));
 NAND2x1_ASAP7_75t_R _20911_ (.A(net339),
    .B(_00694_),
    .Y(_15542_));
 BUFx2_ASAP7_75t_R input58 (.A(net4033),
    .Y(net58));
 OA211x2_ASAP7_75t_R _20913_ (.A1(net339),
    .A2(_15541_),
    .B(_15542_),
    .C(net369),
    .Y(_15544_));
 OR3x1_ASAP7_75t_R _20914_ (.A(net331),
    .B(_15540_),
    .C(_15544_),
    .Y(_15545_));
 OA211x2_ASAP7_75t_R _20915_ (.A1(_13373_),
    .A2(_15535_),
    .B(_15545_),
    .C(net337),
    .Y(_15546_));
 AO21x1_ASAP7_75t_R _20916_ (.A1(_13350_),
    .A2(_15528_),
    .B(_15546_),
    .Y(_15547_));
 BUFx2_ASAP7_75t_R input57 (.A(net3982),
    .Y(net57));
 BUFx2_ASAP7_75t_R input56 (.A(net3762),
    .Y(net56));
 BUFx2_ASAP7_75t_R input55 (.A(net3768),
    .Y(net55));
 INVx1_ASAP7_75t_R _20920_ (.A(_00705_),
    .Y(_15551_));
 BUFx2_ASAP7_75t_R input54 (.A(net3774),
    .Y(net54));
 NAND2x1_ASAP7_75t_R _20922_ (.A(net348),
    .B(_00703_),
    .Y(_15553_));
 BUFx2_ASAP7_75t_R input53 (.A(net3785),
    .Y(net53));
 OA211x2_ASAP7_75t_R _20924_ (.A1(net348),
    .A2(_15551_),
    .B(_15553_),
    .C(net325),
    .Y(_15555_));
 BUFx2_ASAP7_75t_R input52 (.A(data_rdata_i[3]),
    .Y(net52));
 INVx1_ASAP7_75t_R _20926_ (.A(_00704_),
    .Y(_15557_));
 BUFx2_ASAP7_75t_R input51 (.A(net4038),
    .Y(net51));
 NAND2x1_ASAP7_75t_R _20928_ (.A(net346),
    .B(_00702_),
    .Y(_15559_));
 BUFx2_ASAP7_75t_R input50 (.A(net3988),
    .Y(net50));
 OA211x2_ASAP7_75t_R _20930_ (.A1(net346),
    .A2(_15557_),
    .B(_15559_),
    .C(net369),
    .Y(_15561_));
 OR3x1_ASAP7_75t_R _20931_ (.A(_13350_),
    .B(_15555_),
    .C(_15561_),
    .Y(_15562_));
 BUFx2_ASAP7_75t_R input49 (.A(net3771),
    .Y(net49));
 INVx1_ASAP7_75t_R _20933_ (.A(_00709_),
    .Y(_15564_));
 NAND2x1_ASAP7_75t_R _20934_ (.A(net339),
    .B(_00707_),
    .Y(_15565_));
 OA211x2_ASAP7_75t_R _20935_ (.A1(net339),
    .A2(_15564_),
    .B(_15565_),
    .C(net325),
    .Y(_15566_));
 INVx1_ASAP7_75t_R _20936_ (.A(_00708_),
    .Y(_15567_));
 BUFx2_ASAP7_75t_R input48 (.A(net3956),
    .Y(net48));
 NAND2x1_ASAP7_75t_R _20938_ (.A(net339),
    .B(_00706_),
    .Y(_15569_));
 OA211x2_ASAP7_75t_R _20939_ (.A1(net339),
    .A2(_15567_),
    .B(_15569_),
    .C(net369),
    .Y(_15570_));
 OR3x1_ASAP7_75t_R _20940_ (.A(net337),
    .B(_15566_),
    .C(_15570_),
    .Y(_15571_));
 AND3x1_ASAP7_75t_R _20941_ (.A(net331),
    .B(_15562_),
    .C(_15571_),
    .Y(_15572_));
 INVx1_ASAP7_75t_R _20942_ (.A(_00712_),
    .Y(_15573_));
 NAND2x1_ASAP7_75t_R _20943_ (.A(net346),
    .B(_00710_),
    .Y(_15574_));
 OA211x2_ASAP7_75t_R _20944_ (.A1(net346),
    .A2(_15573_),
    .B(_15574_),
    .C(net369),
    .Y(_15575_));
 BUFx2_ASAP7_75t_R input47 (.A(net3907),
    .Y(net47));
 INVx1_ASAP7_75t_R _20946_ (.A(_00713_),
    .Y(_15577_));
 NAND2x1_ASAP7_75t_R _20947_ (.A(net346),
    .B(_00711_),
    .Y(_15578_));
 OA211x2_ASAP7_75t_R _20948_ (.A1(net346),
    .A2(_15577_),
    .B(_15578_),
    .C(net325),
    .Y(_15579_));
 OR3x1_ASAP7_75t_R _20949_ (.A(_13350_),
    .B(_15575_),
    .C(_15579_),
    .Y(_15580_));
 INVx1_ASAP7_75t_R _20950_ (.A(_00717_),
    .Y(_15581_));
 NAND2x1_ASAP7_75t_R _20951_ (.A(net346),
    .B(_00715_),
    .Y(_15582_));
 OA211x2_ASAP7_75t_R _20952_ (.A1(net346),
    .A2(_15581_),
    .B(_15582_),
    .C(net325),
    .Y(_15583_));
 INVx1_ASAP7_75t_R _20953_ (.A(_00716_),
    .Y(_15584_));
 NAND2x1_ASAP7_75t_R _20954_ (.A(net348),
    .B(_00714_),
    .Y(_15585_));
 OA211x2_ASAP7_75t_R _20955_ (.A1(net348),
    .A2(_15584_),
    .B(_15585_),
    .C(net369),
    .Y(_15586_));
 OR3x1_ASAP7_75t_R _20956_ (.A(net337),
    .B(_15583_),
    .C(_15586_),
    .Y(_15587_));
 AND3x1_ASAP7_75t_R _20957_ (.A(_13373_),
    .B(_15580_),
    .C(_15587_),
    .Y(_15588_));
 OR3x1_ASAP7_75t_R _20958_ (.A(net328),
    .B(_15572_),
    .C(_15588_),
    .Y(_15589_));
 OAI21x1_ASAP7_75t_R _20959_ (.A1(_13355_),
    .A2(_15547_),
    .B(_15589_),
    .Y(_15590_));
 OA21x2_ASAP7_75t_R _20960_ (.A1(_00282_),
    .A2(_15490_),
    .B(_15492_),
    .Y(_15591_));
 AOI21x1_ASAP7_75t_R _20961_ (.A1(_13474_),
    .A2(_15590_),
    .B(_15591_),
    .Y(_18389_));
 XOR2x1_ASAP7_75t_R _20962_ (.A(_13620_),
    .Y(_15592_),
    .B(_18389_));
 NOR2x1_ASAP7_75t_R _20963_ (.A(_13986_),
    .B(_15590_),
    .Y(_15593_));
 NAND2x1_ASAP7_75t_R _20964_ (.A(net413),
    .B(_00703_),
    .Y(_15594_));
 OA211x2_ASAP7_75t_R _20965_ (.A1(net413),
    .A2(_15551_),
    .B(_15594_),
    .C(_13649_),
    .Y(_15595_));
 NAND2x1_ASAP7_75t_R _20966_ (.A(net413),
    .B(_00702_),
    .Y(_15596_));
 OA211x2_ASAP7_75t_R _20967_ (.A1(net413),
    .A2(_15557_),
    .B(_15596_),
    .C(net426),
    .Y(_15597_));
 OR3x1_ASAP7_75t_R _20968_ (.A(net321),
    .B(_15595_),
    .C(_15597_),
    .Y(_15598_));
 NAND2x1_ASAP7_75t_R _20969_ (.A(net415),
    .B(_00707_),
    .Y(_15599_));
 OA211x2_ASAP7_75t_R _20970_ (.A1(net415),
    .A2(_15564_),
    .B(_15599_),
    .C(_13649_),
    .Y(_15600_));
 NAND2x1_ASAP7_75t_R _20971_ (.A(net415),
    .B(_00706_),
    .Y(_15601_));
 OA211x2_ASAP7_75t_R _20972_ (.A1(net415),
    .A2(_15567_),
    .B(_15601_),
    .C(net426),
    .Y(_15602_));
 OR3x1_ASAP7_75t_R _20973_ (.A(net387),
    .B(_15600_),
    .C(_15602_),
    .Y(_15603_));
 NAND2x1_ASAP7_75t_R _20974_ (.A(net415),
    .B(_00690_),
    .Y(_15604_));
 OA211x2_ASAP7_75t_R _20975_ (.A1(net415),
    .A2(_15523_),
    .B(_15604_),
    .C(net426),
    .Y(_15605_));
 BUFx2_ASAP7_75t_R input46 (.A(net4003),
    .Y(net46));
 NAND2x1_ASAP7_75t_R _20977_ (.A(net415),
    .B(_00691_),
    .Y(_15607_));
 OA211x2_ASAP7_75t_R _20978_ (.A1(net415),
    .A2(_15518_),
    .B(_15607_),
    .C(_13649_),
    .Y(_15608_));
 OR3x1_ASAP7_75t_R _20979_ (.A(_14015_),
    .B(_15605_),
    .C(_15608_),
    .Y(_15609_));
 INVx1_ASAP7_75t_R _20980_ (.A(_00689_),
    .Y(_15610_));
 NAND2x1_ASAP7_75t_R _20981_ (.A(net413),
    .B(_01696_),
    .Y(_15611_));
 OA211x2_ASAP7_75t_R _20982_ (.A1(net413),
    .A2(_15610_),
    .B(_15611_),
    .C(net319),
    .Y(_15612_));
 NOR2x1_ASAP7_75t_R _20983_ (.A(net413),
    .B(_00688_),
    .Y(_15613_));
 AO21x1_ASAP7_75t_R _20984_ (.A1(net426),
    .A2(_15613_),
    .B(net315),
    .Y(_15614_));
 OA21x2_ASAP7_75t_R _20985_ (.A1(_15612_),
    .A2(_15614_),
    .B(net378),
    .Y(_15615_));
 AO32x1_ASAP7_75t_R _20986_ (.A1(_13626_),
    .A2(_15598_),
    .A3(_15603_),
    .B1(_15609_),
    .B2(_15615_),
    .Y(_15616_));
 NOR2x1_ASAP7_75t_R _20987_ (.A(net415),
    .B(_00700_),
    .Y(_15617_));
 AO21x1_ASAP7_75t_R _20988_ (.A1(net415),
    .A2(_15505_),
    .B(_15617_),
    .Y(_15618_));
 NAND2x1_ASAP7_75t_R _20989_ (.A(net415),
    .B(_00699_),
    .Y(_15619_));
 OA211x2_ASAP7_75t_R _20990_ (.A1(net415),
    .A2(_15510_),
    .B(_15619_),
    .C(_13649_),
    .Y(_15620_));
 AO21x1_ASAP7_75t_R _20991_ (.A1(net426),
    .A2(_15618_),
    .B(_15620_),
    .Y(_15621_));
 BUFx2_ASAP7_75t_R input45 (.A(net3970),
    .Y(net45));
 BUFx2_ASAP7_75t_R input44 (.A(net3998),
    .Y(net44));
 NAND2x1_ASAP7_75t_R _20994_ (.A(net415),
    .B(_00695_),
    .Y(_15624_));
 OA211x2_ASAP7_75t_R _20995_ (.A1(net415),
    .A2(_15537_),
    .B(_15624_),
    .C(_13649_),
    .Y(_15625_));
 NAND2x1_ASAP7_75t_R _20996_ (.A(net415),
    .B(_00694_),
    .Y(_15626_));
 OA211x2_ASAP7_75t_R _20997_ (.A1(net415),
    .A2(_15541_),
    .B(_15626_),
    .C(net426),
    .Y(_15627_));
 OA21x2_ASAP7_75t_R _20998_ (.A1(_15625_),
    .A2(_15627_),
    .B(net387),
    .Y(_15628_));
 AO21x1_ASAP7_75t_R _20999_ (.A1(net321),
    .A2(_15621_),
    .B(_15628_),
    .Y(_15629_));
 AND2x2_ASAP7_75t_R _21000_ (.A(_15609_),
    .B(_15615_),
    .Y(_15630_));
 BUFx2_ASAP7_75t_R input43 (.A(net3940),
    .Y(net43));
 NAND2x1_ASAP7_75t_R _21002_ (.A(net413),
    .B(_00715_),
    .Y(_15632_));
 OA211x2_ASAP7_75t_R _21003_ (.A1(net413),
    .A2(_15581_),
    .B(_15632_),
    .C(_13649_),
    .Y(_15633_));
 NAND2x1_ASAP7_75t_R _21004_ (.A(net413),
    .B(_00714_),
    .Y(_15634_));
 OA211x2_ASAP7_75t_R _21005_ (.A1(net413),
    .A2(_15584_),
    .B(_15634_),
    .C(net426),
    .Y(_15635_));
 OR3x1_ASAP7_75t_R _21006_ (.A(net387),
    .B(_15633_),
    .C(_15635_),
    .Y(_15636_));
 NAND2x1_ASAP7_75t_R _21007_ (.A(net413),
    .B(_00711_),
    .Y(_15637_));
 OA211x2_ASAP7_75t_R _21008_ (.A1(net413),
    .A2(_15577_),
    .B(_15637_),
    .C(net319),
    .Y(_15638_));
 NAND2x1_ASAP7_75t_R _21009_ (.A(net413),
    .B(_00710_),
    .Y(_15639_));
 OA211x2_ASAP7_75t_R _21010_ (.A1(net413),
    .A2(_15573_),
    .B(_15639_),
    .C(net426),
    .Y(_15640_));
 OR3x1_ASAP7_75t_R _21011_ (.A(net321),
    .B(_15638_),
    .C(_15640_),
    .Y(_15641_));
 AND3x1_ASAP7_75t_R _21012_ (.A(_14780_),
    .B(_15636_),
    .C(_15641_),
    .Y(_15642_));
 AO221x2_ASAP7_75t_R _21013_ (.A1(net382),
    .A2(_15616_),
    .B1(_15629_),
    .B2(_15630_),
    .C(_15642_),
    .Y(_15643_));
 BUFx2_ASAP7_75t_R input42 (.A(net3932),
    .Y(net42));
 AOI22x1_ASAP7_75t_R _21015_ (.A1(_13775_),
    .A2(_00718_),
    .B1(_02220_),
    .B2(_13778_),
    .Y(_15645_));
 OA211x2_ASAP7_75t_R _21016_ (.A1(_00284_),
    .A2(_15643_),
    .B(_15645_),
    .C(_13986_),
    .Y(_15646_));
 OA21x2_ASAP7_75t_R _21017_ (.A1(_15593_),
    .A2(_15646_),
    .B(_13817_),
    .Y(_15647_));
 AOI21x1_ASAP7_75t_R _21018_ (.A1(net309),
    .A2(_15592_),
    .B(_15647_),
    .Y(_17779_));
 INVx1_ASAP7_75t_R _21019_ (.A(_17779_),
    .Y(_16738_));
 INVx2_ASAP7_75t_R _21020_ (.A(_00201_),
    .Y(\cs_registers_i.pc_id_i[13] ));
 OA21x2_ASAP7_75t_R _21021_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_13808_),
    .B(_13794_),
    .Y(_15648_));
 INVx1_ASAP7_75t_R _21022_ (.A(_01628_),
    .Y(_15649_));
 AO32x1_ASAP7_75t_R _21023_ (.A1(\cs_registers_i.pc_id_i[13] ),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_15649_),
    .B2(_13450_),
    .Y(_15650_));
 AOI21x1_ASAP7_75t_R _21024_ (.A1(_15643_),
    .A2(_15648_),
    .B(_15650_),
    .Y(_18390_));
 OA21x2_ASAP7_75t_R _21025_ (.A1(_00718_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_15651_));
 AOI21x1_ASAP7_75t_R _21026_ (.A1(net309),
    .A2(_18390_),
    .B(_15651_),
    .Y(_17778_));
 INVx1_ASAP7_75t_R _21027_ (.A(_17778_),
    .Y(_16737_));
 OR4x2_ASAP7_75t_R _21028_ (.A(_00681_),
    .B(_00685_),
    .C(_02270_),
    .D(_02272_),
    .Y(_15652_));
 OA21x2_ASAP7_75t_R _21029_ (.A1(_00683_),
    .A2(_02270_),
    .B(_02269_),
    .Y(_15653_));
 OR3x1_ASAP7_75t_R _21030_ (.A(_00685_),
    .B(_02272_),
    .C(_15653_),
    .Y(_15654_));
 OA21x2_ASAP7_75t_R _21031_ (.A1(_00687_),
    .A2(_02272_),
    .B(_02271_),
    .Y(_15655_));
 OA211x2_ASAP7_75t_R _21032_ (.A1(_15340_),
    .A2(_15652_),
    .B(_15654_),
    .C(_15655_),
    .Y(_15656_));
 OA21x2_ASAP7_75t_R _21033_ (.A1(_15344_),
    .A2(_15652_),
    .B(_15656_),
    .Y(_16739_));
 BUFx2_ASAP7_75t_R input41 (.A(net4043),
    .Y(net41));
 BUFx2_ASAP7_75t_R input40 (.A(net4018),
    .Y(net40));
 AND2x2_ASAP7_75t_R _21036_ (.A(net350),
    .B(_01695_),
    .Y(_15659_));
 AO21x1_ASAP7_75t_R _21037_ (.A1(_13359_),
    .A2(_00721_),
    .B(_15659_),
    .Y(_15660_));
 OAI22x1_ASAP7_75t_R _21038_ (.A1(_00720_),
    .A2(net311),
    .B1(_15660_),
    .B2(net373),
    .Y(_15661_));
 BUFx2_ASAP7_75t_R input39 (.A(net3924),
    .Y(net39));
 INVx1_ASAP7_75t_R _21040_ (.A(_00729_),
    .Y(_15663_));
 NAND2x1_ASAP7_75t_R _21041_ (.A(net350),
    .B(_00727_),
    .Y(_15664_));
 OA211x2_ASAP7_75t_R _21042_ (.A1(net350),
    .A2(_15663_),
    .B(_15664_),
    .C(net324),
    .Y(_15665_));
 INVx1_ASAP7_75t_R _21043_ (.A(_00728_),
    .Y(_15666_));
 BUFx2_ASAP7_75t_R input38 (.A(net3786),
    .Y(net38));
 NAND2x1_ASAP7_75t_R _21045_ (.A(net350),
    .B(_00726_),
    .Y(_15668_));
 OA211x2_ASAP7_75t_R _21046_ (.A1(net350),
    .A2(_15666_),
    .B(_15668_),
    .C(net373),
    .Y(_15669_));
 OR3x1_ASAP7_75t_R _21047_ (.A(net330),
    .B(_15665_),
    .C(_15669_),
    .Y(_15670_));
 OA21x2_ASAP7_75t_R _21048_ (.A1(_13373_),
    .A2(_15661_),
    .B(_15670_),
    .Y(_15671_));
 BUFx2_ASAP7_75t_R input37 (.A(net4058),
    .Y(net37));
 BUFx2_ASAP7_75t_R input36 (.A(net4013),
    .Y(net36));
 INVx1_ASAP7_75t_R _21051_ (.A(_00725_),
    .Y(_15674_));
 BUFx2_ASAP7_75t_R input35 (.A(net4048),
    .Y(net35));
 NAND2x1_ASAP7_75t_R _21053_ (.A(net349),
    .B(_00723_),
    .Y(_15676_));
 OA211x2_ASAP7_75t_R _21054_ (.A1(net349),
    .A2(_15674_),
    .B(_15676_),
    .C(net324),
    .Y(_15677_));
 BUFx2_ASAP7_75t_R input34 (.A(net4023),
    .Y(net34));
 INVx1_ASAP7_75t_R _21056_ (.A(_00724_),
    .Y(_15679_));
 NAND2x1_ASAP7_75t_R _21057_ (.A(net349),
    .B(_00722_),
    .Y(_15680_));
 OA211x2_ASAP7_75t_R _21058_ (.A1(net349),
    .A2(_15679_),
    .B(_15680_),
    .C(net369),
    .Y(_15681_));
 OR3x1_ASAP7_75t_R _21059_ (.A(_13373_),
    .B(_15677_),
    .C(_15681_),
    .Y(_15682_));
 INVx1_ASAP7_75t_R _21060_ (.A(_00733_),
    .Y(_15683_));
 NAND2x1_ASAP7_75t_R _21061_ (.A(net349),
    .B(_00731_),
    .Y(_15684_));
 OA211x2_ASAP7_75t_R _21062_ (.A1(net349),
    .A2(_15683_),
    .B(_15684_),
    .C(net325),
    .Y(_15685_));
 INVx1_ASAP7_75t_R _21063_ (.A(_00732_),
    .Y(_15686_));
 NAND2x1_ASAP7_75t_R _21064_ (.A(net349),
    .B(_00730_),
    .Y(_15687_));
 OA211x2_ASAP7_75t_R _21065_ (.A1(net349),
    .A2(_15686_),
    .B(_15687_),
    .C(net369),
    .Y(_15688_));
 OR3x1_ASAP7_75t_R _21066_ (.A(net331),
    .B(_15685_),
    .C(_15688_),
    .Y(_15689_));
 AO21x1_ASAP7_75t_R _21067_ (.A1(_15682_),
    .A2(_15689_),
    .B(net335),
    .Y(_15690_));
 OA211x2_ASAP7_75t_R _21068_ (.A1(_13350_),
    .A2(_15671_),
    .B(_15690_),
    .C(net327),
    .Y(_15691_));
 INVx1_ASAP7_75t_R _21069_ (.A(_00741_),
    .Y(_15692_));
 NAND2x1_ASAP7_75t_R _21070_ (.A(net349),
    .B(_00739_),
    .Y(_15693_));
 OA211x2_ASAP7_75t_R _21071_ (.A1(net349),
    .A2(_15692_),
    .B(_15693_),
    .C(net324),
    .Y(_15694_));
 INVx1_ASAP7_75t_R _21072_ (.A(_00740_),
    .Y(_15695_));
 NAND2x1_ASAP7_75t_R _21073_ (.A(net349),
    .B(_00738_),
    .Y(_15696_));
 OA211x2_ASAP7_75t_R _21074_ (.A1(net349),
    .A2(_15695_),
    .B(_15696_),
    .C(net369),
    .Y(_15697_));
 OR3x1_ASAP7_75t_R _21075_ (.A(net335),
    .B(_15694_),
    .C(_15697_),
    .Y(_15698_));
 INVx1_ASAP7_75t_R _21076_ (.A(_00737_),
    .Y(_15699_));
 NAND2x1_ASAP7_75t_R _21077_ (.A(net349),
    .B(_00735_),
    .Y(_15700_));
 OA211x2_ASAP7_75t_R _21078_ (.A1(net349),
    .A2(_15699_),
    .B(_15700_),
    .C(net324),
    .Y(_15701_));
 INVx1_ASAP7_75t_R _21079_ (.A(_00736_),
    .Y(_15702_));
 NAND2x1_ASAP7_75t_R _21080_ (.A(net349),
    .B(_00734_),
    .Y(_15703_));
 OA211x2_ASAP7_75t_R _21081_ (.A1(net349),
    .A2(_15702_),
    .B(_15703_),
    .C(net369),
    .Y(_15704_));
 OR3x1_ASAP7_75t_R _21082_ (.A(_13350_),
    .B(_15701_),
    .C(_15704_),
    .Y(_15705_));
 AND3x1_ASAP7_75t_R _21083_ (.A(net330),
    .B(_15698_),
    .C(_15705_),
    .Y(_15706_));
 INVx1_ASAP7_75t_R _21084_ (.A(_00744_),
    .Y(_15707_));
 NAND2x1_ASAP7_75t_R _21085_ (.A(net350),
    .B(_00742_),
    .Y(_15708_));
 OA211x2_ASAP7_75t_R _21086_ (.A1(net350),
    .A2(_15707_),
    .B(_15708_),
    .C(net373),
    .Y(_15709_));
 INVx1_ASAP7_75t_R _21087_ (.A(_00745_),
    .Y(_15710_));
 NAND2x1_ASAP7_75t_R _21088_ (.A(net350),
    .B(_00743_),
    .Y(_15711_));
 OA211x2_ASAP7_75t_R _21089_ (.A1(net350),
    .A2(_15710_),
    .B(_15711_),
    .C(net324),
    .Y(_15712_));
 OR3x1_ASAP7_75t_R _21090_ (.A(_13350_),
    .B(_15709_),
    .C(_15712_),
    .Y(_15713_));
 INVx1_ASAP7_75t_R _21091_ (.A(_00749_),
    .Y(_15714_));
 NAND2x1_ASAP7_75t_R _21092_ (.A(net350),
    .B(_00747_),
    .Y(_15715_));
 OA211x2_ASAP7_75t_R _21093_ (.A1(net350),
    .A2(_15714_),
    .B(_15715_),
    .C(net324),
    .Y(_15716_));
 INVx1_ASAP7_75t_R _21094_ (.A(_00748_),
    .Y(_15717_));
 NAND2x1_ASAP7_75t_R _21095_ (.A(net349),
    .B(_00746_),
    .Y(_15718_));
 OA211x2_ASAP7_75t_R _21096_ (.A1(net349),
    .A2(_15717_),
    .B(_15718_),
    .C(net369),
    .Y(_15719_));
 OR3x1_ASAP7_75t_R _21097_ (.A(net335),
    .B(_15716_),
    .C(_15719_),
    .Y(_15720_));
 AND3x1_ASAP7_75t_R _21098_ (.A(_13373_),
    .B(_15713_),
    .C(_15720_),
    .Y(_15721_));
 OA21x2_ASAP7_75t_R _21099_ (.A1(_15706_),
    .A2(_15721_),
    .B(_13355_),
    .Y(_15722_));
 NOR2x2_ASAP7_75t_R _21100_ (.A(_15691_),
    .B(_15722_),
    .Y(_15723_));
 OA21x2_ASAP7_75t_R _21101_ (.A1(_00279_),
    .A2(_15490_),
    .B(_15492_),
    .Y(_15724_));
 AO21x1_ASAP7_75t_R _21102_ (.A1(_13474_),
    .A2(_15723_),
    .B(_15724_),
    .Y(_18393_));
 INVx1_ASAP7_75t_R _21103_ (.A(_18393_),
    .Y(_18395_));
 NAND2x1_ASAP7_75t_R _21104_ (.A(net395),
    .B(_00735_),
    .Y(_15725_));
 OA211x2_ASAP7_75t_R _21105_ (.A1(net395),
    .A2(_15699_),
    .B(_15725_),
    .C(net317),
    .Y(_15726_));
 NAND2x1_ASAP7_75t_R _21106_ (.A(net395),
    .B(_00734_),
    .Y(_15727_));
 OA211x2_ASAP7_75t_R _21107_ (.A1(net395),
    .A2(_15702_),
    .B(_15727_),
    .C(net423),
    .Y(_15728_));
 OR3x1_ASAP7_75t_R _21108_ (.A(net321),
    .B(_15726_),
    .C(_15728_),
    .Y(_15729_));
 NAND2x1_ASAP7_75t_R _21109_ (.A(net395),
    .B(_00739_),
    .Y(_15730_));
 OA211x2_ASAP7_75t_R _21110_ (.A1(net395),
    .A2(_15692_),
    .B(_15730_),
    .C(net317),
    .Y(_15731_));
 NAND2x1_ASAP7_75t_R _21111_ (.A(net395),
    .B(_00738_),
    .Y(_15732_));
 OA211x2_ASAP7_75t_R _21112_ (.A1(net395),
    .A2(_15695_),
    .B(_15732_),
    .C(net423),
    .Y(_15733_));
 OR3x1_ASAP7_75t_R _21113_ (.A(net385),
    .B(_15731_),
    .C(_15733_),
    .Y(_15734_));
 NAND2x1_ASAP7_75t_R _21114_ (.A(net395),
    .B(_00723_),
    .Y(_15735_));
 OA211x2_ASAP7_75t_R _21115_ (.A1(net395),
    .A2(_15674_),
    .B(_15735_),
    .C(net317),
    .Y(_15736_));
 NAND2x1_ASAP7_75t_R _21116_ (.A(net395),
    .B(_00722_),
    .Y(_15737_));
 OA211x2_ASAP7_75t_R _21117_ (.A1(net395),
    .A2(_15679_),
    .B(_15737_),
    .C(net423),
    .Y(_15738_));
 OR3x1_ASAP7_75t_R _21118_ (.A(net312),
    .B(_15736_),
    .C(_15738_),
    .Y(_15739_));
 INVx1_ASAP7_75t_R _21119_ (.A(_00721_),
    .Y(_15740_));
 NAND2x1_ASAP7_75t_R _21120_ (.A(net407),
    .B(_01695_),
    .Y(_15741_));
 OA211x2_ASAP7_75t_R _21121_ (.A1(net407),
    .A2(_15740_),
    .B(_15741_),
    .C(net317),
    .Y(_15742_));
 NOR2x1_ASAP7_75t_R _21122_ (.A(net407),
    .B(_00720_),
    .Y(_15743_));
 AO21x1_ASAP7_75t_R _21123_ (.A1(net423),
    .A2(_15743_),
    .B(_14005_),
    .Y(_15744_));
 OA21x2_ASAP7_75t_R _21124_ (.A1(_15742_),
    .A2(_15744_),
    .B(net377),
    .Y(_15745_));
 AO32x1_ASAP7_75t_R _21125_ (.A1(_13626_),
    .A2(_15729_),
    .A3(_15734_),
    .B1(_15739_),
    .B2(_15745_),
    .Y(_15746_));
 NAND2x1_ASAP7_75t_R _21126_ (.A(net395),
    .B(_00731_),
    .Y(_15747_));
 OA211x2_ASAP7_75t_R _21127_ (.A1(net395),
    .A2(_15683_),
    .B(_15747_),
    .C(_13649_),
    .Y(_15748_));
 NAND2x1_ASAP7_75t_R _21128_ (.A(net395),
    .B(_00730_),
    .Y(_15749_));
 OA211x2_ASAP7_75t_R _21129_ (.A1(net395),
    .A2(_15686_),
    .B(_15749_),
    .C(net423),
    .Y(_15750_));
 OR3x1_ASAP7_75t_R _21130_ (.A(net386),
    .B(_15748_),
    .C(_15750_),
    .Y(_15751_));
 NAND2x1_ASAP7_75t_R _21131_ (.A(net396),
    .B(_00727_),
    .Y(_15752_));
 OA211x2_ASAP7_75t_R _21132_ (.A1(net396),
    .A2(_15663_),
    .B(_15752_),
    .C(net317),
    .Y(_15753_));
 NAND2x1_ASAP7_75t_R _21133_ (.A(net407),
    .B(_00726_),
    .Y(_15754_));
 OA211x2_ASAP7_75t_R _21134_ (.A1(net407),
    .A2(_15666_),
    .B(_15754_),
    .C(net423),
    .Y(_15755_));
 OR3x1_ASAP7_75t_R _21135_ (.A(net321),
    .B(_15753_),
    .C(_15755_),
    .Y(_15756_));
 AND2x2_ASAP7_75t_R _21136_ (.A(_15751_),
    .B(_15756_),
    .Y(_15757_));
 AND2x2_ASAP7_75t_R _21137_ (.A(_15739_),
    .B(_15745_),
    .Y(_15758_));
 BUFx2_ASAP7_75t_R input33 (.A(net4053),
    .Y(net33));
 INVx1_ASAP7_75t_R _21139_ (.A(_00742_),
    .Y(_15760_));
 NOR2x1_ASAP7_75t_R _21140_ (.A(net385),
    .B(_00746_),
    .Y(_15761_));
 AO21x1_ASAP7_75t_R _21141_ (.A1(net385),
    .A2(_15760_),
    .B(_15761_),
    .Y(_15762_));
 INVx1_ASAP7_75t_R _21142_ (.A(_00747_),
    .Y(_15763_));
 NAND2x1_ASAP7_75t_R _21143_ (.A(net385),
    .B(_00743_),
    .Y(_15764_));
 OA211x2_ASAP7_75t_R _21144_ (.A1(net385),
    .A2(_15763_),
    .B(_15764_),
    .C(net317),
    .Y(_15765_));
 AO21x1_ASAP7_75t_R _21145_ (.A1(net423),
    .A2(_15762_),
    .B(_15765_),
    .Y(_15766_));
 NAND2x1_ASAP7_75t_R _21146_ (.A(net423),
    .B(_00744_),
    .Y(_15767_));
 OA211x2_ASAP7_75t_R _21147_ (.A1(net423),
    .A2(_15710_),
    .B(_15767_),
    .C(net385),
    .Y(_15768_));
 NAND2x1_ASAP7_75t_R _21148_ (.A(net423),
    .B(_00748_),
    .Y(_15769_));
 OA211x2_ASAP7_75t_R _21149_ (.A1(net423),
    .A2(_15714_),
    .B(_15769_),
    .C(net321),
    .Y(_15770_));
 OR3x1_ASAP7_75t_R _21150_ (.A(net407),
    .B(_15768_),
    .C(_15770_),
    .Y(_15771_));
 OA211x2_ASAP7_75t_R _21151_ (.A1(net316),
    .A2(_15766_),
    .B(_15771_),
    .C(_14780_),
    .Y(_15772_));
 AO221x2_ASAP7_75t_R _21152_ (.A1(net379),
    .A2(_15746_),
    .B1(_15757_),
    .B2(_15758_),
    .C(_15772_),
    .Y(_15773_));
 BUFx2_ASAP7_75t_R input32 (.A(net4008),
    .Y(net32));
 INVx2_ASAP7_75t_R _21154_ (.A(_00204_),
    .Y(_15775_));
 INVx1_ASAP7_75t_R _21155_ (.A(_01627_),
    .Y(_15776_));
 AO32x2_ASAP7_75t_R _21156_ (.A1(_15775_),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_15776_),
    .B2(_13450_),
    .Y(_15777_));
 AOI21x1_ASAP7_75t_R _21157_ (.A1(_13810_),
    .A2(_15773_),
    .B(_15777_),
    .Y(_18394_));
 XOR2x2_ASAP7_75t_R _21158_ (.A(_00751_),
    .B(_02227_),
    .Y(_15778_));
 INVx5_ASAP7_75t_R _21159_ (.A(_15778_),
    .Y(net155));
 BUFx2_ASAP7_75t_R input31 (.A(net3916),
    .Y(net31));
 AND2x2_ASAP7_75t_R _21161_ (.A(net342),
    .B(_01694_),
    .Y(_15780_));
 AO21x1_ASAP7_75t_R _21162_ (.A1(net2278),
    .A2(_00754_),
    .B(_15780_),
    .Y(_15781_));
 OAI22x1_ASAP7_75t_R _21163_ (.A1(_00753_),
    .A2(net311),
    .B1(_15781_),
    .B2(net376),
    .Y(_15782_));
 BUFx2_ASAP7_75t_R input30 (.A(net3976),
    .Y(net30));
 INVx1_ASAP7_75t_R _21165_ (.A(_00762_),
    .Y(_15784_));
 NAND2x1_ASAP7_75t_R _21166_ (.A(net343),
    .B(_00760_),
    .Y(_15785_));
 OA211x2_ASAP7_75t_R _21167_ (.A1(net343),
    .A2(_15784_),
    .B(_15785_),
    .C(_13376_),
    .Y(_15786_));
 INVx1_ASAP7_75t_R _21168_ (.A(_00761_),
    .Y(_15787_));
 NAND2x1_ASAP7_75t_R _21169_ (.A(net345),
    .B(_00759_),
    .Y(_15788_));
 OA211x2_ASAP7_75t_R _21170_ (.A1(net345),
    .A2(_15787_),
    .B(_15788_),
    .C(net376),
    .Y(_15789_));
 OR3x1_ASAP7_75t_R _21171_ (.A(net332),
    .B(_15786_),
    .C(_15789_),
    .Y(_15790_));
 OA211x2_ASAP7_75t_R _21172_ (.A1(_13373_),
    .A2(_15782_),
    .B(_15790_),
    .C(net338),
    .Y(_15791_));
 INVx1_ASAP7_75t_R _21173_ (.A(_00758_),
    .Y(_15792_));
 NAND2x1_ASAP7_75t_R _21174_ (.A(net344),
    .B(_00756_),
    .Y(_15793_));
 OA211x2_ASAP7_75t_R _21175_ (.A1(net344),
    .A2(_15792_),
    .B(_15793_),
    .C(_13376_),
    .Y(_15794_));
 INVx1_ASAP7_75t_R _21176_ (.A(_00757_),
    .Y(_15795_));
 NAND2x1_ASAP7_75t_R _21177_ (.A(net344),
    .B(_00755_),
    .Y(_15796_));
 OA211x2_ASAP7_75t_R _21178_ (.A1(net344),
    .A2(_15795_),
    .B(_15796_),
    .C(net2313),
    .Y(_15797_));
 OR3x1_ASAP7_75t_R _21179_ (.A(_13373_),
    .B(_15794_),
    .C(_15797_),
    .Y(_15798_));
 INVx1_ASAP7_75t_R _21180_ (.A(_00766_),
    .Y(_15799_));
 NAND2x1_ASAP7_75t_R _21181_ (.A(net344),
    .B(_00764_),
    .Y(_15800_));
 OA211x2_ASAP7_75t_R _21182_ (.A1(net344),
    .A2(_15799_),
    .B(_15800_),
    .C(_13376_),
    .Y(_15801_));
 INVx1_ASAP7_75t_R _21183_ (.A(_00765_),
    .Y(_15802_));
 NAND2x1_ASAP7_75t_R _21184_ (.A(net344),
    .B(_00763_),
    .Y(_15803_));
 OA211x2_ASAP7_75t_R _21185_ (.A1(net344),
    .A2(_15802_),
    .B(_15803_),
    .C(net2315),
    .Y(_15804_));
 OR3x1_ASAP7_75t_R _21186_ (.A(_00245_),
    .B(_15801_),
    .C(_15804_),
    .Y(_15805_));
 AND3x1_ASAP7_75t_R _21187_ (.A(_13350_),
    .B(_15798_),
    .C(_15805_),
    .Y(_15806_));
 OR3x4_ASAP7_75t_R _21188_ (.A(_13355_),
    .B(_15791_),
    .C(_15806_),
    .Y(_15807_));
 INVx1_ASAP7_75t_R _21189_ (.A(_00770_),
    .Y(_15808_));
 NAND2x1_ASAP7_75t_R _21190_ (.A(net341),
    .B(_00768_),
    .Y(_15809_));
 OA211x2_ASAP7_75t_R _21191_ (.A1(net341),
    .A2(_15808_),
    .B(_15809_),
    .C(net323),
    .Y(_15810_));
 INVx1_ASAP7_75t_R _21192_ (.A(_00769_),
    .Y(_15811_));
 NAND2x1_ASAP7_75t_R _21193_ (.A(net341),
    .B(_00767_),
    .Y(_15812_));
 OA211x2_ASAP7_75t_R _21194_ (.A1(net341),
    .A2(_15811_),
    .B(_15812_),
    .C(net370),
    .Y(_15813_));
 OR3x1_ASAP7_75t_R _21195_ (.A(_13350_),
    .B(_15810_),
    .C(_15813_),
    .Y(_15814_));
 INVx1_ASAP7_75t_R _21196_ (.A(_00774_),
    .Y(_15815_));
 NAND2x1_ASAP7_75t_R _21197_ (.A(net341),
    .B(_00772_),
    .Y(_15816_));
 OA211x2_ASAP7_75t_R _21198_ (.A1(net341),
    .A2(_15815_),
    .B(_15816_),
    .C(net323),
    .Y(_15817_));
 INVx1_ASAP7_75t_R _21199_ (.A(_00773_),
    .Y(_15818_));
 NAND2x1_ASAP7_75t_R _21200_ (.A(net341),
    .B(_00771_),
    .Y(_15819_));
 OA211x2_ASAP7_75t_R _21201_ (.A1(net341),
    .A2(_15818_),
    .B(_15819_),
    .C(net370),
    .Y(_15820_));
 OR3x1_ASAP7_75t_R _21202_ (.A(net337),
    .B(_15817_),
    .C(_15820_),
    .Y(_15821_));
 AND3x1_ASAP7_75t_R _21203_ (.A(net332),
    .B(_15814_),
    .C(_15821_),
    .Y(_15822_));
 INVx1_ASAP7_75t_R _21204_ (.A(_00782_),
    .Y(_15823_));
 NAND2x1_ASAP7_75t_R _21205_ (.A(net344),
    .B(_00780_),
    .Y(_15824_));
 OA211x2_ASAP7_75t_R _21206_ (.A1(net344),
    .A2(_15823_),
    .B(_15824_),
    .C(_13376_),
    .Y(_15825_));
 INVx1_ASAP7_75t_R _21207_ (.A(_00781_),
    .Y(_15826_));
 NAND2x1_ASAP7_75t_R _21208_ (.A(net344),
    .B(_00779_),
    .Y(_15827_));
 OA211x2_ASAP7_75t_R _21209_ (.A1(net344),
    .A2(_15826_),
    .B(_15827_),
    .C(net2315),
    .Y(_15828_));
 OR3x1_ASAP7_75t_R _21210_ (.A(net338),
    .B(_15825_),
    .C(_15828_),
    .Y(_15829_));
 INVx1_ASAP7_75t_R _21211_ (.A(_00778_),
    .Y(_15830_));
 NAND2x1_ASAP7_75t_R _21212_ (.A(net368),
    .B(_00776_),
    .Y(_15831_));
 OA211x2_ASAP7_75t_R _21213_ (.A1(net368),
    .A2(_15830_),
    .B(_15831_),
    .C(_13376_),
    .Y(_15832_));
 INVx1_ASAP7_75t_R _21214_ (.A(_00777_),
    .Y(_15833_));
 NAND2x1_ASAP7_75t_R _21215_ (.A(net368),
    .B(_00775_),
    .Y(_15834_));
 OA211x2_ASAP7_75t_R _21216_ (.A1(net368),
    .A2(_15833_),
    .B(_15834_),
    .C(net2314),
    .Y(_15835_));
 OR3x1_ASAP7_75t_R _21217_ (.A(_13350_),
    .B(_15832_),
    .C(_15835_),
    .Y(_15836_));
 AND3x2_ASAP7_75t_R _21218_ (.A(_13373_),
    .B(_15829_),
    .C(_15836_),
    .Y(_15837_));
 OR3x4_ASAP7_75t_R _21219_ (.A(net328),
    .B(_15822_),
    .C(_15837_),
    .Y(_15838_));
 NAND2x2_ASAP7_75t_R _21220_ (.A(_15807_),
    .B(_15838_),
    .Y(_15839_));
 OA21x2_ASAP7_75t_R _21221_ (.A1(net422),
    .A2(_15490_),
    .B(_15492_),
    .Y(_15840_));
 AO21x2_ASAP7_75t_R _21222_ (.A1(_13474_),
    .A2(_15839_),
    .B(_15840_),
    .Y(_15841_));
 BUFx2_ASAP7_75t_R input29 (.A(net4028),
    .Y(net29));
 INVx1_ASAP7_75t_R _21224_ (.A(_15841_),
    .Y(_18399_));
 INVx1_ASAP7_75t_R _21225_ (.A(_00206_),
    .Y(\cs_registers_i.pc_id_i[15] ));
 NAND2x1_ASAP7_75t_R _21226_ (.A(_00206_),
    .B(_13993_),
    .Y(_15842_));
 NAND2x1_ASAP7_75t_R _21227_ (.A(net418),
    .B(_00756_),
    .Y(_15843_));
 OA211x2_ASAP7_75t_R _21228_ (.A1(net418),
    .A2(_15792_),
    .B(_15843_),
    .C(_13649_),
    .Y(_15844_));
 NAND2x1_ASAP7_75t_R _21229_ (.A(net418),
    .B(_00755_),
    .Y(_15845_));
 OA211x2_ASAP7_75t_R _21230_ (.A1(net418),
    .A2(_15795_),
    .B(_15845_),
    .C(net419),
    .Y(_15846_));
 OR3x1_ASAP7_75t_R _21231_ (.A(_13636_),
    .B(_15844_),
    .C(_15846_),
    .Y(_15847_));
 NAND2x1_ASAP7_75t_R _21232_ (.A(net418),
    .B(_00764_),
    .Y(_15848_));
 OA211x2_ASAP7_75t_R _21233_ (.A1(net418),
    .A2(_15799_),
    .B(_15848_),
    .C(_13649_),
    .Y(_15849_));
 NAND2x1_ASAP7_75t_R _21234_ (.A(net418),
    .B(_00763_),
    .Y(_15850_));
 OA211x2_ASAP7_75t_R _21235_ (.A1(net418),
    .A2(_15802_),
    .B(_15850_),
    .C(net419),
    .Y(_15851_));
 OR3x1_ASAP7_75t_R _21236_ (.A(net381),
    .B(_15849_),
    .C(_15851_),
    .Y(_15852_));
 AO21x1_ASAP7_75t_R _21237_ (.A1(_15847_),
    .A2(_15852_),
    .B(net388),
    .Y(_15853_));
 AND2x2_ASAP7_75t_R _21238_ (.A(net393),
    .B(_01694_),
    .Y(_15854_));
 AO21x1_ASAP7_75t_R _21239_ (.A1(_13675_),
    .A2(_00754_),
    .B(_15854_),
    .Y(_15855_));
 OAI22x1_ASAP7_75t_R _21240_ (.A1(_00753_),
    .A2(net2291),
    .B1(_15855_),
    .B2(net427),
    .Y(_15856_));
 NAND2x1_ASAP7_75t_R _21241_ (.A(net390),
    .B(_00760_),
    .Y(_15857_));
 OA211x2_ASAP7_75t_R _21242_ (.A1(net390),
    .A2(_15784_),
    .B(_15857_),
    .C(_13649_),
    .Y(_15858_));
 NAND2x1_ASAP7_75t_R _21243_ (.A(net391),
    .B(_00759_),
    .Y(_15859_));
 OA211x2_ASAP7_75t_R _21244_ (.A1(net393),
    .A2(_15787_),
    .B(_15859_),
    .C(net427),
    .Y(_15860_));
 OR3x1_ASAP7_75t_R _21245_ (.A(_14942_),
    .B(_15858_),
    .C(_15860_),
    .Y(_15861_));
 OA211x2_ASAP7_75t_R _21246_ (.A1(net315),
    .A2(_15856_),
    .B(_15861_),
    .C(_00286_),
    .Y(_15862_));
 NAND2x1_ASAP7_75t_R _21247_ (.A(net392),
    .B(_00776_),
    .Y(_15863_));
 OA211x2_ASAP7_75t_R _21248_ (.A1(net392),
    .A2(_15830_),
    .B(_15863_),
    .C(_13649_),
    .Y(_15864_));
 NAND2x1_ASAP7_75t_R _21249_ (.A(net392),
    .B(_00775_),
    .Y(_15865_));
 OA211x2_ASAP7_75t_R _21250_ (.A1(net392),
    .A2(_15833_),
    .B(_15865_),
    .C(net419),
    .Y(_15866_));
 OR3x1_ASAP7_75t_R _21251_ (.A(_13630_),
    .B(_15864_),
    .C(_15866_),
    .Y(_15867_));
 NAND2x1_ASAP7_75t_R _21252_ (.A(net392),
    .B(_00780_),
    .Y(_15868_));
 OA211x2_ASAP7_75t_R _21253_ (.A1(net392),
    .A2(_15823_),
    .B(_15868_),
    .C(_13649_),
    .Y(_15869_));
 NAND2x1_ASAP7_75t_R _21254_ (.A(net392),
    .B(_00779_),
    .Y(_15870_));
 OA211x2_ASAP7_75t_R _21255_ (.A1(net392),
    .A2(_15826_),
    .B(_15870_),
    .C(net419),
    .Y(_15871_));
 OR3x1_ASAP7_75t_R _21256_ (.A(net388),
    .B(_15869_),
    .C(_15871_),
    .Y(_15872_));
 AO21x1_ASAP7_75t_R _21257_ (.A1(_15867_),
    .A2(_15872_),
    .B(net381),
    .Y(_15873_));
 NAND2x1_ASAP7_75t_R _21258_ (.A(net417),
    .B(_00768_),
    .Y(_15874_));
 OA211x2_ASAP7_75t_R _21259_ (.A1(net417),
    .A2(_15808_),
    .B(_15874_),
    .C(net319),
    .Y(_15875_));
 NAND2x1_ASAP7_75t_R _21260_ (.A(net417),
    .B(_00767_),
    .Y(_15876_));
 OA211x2_ASAP7_75t_R _21261_ (.A1(net417),
    .A2(_15811_),
    .B(_15876_),
    .C(net426),
    .Y(_15877_));
 OR3x1_ASAP7_75t_R _21262_ (.A(net315),
    .B(_15875_),
    .C(_15877_),
    .Y(_15878_));
 NAND2x1_ASAP7_75t_R _21263_ (.A(net417),
    .B(_00772_),
    .Y(_15879_));
 OA211x2_ASAP7_75t_R _21264_ (.A1(net417),
    .A2(_15815_),
    .B(_15879_),
    .C(net319),
    .Y(_15880_));
 NAND2x1_ASAP7_75t_R _21265_ (.A(net417),
    .B(_00771_),
    .Y(_15881_));
 OA211x2_ASAP7_75t_R _21266_ (.A1(net417),
    .A2(_15818_),
    .B(_15881_),
    .C(net426),
    .Y(_15882_));
 OR3x1_ASAP7_75t_R _21267_ (.A(_14015_),
    .B(_15880_),
    .C(_15882_),
    .Y(_15883_));
 AND3x1_ASAP7_75t_R _21268_ (.A(_13626_),
    .B(_15878_),
    .C(_15883_),
    .Y(_15884_));
 AO221x2_ASAP7_75t_R _21269_ (.A1(_15853_),
    .A2(_15862_),
    .B1(_15873_),
    .B2(_15884_),
    .C(_13993_),
    .Y(_15885_));
 INVx1_ASAP7_75t_R _21270_ (.A(_01626_),
    .Y(_15886_));
 AO32x2_ASAP7_75t_R _21271_ (.A1(_13794_),
    .A2(_15842_),
    .A3(_15885_),
    .B1(_13450_),
    .B2(_15886_),
    .Y(_15887_));
 BUFx2_ASAP7_75t_R input28 (.A(net3993),
    .Y(net28));
 INVx2_ASAP7_75t_R _21273_ (.A(_15887_),
    .Y(_18400_));
 OR2x2_ASAP7_75t_R _21274_ (.A(_00719_),
    .B(_16739_),
    .Y(_15888_));
 OA21x2_ASAP7_75t_R _21275_ (.A1(_00751_),
    .A2(_00752_),
    .B(_02273_),
    .Y(_15889_));
 OA21x2_ASAP7_75t_R _21276_ (.A1(_00751_),
    .A2(_15888_),
    .B(_15889_),
    .Y(_15890_));
 INVx1_ASAP7_75t_R _21277_ (.A(_15890_),
    .Y(_16741_));
 CKINVDCx8_ASAP7_75t_R _21278_ (.A(net260),
    .Y(net156));
 BUFx2_ASAP7_75t_R input27 (.A(net3779),
    .Y(net27));
 AND2x2_ASAP7_75t_R _21280_ (.A(net363),
    .B(_01693_),
    .Y(_15892_));
 AO21x1_ASAP7_75t_R _21281_ (.A1(net2278),
    .A2(_00787_),
    .B(_15892_),
    .Y(_15893_));
 BUFx3_ASAP7_75t_R input26 (.A(net3048),
    .Y(net26));
 BUFx3_ASAP7_75t_R input25 (.A(net3729),
    .Y(net25));
 BUFx2_ASAP7_75t_R input24 (.A(net3434),
    .Y(net24));
 OAI22x1_ASAP7_75t_R _21285_ (.A1(_00786_),
    .A2(net311),
    .B1(_15893_),
    .B2(net373),
    .Y(_15897_));
 BUFx2_ASAP7_75t_R input23 (.A(net3418),
    .Y(net23));
 INVx1_ASAP7_75t_R _21287_ (.A(_00795_),
    .Y(_15899_));
 NAND2x1_ASAP7_75t_R _21288_ (.A(net363),
    .B(_00793_),
    .Y(_15900_));
 BUFx2_ASAP7_75t_R input22 (.A(net3264),
    .Y(net22));
 OA211x2_ASAP7_75t_R _21290_ (.A1(net2333),
    .A2(_15899_),
    .B(_15900_),
    .C(net325),
    .Y(_15902_));
 BUFx2_ASAP7_75t_R input21 (.A(net3257),
    .Y(net21));
 INVx1_ASAP7_75t_R _21292_ (.A(_00794_),
    .Y(_15904_));
 NAND2x1_ASAP7_75t_R _21293_ (.A(net363),
    .B(_00792_),
    .Y(_15905_));
 OA211x2_ASAP7_75t_R _21294_ (.A1(net2333),
    .A2(_15904_),
    .B(_15905_),
    .C(net372),
    .Y(_15906_));
 OR3x1_ASAP7_75t_R _21295_ (.A(net330),
    .B(_15902_),
    .C(_15906_),
    .Y(_15907_));
 BUFx2_ASAP7_75t_R input20 (.A(net3395),
    .Y(net20));
 OA211x2_ASAP7_75t_R _21297_ (.A1(_13373_),
    .A2(_15897_),
    .B(_15907_),
    .C(net335),
    .Y(_15909_));
 BUFx2_ASAP7_75t_R input19 (.A(net3241),
    .Y(net19));
 INVx1_ASAP7_75t_R _21299_ (.A(_00791_),
    .Y(_15911_));
 NAND2x1_ASAP7_75t_R _21300_ (.A(net351),
    .B(_00789_),
    .Y(_15912_));
 BUFx2_ASAP7_75t_R input18 (.A(net3324),
    .Y(net18));
 BUFx2_ASAP7_75t_R input17 (.A(net3348),
    .Y(net17));
 OA211x2_ASAP7_75t_R _21303_ (.A1(net351),
    .A2(_15911_),
    .B(_15912_),
    .C(net325),
    .Y(_15915_));
 BUFx2_ASAP7_75t_R input16 (.A(net3362),
    .Y(net16));
 INVx1_ASAP7_75t_R _21305_ (.A(_00790_),
    .Y(_15917_));
 BUFx2_ASAP7_75t_R input15 (.A(net3441),
    .Y(net15));
 NAND2x1_ASAP7_75t_R _21307_ (.A(net351),
    .B(_00788_),
    .Y(_15919_));
 BUFx2_ASAP7_75t_R input14 (.A(net3402),
    .Y(net14));
 OA211x2_ASAP7_75t_R _21309_ (.A1(net351),
    .A2(_15917_),
    .B(_15919_),
    .C(net373),
    .Y(_15921_));
 OR3x1_ASAP7_75t_R _21310_ (.A(_13373_),
    .B(_15915_),
    .C(_15921_),
    .Y(_15922_));
 BUFx2_ASAP7_75t_R input13 (.A(net3309),
    .Y(net13));
 INVx1_ASAP7_75t_R _21312_ (.A(_00799_),
    .Y(_15924_));
 BUFx2_ASAP7_75t_R input12 (.A(net3340),
    .Y(net12));
 NAND2x1_ASAP7_75t_R _21314_ (.A(net350),
    .B(_00797_),
    .Y(_15926_));
 OA211x2_ASAP7_75t_R _21315_ (.A1(net350),
    .A2(_15924_),
    .B(_15926_),
    .C(net325),
    .Y(_15927_));
 INVx1_ASAP7_75t_R _21316_ (.A(_00798_),
    .Y(_15928_));
 NAND2x1_ASAP7_75t_R _21317_ (.A(net350),
    .B(_00796_),
    .Y(_15929_));
 OA211x2_ASAP7_75t_R _21318_ (.A1(net350),
    .A2(_15928_),
    .B(_15929_),
    .C(net373),
    .Y(_15930_));
 OR3x1_ASAP7_75t_R _21319_ (.A(net330),
    .B(_15927_),
    .C(_15930_),
    .Y(_15931_));
 AND3x1_ASAP7_75t_R _21320_ (.A(_13350_),
    .B(_15922_),
    .C(_15931_),
    .Y(_15932_));
 OR3x2_ASAP7_75t_R _21321_ (.A(_13355_),
    .B(_15909_),
    .C(_15932_),
    .Y(_15933_));
 BUFx2_ASAP7_75t_R input11 (.A(net3272),
    .Y(net11));
 BUFx2_ASAP7_75t_R input10 (.A(net3426),
    .Y(net10));
 INVx1_ASAP7_75t_R _21324_ (.A(_00807_),
    .Y(_15936_));
 NAND2x1_ASAP7_75t_R _21325_ (.A(net350),
    .B(_00805_),
    .Y(_15937_));
 OA211x2_ASAP7_75t_R _21326_ (.A1(net350),
    .A2(_15936_),
    .B(_15937_),
    .C(net325),
    .Y(_15938_));
 INVx1_ASAP7_75t_R _21327_ (.A(_00806_),
    .Y(_15939_));
 NAND2x1_ASAP7_75t_R _21328_ (.A(net350),
    .B(_00804_),
    .Y(_15940_));
 OA211x2_ASAP7_75t_R _21329_ (.A1(net350),
    .A2(_15939_),
    .B(_15940_),
    .C(net373),
    .Y(_15941_));
 OR3x1_ASAP7_75t_R _21330_ (.A(_13373_),
    .B(_15938_),
    .C(_15941_),
    .Y(_15942_));
 INVx1_ASAP7_75t_R _21331_ (.A(_00815_),
    .Y(_15943_));
 NAND2x1_ASAP7_75t_R _21332_ (.A(net2374),
    .B(_00813_),
    .Y(_15944_));
 BUFx2_ASAP7_75t_R input9 (.A(net3332),
    .Y(net9));
 OA211x2_ASAP7_75t_R _21334_ (.A1(net2374),
    .A2(_15943_),
    .B(_15944_),
    .C(net325),
    .Y(_15946_));
 BUFx2_ASAP7_75t_R input8 (.A(net3464),
    .Y(net8));
 BUFx2_ASAP7_75t_R input7 (.A(net3316),
    .Y(net7));
 INVx1_ASAP7_75t_R _21337_ (.A(_00814_),
    .Y(_15949_));
 NAND2x1_ASAP7_75t_R _21338_ (.A(net2374),
    .B(_00812_),
    .Y(_15950_));
 BUFx2_ASAP7_75t_R input6 (.A(net3448),
    .Y(net6));
 OA211x2_ASAP7_75t_R _21340_ (.A1(net2374),
    .A2(_15949_),
    .B(_15950_),
    .C(net372),
    .Y(_15952_));
 OR3x1_ASAP7_75t_R _21341_ (.A(net330),
    .B(_15946_),
    .C(_15952_),
    .Y(_15953_));
 AND3x1_ASAP7_75t_R _21342_ (.A(_13350_),
    .B(_15942_),
    .C(_15953_),
    .Y(_15954_));
 INVx1_ASAP7_75t_R _21343_ (.A(_00803_),
    .Y(_15955_));
 NAND2x1_ASAP7_75t_R _21344_ (.A(net359),
    .B(_00801_),
    .Y(_15956_));
 OA211x2_ASAP7_75t_R _21345_ (.A1(net2332),
    .A2(_15955_),
    .B(_15956_),
    .C(net325),
    .Y(_15957_));
 BUFx2_ASAP7_75t_R input5 (.A(net3471),
    .Y(net5));
 INVx1_ASAP7_75t_R _21347_ (.A(_00802_),
    .Y(_15959_));
 NAND2x1_ASAP7_75t_R _21348_ (.A(net359),
    .B(_00800_),
    .Y(_15960_));
 OA211x2_ASAP7_75t_R _21349_ (.A1(net2332),
    .A2(_15959_),
    .B(_15960_),
    .C(net372),
    .Y(_15961_));
 OR3x1_ASAP7_75t_R _21350_ (.A(_13373_),
    .B(_15957_),
    .C(_15961_),
    .Y(_15962_));
 INVx1_ASAP7_75t_R _21351_ (.A(_00811_),
    .Y(_15963_));
 NAND2x1_ASAP7_75t_R _21352_ (.A(net2374),
    .B(_00809_),
    .Y(_15964_));
 OA211x2_ASAP7_75t_R _21353_ (.A1(net2333),
    .A2(_15963_),
    .B(_15964_),
    .C(net325),
    .Y(_15965_));
 INVx1_ASAP7_75t_R _21354_ (.A(_00810_),
    .Y(_15966_));
 NAND2x1_ASAP7_75t_R _21355_ (.A(net2374),
    .B(_00808_),
    .Y(_15967_));
 OA211x2_ASAP7_75t_R _21356_ (.A1(net2374),
    .A2(_15966_),
    .B(_15967_),
    .C(net372),
    .Y(_15968_));
 OR3x1_ASAP7_75t_R _21357_ (.A(net330),
    .B(_15965_),
    .C(_15968_),
    .Y(_15969_));
 AND3x1_ASAP7_75t_R _21358_ (.A(net335),
    .B(_15962_),
    .C(_15969_),
    .Y(_15970_));
 OR3x2_ASAP7_75t_R _21359_ (.A(net327),
    .B(_15954_),
    .C(_15970_),
    .Y(_15971_));
 NAND2x2_ASAP7_75t_R _21360_ (.A(_15933_),
    .B(_15971_),
    .Y(_15972_));
 OA21x2_ASAP7_75t_R _21361_ (.A1(net409),
    .A2(_15490_),
    .B(_15492_),
    .Y(_15973_));
 AOI21x1_ASAP7_75t_R _21362_ (.A1(_13474_),
    .A2(_15972_),
    .B(_15973_),
    .Y(_18405_));
 AND2x2_ASAP7_75t_R _21363_ (.A(net407),
    .B(_01693_),
    .Y(_15974_));
 AO21x1_ASAP7_75t_R _21364_ (.A1(net316),
    .A2(_00787_),
    .B(_15974_),
    .Y(_15975_));
 OAI22x1_ASAP7_75t_R _21365_ (.A1(_00786_),
    .A2(net2292),
    .B1(_15975_),
    .B2(net422),
    .Y(_15976_));
 NAND2x1_ASAP7_75t_R _21366_ (.A(net400),
    .B(_00801_),
    .Y(_15977_));
 OA211x2_ASAP7_75t_R _21367_ (.A1(net400),
    .A2(_15955_),
    .B(_15977_),
    .C(net317),
    .Y(_15978_));
 NAND2x1_ASAP7_75t_R _21368_ (.A(net400),
    .B(_00800_),
    .Y(_15979_));
 OA211x2_ASAP7_75t_R _21369_ (.A1(net400),
    .A2(_15959_),
    .B(_15979_),
    .C(net422),
    .Y(_15980_));
 OR3x1_ASAP7_75t_R _21370_ (.A(net377),
    .B(_15978_),
    .C(_15980_),
    .Y(_15981_));
 OA211x2_ASAP7_75t_R _21371_ (.A1(_13626_),
    .A2(_15976_),
    .B(_15981_),
    .C(net385),
    .Y(_15982_));
 NAND2x1_ASAP7_75t_R _21372_ (.A(net397),
    .B(_00789_),
    .Y(_15983_));
 OA211x2_ASAP7_75t_R _21373_ (.A1(net397),
    .A2(_15911_),
    .B(_15983_),
    .C(net318),
    .Y(_15984_));
 NAND2x1_ASAP7_75t_R _21374_ (.A(net397),
    .B(_00788_),
    .Y(_15985_));
 OA211x2_ASAP7_75t_R _21375_ (.A1(net397),
    .A2(_15917_),
    .B(_15985_),
    .C(net423),
    .Y(_15986_));
 OR3x1_ASAP7_75t_R _21376_ (.A(_13626_),
    .B(_15984_),
    .C(_15986_),
    .Y(_15987_));
 NAND2x1_ASAP7_75t_R _21377_ (.A(net397),
    .B(_00805_),
    .Y(_15988_));
 OA211x2_ASAP7_75t_R _21378_ (.A1(net397),
    .A2(_15936_),
    .B(_15988_),
    .C(net317),
    .Y(_15989_));
 NAND2x1_ASAP7_75t_R _21379_ (.A(net397),
    .B(_00804_),
    .Y(_15990_));
 OA211x2_ASAP7_75t_R _21380_ (.A1(net397),
    .A2(_15939_),
    .B(_15990_),
    .C(net423),
    .Y(_15991_));
 OR3x1_ASAP7_75t_R _21381_ (.A(net378),
    .B(_15989_),
    .C(_15991_),
    .Y(_15992_));
 AND3x1_ASAP7_75t_R _21382_ (.A(net320),
    .B(_15987_),
    .C(_15992_),
    .Y(_15993_));
 OR3x2_ASAP7_75t_R _21383_ (.A(_13636_),
    .B(_15982_),
    .C(_15993_),
    .Y(_15994_));
 NAND2x1_ASAP7_75t_R _21384_ (.A(net407),
    .B(_00797_),
    .Y(_15995_));
 OA211x2_ASAP7_75t_R _21385_ (.A1(net407),
    .A2(_15924_),
    .B(_15995_),
    .C(net377),
    .Y(_15996_));
 NAND2x1_ASAP7_75t_R _21386_ (.A(net401),
    .B(_00813_),
    .Y(_15997_));
 OA211x2_ASAP7_75t_R _21387_ (.A1(net401),
    .A2(_15943_),
    .B(_15997_),
    .C(_13626_),
    .Y(_15998_));
 OR3x1_ASAP7_75t_R _21388_ (.A(net422),
    .B(_15996_),
    .C(_15998_),
    .Y(_15999_));
 NAND2x1_ASAP7_75t_R _21389_ (.A(net407),
    .B(_00796_),
    .Y(_16000_));
 OA211x2_ASAP7_75t_R _21390_ (.A1(net407),
    .A2(_15928_),
    .B(_16000_),
    .C(net377),
    .Y(_16001_));
 NAND2x1_ASAP7_75t_R _21391_ (.A(net401),
    .B(_00812_),
    .Y(_16002_));
 OA211x2_ASAP7_75t_R _21392_ (.A1(net401),
    .A2(_15949_),
    .B(_16002_),
    .C(_13626_),
    .Y(_16003_));
 OR3x1_ASAP7_75t_R _21393_ (.A(net317),
    .B(_16001_),
    .C(_16003_),
    .Y(_16004_));
 AND3x1_ASAP7_75t_R _21394_ (.A(net321),
    .B(_15999_),
    .C(_16004_),
    .Y(_16005_));
 NAND2x1_ASAP7_75t_R _21395_ (.A(net401),
    .B(_00792_),
    .Y(_16006_));
 OA211x2_ASAP7_75t_R _21396_ (.A1(net401),
    .A2(_15904_),
    .B(_16006_),
    .C(net377),
    .Y(_16007_));
 NAND2x1_ASAP7_75t_R _21397_ (.A(net401),
    .B(_00808_),
    .Y(_16008_));
 OA211x2_ASAP7_75t_R _21398_ (.A1(net401),
    .A2(_15966_),
    .B(_16008_),
    .C(_13626_),
    .Y(_16009_));
 OR3x1_ASAP7_75t_R _21399_ (.A(net317),
    .B(_16007_),
    .C(_16009_),
    .Y(_16010_));
 NAND2x1_ASAP7_75t_R _21400_ (.A(net407),
    .B(_00793_),
    .Y(_16011_));
 OA211x2_ASAP7_75t_R _21401_ (.A1(net407),
    .A2(_15899_),
    .B(_16011_),
    .C(net377),
    .Y(_16012_));
 NAND2x1_ASAP7_75t_R _21402_ (.A(net401),
    .B(_00809_),
    .Y(_16013_));
 OA211x2_ASAP7_75t_R _21403_ (.A1(net401),
    .A2(_15963_),
    .B(_16013_),
    .C(_13626_),
    .Y(_16014_));
 OR3x1_ASAP7_75t_R _21404_ (.A(net422),
    .B(_16012_),
    .C(_16014_),
    .Y(_16015_));
 AND3x1_ASAP7_75t_R _21405_ (.A(net385),
    .B(_16010_),
    .C(_16015_),
    .Y(_16016_));
 OR3x4_ASAP7_75t_R _21406_ (.A(net379),
    .B(_16005_),
    .C(_16016_),
    .Y(_16017_));
 AND3x2_ASAP7_75t_R _21407_ (.A(_13810_),
    .B(_15994_),
    .C(_16017_),
    .Y(_16018_));
 OAI22x1_ASAP7_75t_R _21408_ (.A1(_01625_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00208_),
    .Y(_16019_));
 OR2x4_ASAP7_75t_R _21409_ (.A(_16018_),
    .B(_16019_),
    .Y(_16020_));
 BUFx2_ASAP7_75t_R input4 (.A(net3249),
    .Y(net4));
 INVx2_ASAP7_75t_R _21411_ (.A(_16020_),
    .Y(_18404_));
 AND2x2_ASAP7_75t_R _21412_ (.A(net358),
    .B(_01692_),
    .Y(_16021_));
 AO21x1_ASAP7_75t_R _21413_ (.A1(_13359_),
    .A2(_00820_),
    .B(_16021_),
    .Y(_16022_));
 OAI22x1_ASAP7_75t_R _21414_ (.A1(_00819_),
    .A2(_14184_),
    .B1(_16022_),
    .B2(net372),
    .Y(_16023_));
 INVx1_ASAP7_75t_R _21415_ (.A(_00828_),
    .Y(_16024_));
 NAND2x1_ASAP7_75t_R _21416_ (.A(net359),
    .B(_00826_),
    .Y(_16025_));
 BUFx2_ASAP7_75t_R input3 (.A(net3456),
    .Y(net3));
 OA211x2_ASAP7_75t_R _21418_ (.A1(net2332),
    .A2(_16024_),
    .B(_16025_),
    .C(net324),
    .Y(_16027_));
 INVx1_ASAP7_75t_R _21419_ (.A(_00827_),
    .Y(_16028_));
 NAND2x1_ASAP7_75t_R _21420_ (.A(net359),
    .B(_00825_),
    .Y(_16029_));
 OA211x2_ASAP7_75t_R _21421_ (.A1(net2332),
    .A2(_16028_),
    .B(_16029_),
    .C(net372),
    .Y(_16030_));
 OR3x1_ASAP7_75t_R _21422_ (.A(net330),
    .B(_16027_),
    .C(_16030_),
    .Y(_16031_));
 BUFx2_ASAP7_75t_R input2 (.A(net3280),
    .Y(net2));
 OA211x2_ASAP7_75t_R _21424_ (.A1(_13373_),
    .A2(_16023_),
    .B(_16031_),
    .C(net334),
    .Y(_16033_));
 INVx1_ASAP7_75t_R _21425_ (.A(_00829_),
    .Y(_16034_));
 BUFx2_ASAP7_75t_R input1 (.A(net3287),
    .Y(net1));
 NOR2x1_ASAP7_75t_R _21427_ (.A(net350),
    .B(_00831_),
    .Y(_16036_));
 AO21x1_ASAP7_75t_R _21428_ (.A1(net350),
    .A2(_16034_),
    .B(_16036_),
    .Y(_16037_));
 INVx1_ASAP7_75t_R _21429_ (.A(_00832_),
    .Y(_16038_));
 NAND2x1_ASAP7_75t_R _21430_ (.A(net350),
    .B(_00830_),
    .Y(_16039_));
 TAPCELL_ASAP7_75t_R TAP_1117 ();
 OA211x2_ASAP7_75t_R _21432_ (.A1(net350),
    .A2(_16038_),
    .B(_16039_),
    .C(net324),
    .Y(_16041_));
 AO21x1_ASAP7_75t_R _21433_ (.A1(net372),
    .A2(_16037_),
    .B(_16041_),
    .Y(_16042_));
 INVx1_ASAP7_75t_R _21434_ (.A(_00824_),
    .Y(_16043_));
 NAND2x1_ASAP7_75t_R _21435_ (.A(net350),
    .B(_00822_),
    .Y(_16044_));
 OA211x2_ASAP7_75t_R _21436_ (.A1(net350),
    .A2(_16043_),
    .B(_16044_),
    .C(net324),
    .Y(_16045_));
 INVx1_ASAP7_75t_R _21437_ (.A(_00823_),
    .Y(_16046_));
 NAND2x1_ASAP7_75t_R _21438_ (.A(net350),
    .B(_00821_),
    .Y(_16047_));
 OA211x2_ASAP7_75t_R _21439_ (.A1(net350),
    .A2(_16046_),
    .B(_16047_),
    .C(net372),
    .Y(_16048_));
 OR3x1_ASAP7_75t_R _21440_ (.A(_13373_),
    .B(_16045_),
    .C(_16048_),
    .Y(_16049_));
 OA211x2_ASAP7_75t_R _21441_ (.A1(net330),
    .A2(_16042_),
    .B(_16049_),
    .C(_13350_),
    .Y(_16050_));
 OR3x1_ASAP7_75t_R _21442_ (.A(_13355_),
    .B(_16033_),
    .C(_16050_),
    .Y(_16051_));
 TAPCELL_ASAP7_75t_R TAP_1116 ();
 INVx1_ASAP7_75t_R _21444_ (.A(_00840_),
    .Y(_16053_));
 TAPCELL_ASAP7_75t_R TAP_1115 ();
 NAND2x1_ASAP7_75t_R _21446_ (.A(net350),
    .B(_00838_),
    .Y(_16055_));
 OA211x2_ASAP7_75t_R _21447_ (.A1(net350),
    .A2(_16053_),
    .B(_16055_),
    .C(net324),
    .Y(_16056_));
 INVx1_ASAP7_75t_R _21448_ (.A(_00839_),
    .Y(_16057_));
 NAND2x1_ASAP7_75t_R _21449_ (.A(net2280),
    .B(_00837_),
    .Y(_16058_));
 OA211x2_ASAP7_75t_R _21450_ (.A1(net2288),
    .A2(_16057_),
    .B(_16058_),
    .C(net371),
    .Y(_16059_));
 OR3x1_ASAP7_75t_R _21451_ (.A(net334),
    .B(_16056_),
    .C(_16059_),
    .Y(_16060_));
 INVx1_ASAP7_75t_R _21452_ (.A(_00836_),
    .Y(_16061_));
 NAND2x1_ASAP7_75t_R _21453_ (.A(net350),
    .B(_00834_),
    .Y(_16062_));
 OA211x2_ASAP7_75t_R _21454_ (.A1(net350),
    .A2(_16061_),
    .B(_16062_),
    .C(net324),
    .Y(_16063_));
 TAPCELL_ASAP7_75t_R TAP_1114 ();
 INVx1_ASAP7_75t_R _21456_ (.A(_00835_),
    .Y(_16065_));
 NAND2x1_ASAP7_75t_R _21457_ (.A(net350),
    .B(_00833_),
    .Y(_16066_));
 OA211x2_ASAP7_75t_R _21458_ (.A1(net350),
    .A2(_16065_),
    .B(_16066_),
    .C(net372),
    .Y(_16067_));
 OR3x1_ASAP7_75t_R _21459_ (.A(_13350_),
    .B(_16063_),
    .C(_16067_),
    .Y(_16068_));
 AND3x1_ASAP7_75t_R _21460_ (.A(net330),
    .B(_16060_),
    .C(_16068_),
    .Y(_16069_));
 INVx1_ASAP7_75t_R _21461_ (.A(_00843_),
    .Y(_16070_));
 NAND2x1_ASAP7_75t_R _21462_ (.A(net2280),
    .B(_00841_),
    .Y(_16071_));
 OA211x2_ASAP7_75t_R _21463_ (.A1(net2288),
    .A2(_16070_),
    .B(_16071_),
    .C(net371),
    .Y(_16072_));
 INVx1_ASAP7_75t_R _21464_ (.A(_00844_),
    .Y(_16073_));
 NAND2x1_ASAP7_75t_R _21465_ (.A(net2280),
    .B(_00842_),
    .Y(_16074_));
 OA211x2_ASAP7_75t_R _21466_ (.A1(net2288),
    .A2(_16073_),
    .B(_16074_),
    .C(net324),
    .Y(_16075_));
 OR3x1_ASAP7_75t_R _21467_ (.A(_13350_),
    .B(_16072_),
    .C(_16075_),
    .Y(_16076_));
 INVx1_ASAP7_75t_R _21468_ (.A(_00848_),
    .Y(_16077_));
 NAND2x1_ASAP7_75t_R _21469_ (.A(net2280),
    .B(_00846_),
    .Y(_16078_));
 OA211x2_ASAP7_75t_R _21470_ (.A1(net2288),
    .A2(_16077_),
    .B(_16078_),
    .C(net324),
    .Y(_16079_));
 TAPCELL_ASAP7_75t_R TAP_1113 ();
 INVx1_ASAP7_75t_R _21472_ (.A(_00847_),
    .Y(_16081_));
 NAND2x1_ASAP7_75t_R _21473_ (.A(net2280),
    .B(_00845_),
    .Y(_16082_));
 OA211x2_ASAP7_75t_R _21474_ (.A1(net2288),
    .A2(_16081_),
    .B(_16082_),
    .C(net371),
    .Y(_16083_));
 OR3x1_ASAP7_75t_R _21475_ (.A(net334),
    .B(_16079_),
    .C(_16083_),
    .Y(_16084_));
 AND3x1_ASAP7_75t_R _21476_ (.A(_13373_),
    .B(_16076_),
    .C(_16084_),
    .Y(_16085_));
 OR3x2_ASAP7_75t_R _21477_ (.A(net327),
    .B(_16069_),
    .C(_16085_),
    .Y(_16086_));
 NAND2x2_ASAP7_75t_R _21478_ (.A(_16051_),
    .B(_16086_),
    .Y(_16087_));
 OA21x2_ASAP7_75t_R _21479_ (.A1(net385),
    .A2(_15490_),
    .B(_15492_),
    .Y(_16088_));
 AOI21x1_ASAP7_75t_R _21480_ (.A1(_13474_),
    .A2(_16087_),
    .B(_16088_),
    .Y(_18410_));
 XOR2x1_ASAP7_75t_R _21481_ (.A(_13620_),
    .Y(_16089_),
    .B(_18410_));
 NOR2x1_ASAP7_75t_R _21482_ (.A(_13986_),
    .B(_16087_),
    .Y(_16090_));
 NAND2x1_ASAP7_75t_R _21483_ (.A(net395),
    .B(_00838_),
    .Y(_16091_));
 OA211x2_ASAP7_75t_R _21484_ (.A1(net395),
    .A2(_16053_),
    .B(_16091_),
    .C(net317),
    .Y(_16092_));
 NAND2x1_ASAP7_75t_R _21485_ (.A(net395),
    .B(_00837_),
    .Y(_16093_));
 OA211x2_ASAP7_75t_R _21486_ (.A1(net395),
    .A2(_16057_),
    .B(_16093_),
    .C(net423),
    .Y(_16094_));
 OR3x1_ASAP7_75t_R _21487_ (.A(net383),
    .B(_16092_),
    .C(_16094_),
    .Y(_16095_));
 NAND2x1_ASAP7_75t_R _21488_ (.A(net395),
    .B(_00834_),
    .Y(_16096_));
 OA211x2_ASAP7_75t_R _21489_ (.A1(net395),
    .A2(_16061_),
    .B(_16096_),
    .C(net317),
    .Y(_16097_));
 NAND2x1_ASAP7_75t_R _21490_ (.A(net395),
    .B(_00833_),
    .Y(_16098_));
 OA211x2_ASAP7_75t_R _21491_ (.A1(net395),
    .A2(_16065_),
    .B(_16098_),
    .C(net423),
    .Y(_16099_));
 OR3x1_ASAP7_75t_R _21492_ (.A(net321),
    .B(_16097_),
    .C(_16099_),
    .Y(_16100_));
 NAND2x1_ASAP7_75t_R _21493_ (.A(net407),
    .B(_00822_),
    .Y(_16101_));
 OA211x2_ASAP7_75t_R _21494_ (.A1(net407),
    .A2(_16043_),
    .B(_16101_),
    .C(net317),
    .Y(_16102_));
 NAND2x1_ASAP7_75t_R _21495_ (.A(net407),
    .B(_00821_),
    .Y(_16103_));
 OA211x2_ASAP7_75t_R _21496_ (.A1(net407),
    .A2(_16046_),
    .B(_16103_),
    .C(net423),
    .Y(_16104_));
 OR3x1_ASAP7_75t_R _21497_ (.A(net312),
    .B(_16102_),
    .C(_16104_),
    .Y(_16105_));
 INVx1_ASAP7_75t_R _21498_ (.A(_00820_),
    .Y(_16106_));
 NAND2x1_ASAP7_75t_R _21499_ (.A(net400),
    .B(_01692_),
    .Y(_16107_));
 OA211x2_ASAP7_75t_R _21500_ (.A1(net400),
    .A2(_16106_),
    .B(_16107_),
    .C(net317),
    .Y(_16108_));
 NOR2x1_ASAP7_75t_R _21501_ (.A(net400),
    .B(_00819_),
    .Y(_16109_));
 AO21x1_ASAP7_75t_R _21502_ (.A1(net423),
    .A2(_16109_),
    .B(_14005_),
    .Y(_16110_));
 OA21x2_ASAP7_75t_R _21503_ (.A1(_16108_),
    .A2(_16110_),
    .B(net377),
    .Y(_16111_));
 AO32x1_ASAP7_75t_R _21504_ (.A1(_13626_),
    .A2(_16095_),
    .A3(_16100_),
    .B1(_16105_),
    .B2(_16111_),
    .Y(_16112_));
 NOR2x1_ASAP7_75t_R _21505_ (.A(net395),
    .B(_00831_),
    .Y(_16113_));
 AO21x1_ASAP7_75t_R _21506_ (.A1(net395),
    .A2(_16034_),
    .B(_16113_),
    .Y(_16114_));
 NAND2x1_ASAP7_75t_R _21507_ (.A(net395),
    .B(_00830_),
    .Y(_16115_));
 OA211x2_ASAP7_75t_R _21508_ (.A1(net395),
    .A2(_16038_),
    .B(_16115_),
    .C(net317),
    .Y(_16116_));
 AO21x1_ASAP7_75t_R _21509_ (.A1(net423),
    .A2(_16114_),
    .B(_16116_),
    .Y(_16117_));
 NAND2x1_ASAP7_75t_R _21510_ (.A(net407),
    .B(_00826_),
    .Y(_16118_));
 OA211x2_ASAP7_75t_R _21511_ (.A1(net407),
    .A2(_16024_),
    .B(_16118_),
    .C(net317),
    .Y(_16119_));
 NAND2x1_ASAP7_75t_R _21512_ (.A(net407),
    .B(_00825_),
    .Y(_16120_));
 OA211x2_ASAP7_75t_R _21513_ (.A1(net407),
    .A2(_16028_),
    .B(_16120_),
    .C(net423),
    .Y(_16121_));
 OA21x2_ASAP7_75t_R _21514_ (.A1(_16119_),
    .A2(_16121_),
    .B(net385),
    .Y(_16122_));
 AO21x1_ASAP7_75t_R _21515_ (.A1(net321),
    .A2(_16117_),
    .B(_16122_),
    .Y(_16123_));
 AND2x2_ASAP7_75t_R _21516_ (.A(_16105_),
    .B(_16111_),
    .Y(_16124_));
 INVx1_ASAP7_75t_R _21517_ (.A(_00841_),
    .Y(_16125_));
 NOR2x1_ASAP7_75t_R _21518_ (.A(net383),
    .B(_00845_),
    .Y(_16126_));
 AO21x1_ASAP7_75t_R _21519_ (.A1(net383),
    .A2(_16125_),
    .B(_16126_),
    .Y(_16127_));
 INVx1_ASAP7_75t_R _21520_ (.A(_00846_),
    .Y(_16128_));
 NAND2x1_ASAP7_75t_R _21521_ (.A(net383),
    .B(_00842_),
    .Y(_16129_));
 OA211x2_ASAP7_75t_R _21522_ (.A1(net383),
    .A2(_16128_),
    .B(_16129_),
    .C(net317),
    .Y(_16130_));
 AO21x1_ASAP7_75t_R _21523_ (.A1(net421),
    .A2(_16127_),
    .B(_16130_),
    .Y(_16131_));
 NAND2x1_ASAP7_75t_R _21524_ (.A(net421),
    .B(_00843_),
    .Y(_16132_));
 OA211x2_ASAP7_75t_R _21525_ (.A1(net421),
    .A2(_16073_),
    .B(_16132_),
    .C(net383),
    .Y(_16133_));
 NAND2x1_ASAP7_75t_R _21526_ (.A(net421),
    .B(_00847_),
    .Y(_16134_));
 OA211x2_ASAP7_75t_R _21527_ (.A1(net421),
    .A2(_16077_),
    .B(_16134_),
    .C(net321),
    .Y(_16135_));
 OR3x1_ASAP7_75t_R _21528_ (.A(net400),
    .B(_16133_),
    .C(_16135_),
    .Y(_16136_));
 OA211x2_ASAP7_75t_R _21529_ (.A1(net316),
    .A2(_16131_),
    .B(_16136_),
    .C(_14780_),
    .Y(_16137_));
 AO221x2_ASAP7_75t_R _21530_ (.A1(net379),
    .A2(_16112_),
    .B1(_16123_),
    .B2(_16124_),
    .C(_16137_),
    .Y(_16138_));
 TAPCELL_ASAP7_75t_R TAP_1112 ();
 AOI22x1_ASAP7_75t_R _21532_ (.A1(_13775_),
    .A2(_00849_),
    .B1(_02216_),
    .B2(_13778_),
    .Y(_16140_));
 OA211x2_ASAP7_75t_R _21533_ (.A1(_00284_),
    .A2(_16138_),
    .B(_16140_),
    .C(_13986_),
    .Y(_16141_));
 OA21x2_ASAP7_75t_R _21534_ (.A1(_16090_),
    .A2(_16141_),
    .B(_13817_),
    .Y(_16142_));
 AOI21x1_ASAP7_75t_R _21535_ (.A1(net308),
    .A2(_16089_),
    .B(_16142_),
    .Y(_17784_));
 INVx1_ASAP7_75t_R _21536_ (.A(_17784_),
    .Y(_16743_));
 INVx2_ASAP7_75t_R _21537_ (.A(_00209_),
    .Y(\cs_registers_i.pc_id_i[17] ));
 INVx1_ASAP7_75t_R _21538_ (.A(_01624_),
    .Y(_16143_));
 AO32x2_ASAP7_75t_R _21539_ (.A1(\cs_registers_i.pc_id_i[17] ),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_16143_),
    .B2(_13450_),
    .Y(_16144_));
 AO21x2_ASAP7_75t_R _21540_ (.A1(_13810_),
    .A2(_16138_),
    .B(_16144_),
    .Y(_16145_));
 TAPCELL_ASAP7_75t_R TAP_1111 ();
 INVx3_ASAP7_75t_R _21542_ (.A(_16145_),
    .Y(_18409_));
 OA21x2_ASAP7_75t_R _21543_ (.A1(_00849_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_16146_));
 AOI21x1_ASAP7_75t_R _21544_ (.A1(net308),
    .A2(_18409_),
    .B(_16146_),
    .Y(_17785_));
 INVx1_ASAP7_75t_R _21545_ (.A(_17785_),
    .Y(_16744_));
 OA21x2_ASAP7_75t_R _21546_ (.A1(_00784_),
    .A2(_15890_),
    .B(_00817_),
    .Y(_16147_));
 OA21x2_ASAP7_75t_R _21547_ (.A1(_02275_),
    .A2(_16147_),
    .B(_02274_),
    .Y(_16745_));
 AND2x2_ASAP7_75t_R _21548_ (.A(net342),
    .B(_01691_),
    .Y(_16148_));
 AO21x1_ASAP7_75t_R _21549_ (.A1(net326),
    .A2(_00852_),
    .B(_16148_),
    .Y(_16149_));
 OAI22x1_ASAP7_75t_R _21550_ (.A1(_00851_),
    .A2(net311),
    .B1(_16149_),
    .B2(net376),
    .Y(_16150_));
 INVx1_ASAP7_75t_R _21551_ (.A(_00860_),
    .Y(_16151_));
 TAPCELL_ASAP7_75t_R TAP_1110 ();
 NAND2x1_ASAP7_75t_R _21553_ (.A(net345),
    .B(_00858_),
    .Y(_16153_));
 TAPCELL_ASAP7_75t_R TAP_1109 ();
 OA211x2_ASAP7_75t_R _21555_ (.A1(net345),
    .A2(_16151_),
    .B(_16153_),
    .C(_13376_),
    .Y(_16155_));
 INVx1_ASAP7_75t_R _21556_ (.A(_00859_),
    .Y(_16156_));
 NAND2x1_ASAP7_75t_R _21557_ (.A(net345),
    .B(_00857_),
    .Y(_16157_));
 OA211x2_ASAP7_75t_R _21558_ (.A1(net345),
    .A2(_16156_),
    .B(_16157_),
    .C(net376),
    .Y(_16158_));
 OR3x1_ASAP7_75t_R _21559_ (.A(net332),
    .B(_16155_),
    .C(_16158_),
    .Y(_16159_));
 OA21x2_ASAP7_75t_R _21560_ (.A1(_13373_),
    .A2(_16150_),
    .B(_16159_),
    .Y(_16160_));
 INVx1_ASAP7_75t_R _21561_ (.A(_00856_),
    .Y(_16161_));
 NAND2x1_ASAP7_75t_R _21562_ (.A(net345),
    .B(_00854_),
    .Y(_16162_));
 OA211x2_ASAP7_75t_R _21563_ (.A1(net345),
    .A2(_16161_),
    .B(_16162_),
    .C(_13376_),
    .Y(_16163_));
 TAPCELL_ASAP7_75t_R TAP_1108 ();
 INVx1_ASAP7_75t_R _21565_ (.A(_00855_),
    .Y(_16165_));
 NAND2x1_ASAP7_75t_R _21566_ (.A(net345),
    .B(_00853_),
    .Y(_16166_));
 OA211x2_ASAP7_75t_R _21567_ (.A1(net345),
    .A2(_16165_),
    .B(_16166_),
    .C(net376),
    .Y(_16167_));
 OR3x1_ASAP7_75t_R _21568_ (.A(_13373_),
    .B(_16163_),
    .C(_16167_),
    .Y(_16168_));
 INVx1_ASAP7_75t_R _21569_ (.A(_00864_),
    .Y(_16169_));
 NAND2x1_ASAP7_75t_R _21570_ (.A(net345),
    .B(_00862_),
    .Y(_16170_));
 OA211x2_ASAP7_75t_R _21571_ (.A1(net345),
    .A2(_16169_),
    .B(_16170_),
    .C(_13376_),
    .Y(_16171_));
 INVx1_ASAP7_75t_R _21572_ (.A(_00863_),
    .Y(_16172_));
 NAND2x1_ASAP7_75t_R _21573_ (.A(net345),
    .B(_00861_),
    .Y(_16173_));
 OA211x2_ASAP7_75t_R _21574_ (.A1(net345),
    .A2(_16172_),
    .B(_16173_),
    .C(net376),
    .Y(_16174_));
 OR3x1_ASAP7_75t_R _21575_ (.A(net332),
    .B(_16171_),
    .C(_16174_),
    .Y(_16175_));
 AND3x1_ASAP7_75t_R _21576_ (.A(_13350_),
    .B(_16168_),
    .C(_16175_),
    .Y(_16176_));
 AO21x1_ASAP7_75t_R _21577_ (.A1(net338),
    .A2(_16160_),
    .B(_16176_),
    .Y(_16177_));
 INVx1_ASAP7_75t_R _21578_ (.A(_00872_),
    .Y(_16178_));
 NAND2x1_ASAP7_75t_R _21579_ (.A(net342),
    .B(_00870_),
    .Y(_16179_));
 OA211x2_ASAP7_75t_R _21580_ (.A1(net342),
    .A2(_16178_),
    .B(_16179_),
    .C(_13376_),
    .Y(_16180_));
 INVx1_ASAP7_75t_R _21581_ (.A(_00871_),
    .Y(_16181_));
 NAND2x1_ASAP7_75t_R _21582_ (.A(net342),
    .B(_00869_),
    .Y(_16182_));
 OA211x2_ASAP7_75t_R _21583_ (.A1(net342),
    .A2(_16181_),
    .B(_16182_),
    .C(net376),
    .Y(_16183_));
 OR3x1_ASAP7_75t_R _21584_ (.A(_13373_),
    .B(_16180_),
    .C(_16183_),
    .Y(_16184_));
 INVx1_ASAP7_75t_R _21585_ (.A(_00880_),
    .Y(_16185_));
 NAND2x1_ASAP7_75t_R _21586_ (.A(net342),
    .B(_00878_),
    .Y(_16186_));
 OA211x2_ASAP7_75t_R _21587_ (.A1(net342),
    .A2(_16185_),
    .B(_16186_),
    .C(_13376_),
    .Y(_16187_));
 INVx1_ASAP7_75t_R _21588_ (.A(_00879_),
    .Y(_16188_));
 NAND2x1_ASAP7_75t_R _21589_ (.A(net342),
    .B(_00877_),
    .Y(_16189_));
 OA211x2_ASAP7_75t_R _21590_ (.A1(net342),
    .A2(_16188_),
    .B(_16189_),
    .C(net376),
    .Y(_16190_));
 OR3x1_ASAP7_75t_R _21591_ (.A(net332),
    .B(_16187_),
    .C(_16190_),
    .Y(_16191_));
 AND3x1_ASAP7_75t_R _21592_ (.A(_13350_),
    .B(_16184_),
    .C(_16191_),
    .Y(_16192_));
 TAPCELL_ASAP7_75t_R TAP_1107 ();
 TAPCELL_ASAP7_75t_R TAP_1106 ();
 INVx1_ASAP7_75t_R _21595_ (.A(_00873_),
    .Y(_16195_));
 TAPCELL_ASAP7_75t_R TAP_1105 ();
 NOR2x1_ASAP7_75t_R _21597_ (.A(net342),
    .B(_00875_),
    .Y(_16197_));
 AO21x1_ASAP7_75t_R _21598_ (.A1(net342),
    .A2(_16195_),
    .B(_16197_),
    .Y(_16198_));
 TAPCELL_ASAP7_75t_R TAP_1104 ();
 INVx1_ASAP7_75t_R _21600_ (.A(_00876_),
    .Y(_16200_));
 NAND2x1_ASAP7_75t_R _21601_ (.A(net342),
    .B(_00874_),
    .Y(_16201_));
 OA211x2_ASAP7_75t_R _21602_ (.A1(net342),
    .A2(_16200_),
    .B(_16201_),
    .C(_13376_),
    .Y(_16202_));
 AO21x1_ASAP7_75t_R _21603_ (.A1(net376),
    .A2(_16198_),
    .B(_16202_),
    .Y(_16203_));
 INVx1_ASAP7_75t_R _21604_ (.A(_00868_),
    .Y(_16204_));
 NAND2x1_ASAP7_75t_R _21605_ (.A(net342),
    .B(_00866_),
    .Y(_16205_));
 OA211x2_ASAP7_75t_R _21606_ (.A1(net342),
    .A2(_16204_),
    .B(_16205_),
    .C(_13376_),
    .Y(_16206_));
 INVx1_ASAP7_75t_R _21607_ (.A(_00867_),
    .Y(_16207_));
 NAND2x1_ASAP7_75t_R _21608_ (.A(net342),
    .B(_00865_),
    .Y(_16208_));
 OA211x2_ASAP7_75t_R _21609_ (.A1(net342),
    .A2(_16207_),
    .B(_16208_),
    .C(net376),
    .Y(_16209_));
 OR3x1_ASAP7_75t_R _21610_ (.A(_13373_),
    .B(_16206_),
    .C(_16209_),
    .Y(_16210_));
 OA211x2_ASAP7_75t_R _21611_ (.A1(net332),
    .A2(_16203_),
    .B(_16210_),
    .C(net338),
    .Y(_16211_));
 OR3x1_ASAP7_75t_R _21612_ (.A(net328),
    .B(_16192_),
    .C(_16211_),
    .Y(_16212_));
 OA21x2_ASAP7_75t_R _21613_ (.A1(_13355_),
    .A2(_16177_),
    .B(_16212_),
    .Y(_16213_));
 OAI21x1_ASAP7_75t_R _21614_ (.A1(net380),
    .A2(_15490_),
    .B(_15492_),
    .Y(_16214_));
 OA21x2_ASAP7_75t_R _21615_ (.A1(_13521_),
    .A2(_16213_),
    .B(_16214_),
    .Y(_18415_));
 AND2x2_ASAP7_75t_R _21616_ (.A(net389),
    .B(_01691_),
    .Y(_16215_));
 AO21x1_ASAP7_75t_R _21617_ (.A1(_13675_),
    .A2(_00852_),
    .B(_16215_),
    .Y(_16216_));
 OAI22x1_ASAP7_75t_R _21618_ (.A1(_00851_),
    .A2(net2290),
    .B1(_16216_),
    .B2(net427),
    .Y(_16217_));
 TAPCELL_ASAP7_75t_R TAP_1103 ();
 NAND2x1_ASAP7_75t_R _21620_ (.A(net391),
    .B(_00858_),
    .Y(_16219_));
 OA211x2_ASAP7_75t_R _21621_ (.A1(net391),
    .A2(_16151_),
    .B(_16219_),
    .C(_13649_),
    .Y(_16220_));
 NAND2x1_ASAP7_75t_R _21622_ (.A(net391),
    .B(_00857_),
    .Y(_16221_));
 OA211x2_ASAP7_75t_R _21623_ (.A1(net391),
    .A2(_16156_),
    .B(_16221_),
    .C(net427),
    .Y(_16222_));
 OR3x1_ASAP7_75t_R _21624_ (.A(net381),
    .B(_16220_),
    .C(_16222_),
    .Y(_16223_));
 OA211x2_ASAP7_75t_R _21625_ (.A1(_13636_),
    .A2(_16217_),
    .B(_16223_),
    .C(net387),
    .Y(_16224_));
 TAPCELL_ASAP7_75t_R TAP_1102 ();
 NAND2x1_ASAP7_75t_R _21627_ (.A(net391),
    .B(_00853_),
    .Y(_16226_));
 OA211x2_ASAP7_75t_R _21628_ (.A1(net391),
    .A2(_16165_),
    .B(_16226_),
    .C(net381),
    .Y(_16227_));
 NAND2x1_ASAP7_75t_R _21629_ (.A(net391),
    .B(_00861_),
    .Y(_16228_));
 OA211x2_ASAP7_75t_R _21630_ (.A1(net391),
    .A2(_16172_),
    .B(_16228_),
    .C(_13636_),
    .Y(_16229_));
 OR3x1_ASAP7_75t_R _21631_ (.A(_13649_),
    .B(_16227_),
    .C(_16229_),
    .Y(_16230_));
 NAND2x1_ASAP7_75t_R _21632_ (.A(net391),
    .B(_00854_),
    .Y(_16231_));
 OA211x2_ASAP7_75t_R _21633_ (.A1(net391),
    .A2(_16161_),
    .B(_16231_),
    .C(net381),
    .Y(_16232_));
 NAND2x1_ASAP7_75t_R _21634_ (.A(net391),
    .B(_00862_),
    .Y(_16233_));
 OA211x2_ASAP7_75t_R _21635_ (.A1(net391),
    .A2(_16169_),
    .B(_16233_),
    .C(_13636_),
    .Y(_16234_));
 OR3x1_ASAP7_75t_R _21636_ (.A(net427),
    .B(_16232_),
    .C(_16234_),
    .Y(_16235_));
 AND3x1_ASAP7_75t_R _21637_ (.A(_13630_),
    .B(_16230_),
    .C(_16235_),
    .Y(_16236_));
 OR3x2_ASAP7_75t_R _21638_ (.A(_13626_),
    .B(_16224_),
    .C(_16236_),
    .Y(_16237_));
 NAND2x1_ASAP7_75t_R _21639_ (.A(net393),
    .B(_00870_),
    .Y(_16238_));
 OA211x2_ASAP7_75t_R _21640_ (.A1(net393),
    .A2(_16178_),
    .B(_16238_),
    .C(_13649_),
    .Y(_16239_));
 NAND2x1_ASAP7_75t_R _21641_ (.A(net389),
    .B(_00869_),
    .Y(_16240_));
 OA211x2_ASAP7_75t_R _21642_ (.A1(net389),
    .A2(_16181_),
    .B(_16240_),
    .C(net427),
    .Y(_16241_));
 OR3x1_ASAP7_75t_R _21643_ (.A(net387),
    .B(_16239_),
    .C(_16241_),
    .Y(_16242_));
 NAND2x1_ASAP7_75t_R _21644_ (.A(net389),
    .B(_00866_),
    .Y(_16243_));
 OA211x2_ASAP7_75t_R _21645_ (.A1(net389),
    .A2(_16204_),
    .B(_16243_),
    .C(_13649_),
    .Y(_16244_));
 NAND2x1_ASAP7_75t_R _21646_ (.A(net389),
    .B(_00865_),
    .Y(_16245_));
 OA211x2_ASAP7_75t_R _21647_ (.A1(net389),
    .A2(_16207_),
    .B(_16245_),
    .C(net427),
    .Y(_16246_));
 OR3x1_ASAP7_75t_R _21648_ (.A(_13630_),
    .B(_16244_),
    .C(_16246_),
    .Y(_16247_));
 AND3x1_ASAP7_75t_R _21649_ (.A(net382),
    .B(_16242_),
    .C(_16247_),
    .Y(_16248_));
 NOR2x1_ASAP7_75t_R _21650_ (.A(net391),
    .B(_00875_),
    .Y(_16249_));
 AO21x1_ASAP7_75t_R _21651_ (.A1(net391),
    .A2(_16195_),
    .B(_16249_),
    .Y(_16250_));
 NAND2x1_ASAP7_75t_R _21652_ (.A(net389),
    .B(_00874_),
    .Y(_16251_));
 OA211x2_ASAP7_75t_R _21653_ (.A1(net389),
    .A2(_16200_),
    .B(_16251_),
    .C(_13649_),
    .Y(_16252_));
 AO21x1_ASAP7_75t_R _21654_ (.A1(net427),
    .A2(_16250_),
    .B(_16252_),
    .Y(_16253_));
 NAND2x1_ASAP7_75t_R _21655_ (.A(net389),
    .B(_00878_),
    .Y(_16254_));
 OA211x2_ASAP7_75t_R _21656_ (.A1(net389),
    .A2(_16185_),
    .B(_16254_),
    .C(_13649_),
    .Y(_16255_));
 NAND2x1_ASAP7_75t_R _21657_ (.A(net391),
    .B(_00877_),
    .Y(_16256_));
 OA211x2_ASAP7_75t_R _21658_ (.A1(net391),
    .A2(_16188_),
    .B(_16256_),
    .C(net427),
    .Y(_16257_));
 OR3x1_ASAP7_75t_R _21659_ (.A(net387),
    .B(_16255_),
    .C(_16257_),
    .Y(_16258_));
 OA211x2_ASAP7_75t_R _21660_ (.A1(_13630_),
    .A2(_16253_),
    .B(_16258_),
    .C(_13636_),
    .Y(_16259_));
 OR3x1_ASAP7_75t_R _21661_ (.A(_00286_),
    .B(_16248_),
    .C(_16259_),
    .Y(_16260_));
 NAND2x2_ASAP7_75t_R _21662_ (.A(_16237_),
    .B(_16260_),
    .Y(_16261_));
 OA222x2_ASAP7_75t_R _21663_ (.A1(_01623_),
    .A2(_13807_),
    .B1(_15112_),
    .B2(_16261_),
    .C1(_14103_),
    .C2(_00211_),
    .Y(_16262_));
 TAPCELL_ASAP7_75t_R TAP_1101 ();
 XOR2x2_ASAP7_75t_R _21665_ (.A(_00882_),
    .B(_02228_),
    .Y(_16263_));
 INVx4_ASAP7_75t_R _21666_ (.A(_16263_),
    .Y(net159));
 TAPCELL_ASAP7_75t_R TAP_1100 ();
 INVx1_ASAP7_75t_R _21668_ (.A(_00905_),
    .Y(_16265_));
 NAND2x1_ASAP7_75t_R _21669_ (.A(net2343),
    .B(_00903_),
    .Y(_16266_));
 OA21x2_ASAP7_75t_R _21670_ (.A1(net2331),
    .A2(_16265_),
    .B(_16266_),
    .Y(_16267_));
 INVx1_ASAP7_75t_R _21671_ (.A(_00904_),
    .Y(_16268_));
 NAND2x1_ASAP7_75t_R _21672_ (.A(net2343),
    .B(_00902_),
    .Y(_16269_));
 OA211x2_ASAP7_75t_R _21673_ (.A1(net2331),
    .A2(_16268_),
    .B(_16269_),
    .C(net371),
    .Y(_16270_));
 AO21x1_ASAP7_75t_R _21674_ (.A1(net324),
    .A2(_16267_),
    .B(_16270_),
    .Y(_16271_));
 INVx1_ASAP7_75t_R _21675_ (.A(_00901_),
    .Y(_16272_));
 NAND2x1_ASAP7_75t_R _21676_ (.A(net2343),
    .B(_00899_),
    .Y(_16273_));
 OA211x2_ASAP7_75t_R _21677_ (.A1(net2331),
    .A2(_16272_),
    .B(_16273_),
    .C(net324),
    .Y(_16274_));
 INVx1_ASAP7_75t_R _21678_ (.A(_00900_),
    .Y(_16275_));
 NAND2x1_ASAP7_75t_R _21679_ (.A(net2343),
    .B(_00898_),
    .Y(_16276_));
 OA211x2_ASAP7_75t_R _21680_ (.A1(net2331),
    .A2(_16275_),
    .B(_16276_),
    .C(net371),
    .Y(_16277_));
 OR3x1_ASAP7_75t_R _21681_ (.A(_13350_),
    .B(_16274_),
    .C(_16277_),
    .Y(_16278_));
 OA21x2_ASAP7_75t_R _21682_ (.A1(net334),
    .A2(_16271_),
    .B(_16278_),
    .Y(_16279_));
 INVx1_ASAP7_75t_R _21683_ (.A(_00908_),
    .Y(_16280_));
 NAND2x1_ASAP7_75t_R _21684_ (.A(net2294),
    .B(_00906_),
    .Y(_16281_));
 OA211x2_ASAP7_75t_R _21685_ (.A1(net2321),
    .A2(_16280_),
    .B(_16281_),
    .C(net371),
    .Y(_16282_));
 INVx1_ASAP7_75t_R _21686_ (.A(_00909_),
    .Y(_16283_));
 NAND2x1_ASAP7_75t_R _21687_ (.A(net2321),
    .B(_00907_),
    .Y(_16284_));
 OA211x2_ASAP7_75t_R _21688_ (.A1(net2321),
    .A2(_16283_),
    .B(_16284_),
    .C(net324),
    .Y(_16285_));
 OR3x1_ASAP7_75t_R _21689_ (.A(_13350_),
    .B(_16282_),
    .C(_16285_),
    .Y(_16286_));
 INVx1_ASAP7_75t_R _21690_ (.A(_00913_),
    .Y(_16287_));
 NAND2x1_ASAP7_75t_R _21691_ (.A(net2321),
    .B(_00911_),
    .Y(_16288_));
 OA211x2_ASAP7_75t_R _21692_ (.A1(net2321),
    .A2(_16287_),
    .B(_16288_),
    .C(net324),
    .Y(_16289_));
 INVx1_ASAP7_75t_R _21693_ (.A(_00912_),
    .Y(_16290_));
 NAND2x1_ASAP7_75t_R _21694_ (.A(net2294),
    .B(_00910_),
    .Y(_16291_));
 OA211x2_ASAP7_75t_R _21695_ (.A1(net2321),
    .A2(_16290_),
    .B(_16291_),
    .C(net371),
    .Y(_16292_));
 OR3x1_ASAP7_75t_R _21696_ (.A(net334),
    .B(_16289_),
    .C(_16292_),
    .Y(_16293_));
 AND3x1_ASAP7_75t_R _21697_ (.A(_13373_),
    .B(_16286_),
    .C(_16293_),
    .Y(_16294_));
 AO21x1_ASAP7_75t_R _21698_ (.A1(net330),
    .A2(_16279_),
    .B(_16294_),
    .Y(_16295_));
 AND2x2_ASAP7_75t_R _21699_ (.A(net2288),
    .B(_01690_),
    .Y(_16296_));
 AO21x1_ASAP7_75t_R _21700_ (.A1(_13359_),
    .A2(_00885_),
    .B(_16296_),
    .Y(_16297_));
 OAI22x1_ASAP7_75t_R _21701_ (.A1(_00884_),
    .A2(_14184_),
    .B1(_16297_),
    .B2(net371),
    .Y(_16298_));
 INVx1_ASAP7_75t_R _21702_ (.A(_00893_),
    .Y(_16299_));
 NAND2x1_ASAP7_75t_R _21703_ (.A(net2342),
    .B(_00891_),
    .Y(_16300_));
 OA211x2_ASAP7_75t_R _21704_ (.A1(net2331),
    .A2(_16299_),
    .B(_16300_),
    .C(net324),
    .Y(_16301_));
 INVx1_ASAP7_75t_R _21705_ (.A(_00892_),
    .Y(_16302_));
 NAND2x1_ASAP7_75t_R _21706_ (.A(net2342),
    .B(_00890_),
    .Y(_16303_));
 OA211x2_ASAP7_75t_R _21707_ (.A1(net2331),
    .A2(_16302_),
    .B(_16303_),
    .C(net371),
    .Y(_16304_));
 OR3x1_ASAP7_75t_R _21708_ (.A(net330),
    .B(_16301_),
    .C(_16304_),
    .Y(_16305_));
 OA211x2_ASAP7_75t_R _21709_ (.A1(_13373_),
    .A2(_16298_),
    .B(_16305_),
    .C(net334),
    .Y(_16306_));
 INVx1_ASAP7_75t_R _21710_ (.A(_00894_),
    .Y(_16307_));
 NOR2x1_ASAP7_75t_R _21711_ (.A(net2344),
    .B(_00896_),
    .Y(_16308_));
 AO21x1_ASAP7_75t_R _21712_ (.A1(net2331),
    .A2(_16307_),
    .B(_16308_),
    .Y(_16309_));
 TAPCELL_ASAP7_75t_R TAP_1099 ();
 INVx1_ASAP7_75t_R _21714_ (.A(_00897_),
    .Y(_16311_));
 NAND2x1_ASAP7_75t_R _21715_ (.A(net2288),
    .B(_00895_),
    .Y(_16312_));
 OA211x2_ASAP7_75t_R _21716_ (.A1(net2288),
    .A2(_16311_),
    .B(_16312_),
    .C(net324),
    .Y(_16313_));
 AO21x1_ASAP7_75t_R _21717_ (.A1(net371),
    .A2(_16309_),
    .B(_16313_),
    .Y(_16314_));
 INVx1_ASAP7_75t_R _21718_ (.A(_00889_),
    .Y(_16315_));
 NAND2x1_ASAP7_75t_R _21719_ (.A(net2342),
    .B(_00887_),
    .Y(_16316_));
 OA211x2_ASAP7_75t_R _21720_ (.A1(net2331),
    .A2(_16315_),
    .B(_16316_),
    .C(net324),
    .Y(_16317_));
 INVx1_ASAP7_75t_R _21721_ (.A(_00888_),
    .Y(_16318_));
 NAND2x1_ASAP7_75t_R _21722_ (.A(net2342),
    .B(_00886_),
    .Y(_16319_));
 OA211x2_ASAP7_75t_R _21723_ (.A1(net2331),
    .A2(_16318_),
    .B(_16319_),
    .C(net371),
    .Y(_16320_));
 OR3x1_ASAP7_75t_R _21724_ (.A(_13373_),
    .B(_16317_),
    .C(_16320_),
    .Y(_16321_));
 OA211x2_ASAP7_75t_R _21725_ (.A1(net330),
    .A2(_16314_),
    .B(_16321_),
    .C(_13350_),
    .Y(_16322_));
 OA21x2_ASAP7_75t_R _21726_ (.A1(_16306_),
    .A2(_16322_),
    .B(net327),
    .Y(_16323_));
 AO21x2_ASAP7_75t_R _21727_ (.A1(_13355_),
    .A2(_16295_),
    .B(_16323_),
    .Y(_16324_));
 TAPCELL_ASAP7_75t_R TAP_1098 ();
 OAI21x1_ASAP7_75t_R _21729_ (.A1(net377),
    .A2(_15490_),
    .B(_15492_),
    .Y(_16326_));
 OA21x2_ASAP7_75t_R _21730_ (.A1(_13521_),
    .A2(_16324_),
    .B(_16326_),
    .Y(_18419_));
 TAPCELL_ASAP7_75t_R TAP_1097 ();
 XOR2x1_ASAP7_75t_R _21732_ (.A(_13620_),
    .Y(_16328_),
    .B(_18419_));
 INVx1_ASAP7_75t_R _21733_ (.A(_16324_),
    .Y(_16329_));
 NAND2x1_ASAP7_75t_R _21734_ (.A(net394),
    .B(_00902_),
    .Y(_16330_));
 OA211x2_ASAP7_75t_R _21735_ (.A1(net394),
    .A2(_16268_),
    .B(_16330_),
    .C(net321),
    .Y(_16331_));
 TAPCELL_ASAP7_75t_R TAP_1096 ();
 NAND2x1_ASAP7_75t_R _21737_ (.A(net394),
    .B(_00898_),
    .Y(_16333_));
 OA211x2_ASAP7_75t_R _21738_ (.A1(net394),
    .A2(_16275_),
    .B(_16333_),
    .C(net383),
    .Y(_16334_));
 OR3x1_ASAP7_75t_R _21739_ (.A(net317),
    .B(_16331_),
    .C(_16334_),
    .Y(_16335_));
 NAND2x1_ASAP7_75t_R _21740_ (.A(net394),
    .B(_00903_),
    .Y(_16336_));
 OA211x2_ASAP7_75t_R _21741_ (.A1(net394),
    .A2(_16265_),
    .B(_16336_),
    .C(net321),
    .Y(_16337_));
 NAND2x1_ASAP7_75t_R _21742_ (.A(net394),
    .B(_00899_),
    .Y(_16338_));
 OA211x2_ASAP7_75t_R _21743_ (.A1(net394),
    .A2(_16272_),
    .B(_16338_),
    .C(net383),
    .Y(_16339_));
 OR3x1_ASAP7_75t_R _21744_ (.A(net421),
    .B(_16337_),
    .C(_16339_),
    .Y(_16340_));
 NAND2x1_ASAP7_75t_R _21745_ (.A(net399),
    .B(_00886_),
    .Y(_16341_));
 OA211x2_ASAP7_75t_R _21746_ (.A1(net399),
    .A2(_16318_),
    .B(_16341_),
    .C(net421),
    .Y(_16342_));
 NAND2x1_ASAP7_75t_R _21747_ (.A(net399),
    .B(_00887_),
    .Y(_16343_));
 OA211x2_ASAP7_75t_R _21748_ (.A1(net399),
    .A2(_16315_),
    .B(_16343_),
    .C(net317),
    .Y(_16344_));
 OR3x1_ASAP7_75t_R _21749_ (.A(net312),
    .B(_16342_),
    .C(_16344_),
    .Y(_16345_));
 INVx1_ASAP7_75t_R _21750_ (.A(_00885_),
    .Y(_16346_));
 NAND2x1_ASAP7_75t_R _21751_ (.A(net399),
    .B(_01690_),
    .Y(_16347_));
 OA211x2_ASAP7_75t_R _21752_ (.A1(net399),
    .A2(_16346_),
    .B(_16347_),
    .C(net317),
    .Y(_16348_));
 NOR2x1_ASAP7_75t_R _21753_ (.A(net399),
    .B(_00884_),
    .Y(_16349_));
 AO21x1_ASAP7_75t_R _21754_ (.A1(net421),
    .A2(_16349_),
    .B(_14005_),
    .Y(_16350_));
 OA21x2_ASAP7_75t_R _21755_ (.A1(_16348_),
    .A2(_16350_),
    .B(net377),
    .Y(_16351_));
 AO32x1_ASAP7_75t_R _21756_ (.A1(_13626_),
    .A2(_16335_),
    .A3(_16340_),
    .B1(_16345_),
    .B2(_16351_),
    .Y(_16352_));
 NOR2x1_ASAP7_75t_R _21757_ (.A(net395),
    .B(_00896_),
    .Y(_16353_));
 AO21x1_ASAP7_75t_R _21758_ (.A1(net395),
    .A2(_16307_),
    .B(_16353_),
    .Y(_16354_));
 NAND2x1_ASAP7_75t_R _21759_ (.A(net395),
    .B(_00895_),
    .Y(_16355_));
 OA211x2_ASAP7_75t_R _21760_ (.A1(net395),
    .A2(_16311_),
    .B(_16355_),
    .C(net317),
    .Y(_16356_));
 AO21x1_ASAP7_75t_R _21761_ (.A1(net421),
    .A2(_16354_),
    .B(_16356_),
    .Y(_16357_));
 NAND2x1_ASAP7_75t_R _21762_ (.A(net399),
    .B(_00891_),
    .Y(_16358_));
 OA211x2_ASAP7_75t_R _21763_ (.A1(net399),
    .A2(_16299_),
    .B(_16358_),
    .C(net317),
    .Y(_16359_));
 NAND2x1_ASAP7_75t_R _21764_ (.A(net399),
    .B(_00890_),
    .Y(_16360_));
 OA211x2_ASAP7_75t_R _21765_ (.A1(net399),
    .A2(_16302_),
    .B(_16360_),
    .C(net421),
    .Y(_16361_));
 OA21x2_ASAP7_75t_R _21766_ (.A1(_16359_),
    .A2(_16361_),
    .B(net383),
    .Y(_16362_));
 AO21x1_ASAP7_75t_R _21767_ (.A1(net321),
    .A2(_16357_),
    .B(_16362_),
    .Y(_16363_));
 AND2x2_ASAP7_75t_R _21768_ (.A(_16345_),
    .B(_16351_),
    .Y(_16364_));
 TAPCELL_ASAP7_75t_R TAP_1095 ();
 INVx1_ASAP7_75t_R _21770_ (.A(_00906_),
    .Y(_16366_));
 NOR2x1_ASAP7_75t_R _21771_ (.A(net383),
    .B(_00910_),
    .Y(_16367_));
 AO21x1_ASAP7_75t_R _21772_ (.A1(net383),
    .A2(_16366_),
    .B(_16367_),
    .Y(_16368_));
 NAND2x1_ASAP7_75t_R _21773_ (.A(net383),
    .B(_00908_),
    .Y(_16369_));
 OA211x2_ASAP7_75t_R _21774_ (.A1(net383),
    .A2(_16290_),
    .B(_16369_),
    .C(net316),
    .Y(_16370_));
 AO21x1_ASAP7_75t_R _21775_ (.A1(net394),
    .A2(_16368_),
    .B(_16370_),
    .Y(_16371_));
 NAND2x1_ASAP7_75t_R _21776_ (.A(net394),
    .B(_00911_),
    .Y(_16372_));
 OA211x2_ASAP7_75t_R _21777_ (.A1(net394),
    .A2(_16287_),
    .B(_16372_),
    .C(net321),
    .Y(_16373_));
 NAND2x1_ASAP7_75t_R _21778_ (.A(net394),
    .B(_00907_),
    .Y(_16374_));
 OA211x2_ASAP7_75t_R _21779_ (.A1(net394),
    .A2(_16283_),
    .B(_16374_),
    .C(net383),
    .Y(_16375_));
 OR3x1_ASAP7_75t_R _21780_ (.A(net421),
    .B(_16373_),
    .C(_16375_),
    .Y(_16376_));
 OA211x2_ASAP7_75t_R _21781_ (.A1(net317),
    .A2(_16371_),
    .B(_16376_),
    .C(_14780_),
    .Y(_16377_));
 AO221x2_ASAP7_75t_R _21782_ (.A1(net379),
    .A2(_16352_),
    .B1(_16363_),
    .B2(_16364_),
    .C(_16377_),
    .Y(_16378_));
 NOR2x1_ASAP7_75t_R _21783_ (.A(_00284_),
    .B(_16378_),
    .Y(_16379_));
 TAPCELL_ASAP7_75t_R TAP_1094 ();
 AO221x1_ASAP7_75t_R _21785_ (.A1(_13775_),
    .A2(_00914_),
    .B1(_02214_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_16381_));
 OA22x2_ASAP7_75t_R _21786_ (.A1(_13986_),
    .A2(_16329_),
    .B1(_16379_),
    .B2(_16381_),
    .Y(_16382_));
 NOR2x1_ASAP7_75t_R _21787_ (.A(net308),
    .B(_16382_),
    .Y(_16383_));
 AOI21x1_ASAP7_75t_R _21788_ (.A1(net308),
    .A2(_16328_),
    .B(_16383_),
    .Y(_17788_));
 INVx1_ASAP7_75t_R _21789_ (.A(_17788_),
    .Y(_16746_));
 INVx2_ASAP7_75t_R _21790_ (.A(_00212_),
    .Y(\cs_registers_i.pc_id_i[19] ));
 INVx1_ASAP7_75t_R _21791_ (.A(_01622_),
    .Y(_16384_));
 AND3x1_ASAP7_75t_R _21792_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_13993_),
    .C(_13794_),
    .Y(_16385_));
 AOI221x1_ASAP7_75t_R _21793_ (.A1(_16384_),
    .A2(_13450_),
    .B1(_13810_),
    .B2(_16378_),
    .C(_16385_),
    .Y(_16386_));
 TAPCELL_ASAP7_75t_R TAP_1093 ();
 OA21x2_ASAP7_75t_R _21795_ (.A1(_00914_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_16387_));
 AOI21x1_ASAP7_75t_R _21796_ (.A1(net308),
    .A2(_16386_),
    .B(_16387_),
    .Y(_17789_));
 INVx1_ASAP7_75t_R _21797_ (.A(_17789_),
    .Y(_16748_));
 OR5x2_ASAP7_75t_R _21798_ (.A(_00751_),
    .B(_00784_),
    .C(_00882_),
    .D(_00850_),
    .E(_02275_),
    .Y(_16388_));
 OA21x2_ASAP7_75t_R _21799_ (.A1(_00817_),
    .A2(_02275_),
    .B(_02274_),
    .Y(_16389_));
 OA21x2_ASAP7_75t_R _21800_ (.A1(_00850_),
    .A2(_16389_),
    .B(_00883_),
    .Y(_16390_));
 OR5x1_ASAP7_75t_R _21801_ (.A(_00784_),
    .B(_00882_),
    .C(_00850_),
    .D(_02275_),
    .E(_15889_),
    .Y(_16391_));
 OA211x2_ASAP7_75t_R _21802_ (.A1(_00882_),
    .A2(_16390_),
    .B(_16391_),
    .C(_02276_),
    .Y(_16392_));
 OA21x2_ASAP7_75t_R _21803_ (.A1(_15888_),
    .A2(_16388_),
    .B(_16392_),
    .Y(_16747_));
 INVx1_ASAP7_75t_R _21804_ (.A(_00916_),
    .Y(_16393_));
 INVx1_ASAP7_75t_R _21805_ (.A(_00917_),
    .Y(_16394_));
 NAND2x1_ASAP7_75t_R _21806_ (.A(net340),
    .B(_01689_),
    .Y(_16395_));
 OA211x2_ASAP7_75t_R _21807_ (.A1(net340),
    .A2(_16394_),
    .B(_16395_),
    .C(_13376_),
    .Y(_16396_));
 AO21x1_ASAP7_75t_R _21808_ (.A1(_16393_),
    .A2(net2216),
    .B(_16396_),
    .Y(_16397_));
 INVx1_ASAP7_75t_R _21809_ (.A(_00925_),
    .Y(_16398_));
 NAND2x1_ASAP7_75t_R _21810_ (.A(net343),
    .B(_00923_),
    .Y(_16399_));
 OA211x2_ASAP7_75t_R _21811_ (.A1(net343),
    .A2(_16398_),
    .B(_16399_),
    .C(_13376_),
    .Y(_16400_));
 INVx1_ASAP7_75t_R _21812_ (.A(_00924_),
    .Y(_16401_));
 NAND2x1_ASAP7_75t_R _21813_ (.A(net345),
    .B(_00922_),
    .Y(_16402_));
 OA211x2_ASAP7_75t_R _21814_ (.A1(net345),
    .A2(_16401_),
    .B(_16402_),
    .C(net376),
    .Y(_16403_));
 OR3x1_ASAP7_75t_R _21815_ (.A(net332),
    .B(_16400_),
    .C(_16403_),
    .Y(_16404_));
 OA21x2_ASAP7_75t_R _21816_ (.A1(_13373_),
    .A2(_16397_),
    .B(_16404_),
    .Y(_16405_));
 TAPCELL_ASAP7_75t_R TAP_1092 ();
 INVx1_ASAP7_75t_R _21818_ (.A(_00921_),
    .Y(_16407_));
 NAND2x1_ASAP7_75t_R _21819_ (.A(net343),
    .B(_00919_),
    .Y(_16408_));
 OA211x2_ASAP7_75t_R _21820_ (.A1(net343),
    .A2(_16407_),
    .B(_16408_),
    .C(_13376_),
    .Y(_16409_));
 INVx1_ASAP7_75t_R _21821_ (.A(_00920_),
    .Y(_16410_));
 NAND2x1_ASAP7_75t_R _21822_ (.A(net343),
    .B(_00918_),
    .Y(_16411_));
 TAPCELL_ASAP7_75t_R TAP_1091 ();
 OA211x2_ASAP7_75t_R _21824_ (.A1(net343),
    .A2(_16410_),
    .B(_16411_),
    .C(net2314),
    .Y(_16413_));
 OR3x1_ASAP7_75t_R _21825_ (.A(_13373_),
    .B(_16409_),
    .C(_16413_),
    .Y(_16414_));
 INVx1_ASAP7_75t_R _21826_ (.A(_00929_),
    .Y(_16415_));
 NAND2x1_ASAP7_75t_R _21827_ (.A(net344),
    .B(_00927_),
    .Y(_16416_));
 OA211x2_ASAP7_75t_R _21828_ (.A1(net344),
    .A2(_16415_),
    .B(_16416_),
    .C(_13376_),
    .Y(_16417_));
 INVx1_ASAP7_75t_R _21829_ (.A(_00928_),
    .Y(_16418_));
 NAND2x1_ASAP7_75t_R _21830_ (.A(net344),
    .B(_00926_),
    .Y(_16419_));
 OA211x2_ASAP7_75t_R _21831_ (.A1(net344),
    .A2(_16418_),
    .B(_16419_),
    .C(net2315),
    .Y(_16420_));
 OR3x1_ASAP7_75t_R _21832_ (.A(_00245_),
    .B(_16417_),
    .C(_16420_),
    .Y(_16421_));
 AND3x1_ASAP7_75t_R _21833_ (.A(_13350_),
    .B(_16414_),
    .C(_16421_),
    .Y(_16422_));
 AO21x1_ASAP7_75t_R _21834_ (.A1(net338),
    .A2(_16405_),
    .B(_16422_),
    .Y(_16423_));
 INVx1_ASAP7_75t_R _21835_ (.A(_00945_),
    .Y(_16424_));
 NAND2x1_ASAP7_75t_R _21836_ (.A(net343),
    .B(_00943_),
    .Y(_16425_));
 OA211x2_ASAP7_75t_R _21837_ (.A1(net343),
    .A2(_16424_),
    .B(_16425_),
    .C(_13376_),
    .Y(_16426_));
 INVx1_ASAP7_75t_R _21838_ (.A(_00944_),
    .Y(_16427_));
 NAND2x1_ASAP7_75t_R _21839_ (.A(net343),
    .B(_00942_),
    .Y(_16428_));
 OA211x2_ASAP7_75t_R _21840_ (.A1(net343),
    .A2(_16427_),
    .B(_16428_),
    .C(net2314),
    .Y(_16429_));
 OR3x1_ASAP7_75t_R _21841_ (.A(net338),
    .B(_16426_),
    .C(_16429_),
    .Y(_16430_));
 INVx1_ASAP7_75t_R _21842_ (.A(_00941_),
    .Y(_16431_));
 NAND2x1_ASAP7_75t_R _21843_ (.A(net343),
    .B(_00939_),
    .Y(_16432_));
 OA211x2_ASAP7_75t_R _21844_ (.A1(net343),
    .A2(_16431_),
    .B(_16432_),
    .C(_13376_),
    .Y(_16433_));
 INVx1_ASAP7_75t_R _21845_ (.A(_00940_),
    .Y(_16434_));
 NAND2x1_ASAP7_75t_R _21846_ (.A(net343),
    .B(_00938_),
    .Y(_16435_));
 OA211x2_ASAP7_75t_R _21847_ (.A1(net343),
    .A2(_16434_),
    .B(_16435_),
    .C(net2314),
    .Y(_16436_));
 OR3x1_ASAP7_75t_R _21848_ (.A(_13350_),
    .B(_16433_),
    .C(_16436_),
    .Y(_16437_));
 AND3x1_ASAP7_75t_R _21849_ (.A(_13373_),
    .B(_16430_),
    .C(_16437_),
    .Y(_16438_));
 INVx1_ASAP7_75t_R _21850_ (.A(_00930_),
    .Y(_16439_));
 NOR2x1_ASAP7_75t_R _21851_ (.A(net340),
    .B(_00932_),
    .Y(_16440_));
 AO21x1_ASAP7_75t_R _21852_ (.A1(net340),
    .A2(_16439_),
    .B(_16440_),
    .Y(_16441_));
 INVx1_ASAP7_75t_R _21853_ (.A(_00933_),
    .Y(_16442_));
 TAPCELL_ASAP7_75t_R TAP_1090 ();
 NAND2x1_ASAP7_75t_R _21855_ (.A(net340),
    .B(_00931_),
    .Y(_16444_));
 OA211x2_ASAP7_75t_R _21856_ (.A1(net340),
    .A2(_16442_),
    .B(_16444_),
    .C(_13376_),
    .Y(_16445_));
 AO21x1_ASAP7_75t_R _21857_ (.A1(net370),
    .A2(_16441_),
    .B(_16445_),
    .Y(_16446_));
 INVx1_ASAP7_75t_R _21858_ (.A(_00937_),
    .Y(_16447_));
 NAND2x1_ASAP7_75t_R _21859_ (.A(net340),
    .B(_00935_),
    .Y(_16448_));
 OA211x2_ASAP7_75t_R _21860_ (.A1(net340),
    .A2(_16447_),
    .B(_16448_),
    .C(_13376_),
    .Y(_16449_));
 INVx1_ASAP7_75t_R _21861_ (.A(_00936_),
    .Y(_16450_));
 NAND2x1_ASAP7_75t_R _21862_ (.A(net340),
    .B(_00934_),
    .Y(_16451_));
 OA211x2_ASAP7_75t_R _21863_ (.A1(net340),
    .A2(_16450_),
    .B(_16451_),
    .C(net370),
    .Y(_16452_));
 OR3x1_ASAP7_75t_R _21864_ (.A(net337),
    .B(_16449_),
    .C(_16452_),
    .Y(_16453_));
 OA211x2_ASAP7_75t_R _21865_ (.A1(_13350_),
    .A2(_16446_),
    .B(_16453_),
    .C(net332),
    .Y(_16454_));
 OR3x1_ASAP7_75t_R _21866_ (.A(net328),
    .B(_16438_),
    .C(_16454_),
    .Y(_16455_));
 OA21x2_ASAP7_75t_R _21867_ (.A1(_13355_),
    .A2(_16423_),
    .B(_16455_),
    .Y(_16456_));
 INVx2_ASAP7_75t_R _21868_ (.A(_16456_),
    .Y(_16457_));
 TAPCELL_ASAP7_75t_R TAP_1089 ();
 OA21x2_ASAP7_75t_R _21870_ (.A1(_00280_),
    .A2(_14543_),
    .B(_13521_),
    .Y(_16459_));
 TAPCELL_ASAP7_75t_R TAP_1088 ();
 OA21x2_ASAP7_75t_R _21872_ (.A1(net374),
    .A2(_15489_),
    .B(_16459_),
    .Y(_16461_));
 AOI21x1_ASAP7_75t_R _21873_ (.A1(_13474_),
    .A2(_16457_),
    .B(_16461_),
    .Y(_18425_));
 NAND2x1_ASAP7_75t_R _21874_ (.A(net393),
    .B(_01689_),
    .Y(_16462_));
 OA211x2_ASAP7_75t_R _21875_ (.A1(net393),
    .A2(_16394_),
    .B(_16462_),
    .C(net319),
    .Y(_16463_));
 AO21x1_ASAP7_75t_R _21876_ (.A1(_16393_),
    .A2(_13687_),
    .B(_16463_),
    .Y(_16464_));
 NAND2x1_ASAP7_75t_R _21877_ (.A(net390),
    .B(_00919_),
    .Y(_16465_));
 OA211x2_ASAP7_75t_R _21878_ (.A1(net390),
    .A2(_16407_),
    .B(_16465_),
    .C(_13649_),
    .Y(_16466_));
 NAND2x1_ASAP7_75t_R _21879_ (.A(net390),
    .B(_00918_),
    .Y(_16467_));
 OA211x2_ASAP7_75t_R _21880_ (.A1(net390),
    .A2(_16410_),
    .B(_16467_),
    .C(net419),
    .Y(_16468_));
 OR3x1_ASAP7_75t_R _21881_ (.A(_13636_),
    .B(_16466_),
    .C(_16468_),
    .Y(_16469_));
 NAND2x1_ASAP7_75t_R _21882_ (.A(net392),
    .B(_00927_),
    .Y(_16470_));
 OA211x2_ASAP7_75t_R _21883_ (.A1(net392),
    .A2(_16415_),
    .B(_16470_),
    .C(_13649_),
    .Y(_16471_));
 NAND2x1_ASAP7_75t_R _21884_ (.A(net392),
    .B(_00926_),
    .Y(_16472_));
 OA211x2_ASAP7_75t_R _21885_ (.A1(net392),
    .A2(_16418_),
    .B(_16472_),
    .C(net419),
    .Y(_16473_));
 OR3x1_ASAP7_75t_R _21886_ (.A(net381),
    .B(_16471_),
    .C(_16473_),
    .Y(_16474_));
 AO21x1_ASAP7_75t_R _21887_ (.A1(_16469_),
    .A2(_16474_),
    .B(net388),
    .Y(_16475_));
 NAND2x1_ASAP7_75t_R _21888_ (.A(net391),
    .B(_00922_),
    .Y(_16476_));
 OA211x2_ASAP7_75t_R _21889_ (.A1(net391),
    .A2(_16401_),
    .B(_16476_),
    .C(net427),
    .Y(_16477_));
 NAND2x1_ASAP7_75t_R _21890_ (.A(net390),
    .B(_00923_),
    .Y(_16478_));
 OA211x2_ASAP7_75t_R _21891_ (.A1(net390),
    .A2(_16398_),
    .B(_16478_),
    .C(_13649_),
    .Y(_16479_));
 OR3x1_ASAP7_75t_R _21892_ (.A(_14942_),
    .B(_16477_),
    .C(_16479_),
    .Y(_16480_));
 OA211x2_ASAP7_75t_R _21893_ (.A1(net315),
    .A2(_16464_),
    .B(_16475_),
    .C(_16480_),
    .Y(_16481_));
 INVx1_ASAP7_75t_R _21894_ (.A(_00935_),
    .Y(_16482_));
 NAND2x1_ASAP7_75t_R _21895_ (.A(net387),
    .B(_00931_),
    .Y(_16483_));
 OA211x2_ASAP7_75t_R _21896_ (.A1(net387),
    .A2(_16482_),
    .B(_16483_),
    .C(net393),
    .Y(_16484_));
 NAND2x1_ASAP7_75t_R _21897_ (.A(net387),
    .B(_00933_),
    .Y(_16485_));
 OA211x2_ASAP7_75t_R _21898_ (.A1(net387),
    .A2(_16447_),
    .B(_16485_),
    .C(_13675_),
    .Y(_16486_));
 OR3x1_ASAP7_75t_R _21899_ (.A(net2263),
    .B(_16484_),
    .C(_16486_),
    .Y(_16487_));
 INVx1_ASAP7_75t_R _21900_ (.A(_00934_),
    .Y(_16488_));
 NAND2x1_ASAP7_75t_R _21901_ (.A(net387),
    .B(_00930_),
    .Y(_16489_));
 OA211x2_ASAP7_75t_R _21902_ (.A1(net387),
    .A2(_16488_),
    .B(_16489_),
    .C(net393),
    .Y(_16490_));
 NAND2x1_ASAP7_75t_R _21903_ (.A(net387),
    .B(_00932_),
    .Y(_16491_));
 OA211x2_ASAP7_75t_R _21904_ (.A1(net387),
    .A2(_16450_),
    .B(_16491_),
    .C(_13675_),
    .Y(_16492_));
 OR3x1_ASAP7_75t_R _21905_ (.A(net319),
    .B(_16490_),
    .C(_16492_),
    .Y(_16493_));
 AND3x1_ASAP7_75t_R _21906_ (.A(net382),
    .B(_16487_),
    .C(_16493_),
    .Y(_16494_));
 NAND2x1_ASAP7_75t_R _21907_ (.A(net390),
    .B(_00938_),
    .Y(_16495_));
 OA211x2_ASAP7_75t_R _21908_ (.A1(net390),
    .A2(_16434_),
    .B(_16495_),
    .C(net388),
    .Y(_16496_));
 NAND2x1_ASAP7_75t_R _21909_ (.A(net390),
    .B(_00942_),
    .Y(_16497_));
 OA211x2_ASAP7_75t_R _21910_ (.A1(net390),
    .A2(_16427_),
    .B(_16497_),
    .C(_13630_),
    .Y(_16498_));
 OR3x1_ASAP7_75t_R _21911_ (.A(_13649_),
    .B(_16496_),
    .C(_16498_),
    .Y(_16499_));
 NAND2x1_ASAP7_75t_R _21912_ (.A(net390),
    .B(_00943_),
    .Y(_16500_));
 OA211x2_ASAP7_75t_R _21913_ (.A1(net390),
    .A2(_16424_),
    .B(_16500_),
    .C(_13630_),
    .Y(_16501_));
 NAND2x1_ASAP7_75t_R _21914_ (.A(net390),
    .B(_00939_),
    .Y(_16502_));
 OA211x2_ASAP7_75t_R _21915_ (.A1(net390),
    .A2(_16431_),
    .B(_16502_),
    .C(net388),
    .Y(_16503_));
 OR3x1_ASAP7_75t_R _21916_ (.A(net419),
    .B(_16501_),
    .C(_16503_),
    .Y(_16504_));
 AND3x1_ASAP7_75t_R _21917_ (.A(_13636_),
    .B(_16499_),
    .C(_16504_),
    .Y(_16505_));
 OR3x2_ASAP7_75t_R _21918_ (.A(_00286_),
    .B(_16494_),
    .C(_16505_),
    .Y(_16506_));
 OA211x2_ASAP7_75t_R _21919_ (.A1(_13626_),
    .A2(_16481_),
    .B(_16506_),
    .C(_13810_),
    .Y(_16507_));
 OAI22x1_ASAP7_75t_R _21920_ (.A1(_01621_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00214_),
    .Y(_16508_));
 NOR2x2_ASAP7_75t_R _21921_ (.A(_16507_),
    .B(_16508_),
    .Y(_18424_));
 XOR2x2_ASAP7_75t_R _21922_ (.A(_00947_),
    .B(_02229_),
    .Y(_16509_));
 INVx3_ASAP7_75t_R _21923_ (.A(_16509_),
    .Y(net161));
 AND2x2_ASAP7_75t_R _21924_ (.A(net2371),
    .B(_01688_),
    .Y(_16510_));
 AO21x1_ASAP7_75t_R _21925_ (.A1(net2260),
    .A2(_00950_),
    .B(_16510_),
    .Y(_16511_));
 OAI22x1_ASAP7_75t_R _21926_ (.A1(_00949_),
    .A2(_14184_),
    .B1(_16511_),
    .B2(net371),
    .Y(_16512_));
 INVx1_ASAP7_75t_R _21927_ (.A(_00958_),
    .Y(_16513_));
 NAND2x1_ASAP7_75t_R _21928_ (.A(net2373),
    .B(_00956_),
    .Y(_16514_));
 OA211x2_ASAP7_75t_R _21929_ (.A1(net2279),
    .A2(_16513_),
    .B(_16514_),
    .C(net324),
    .Y(_16515_));
 INVx1_ASAP7_75t_R _21930_ (.A(_00957_),
    .Y(_16516_));
 NAND2x1_ASAP7_75t_R _21931_ (.A(net2375),
    .B(_00955_),
    .Y(_16517_));
 OA211x2_ASAP7_75t_R _21932_ (.A1(net2279),
    .A2(_16516_),
    .B(_16517_),
    .C(net372),
    .Y(_16518_));
 OR3x1_ASAP7_75t_R _21933_ (.A(net330),
    .B(_16515_),
    .C(_16518_),
    .Y(_16519_));
 OA211x2_ASAP7_75t_R _21934_ (.A1(_13373_),
    .A2(_16512_),
    .B(_16519_),
    .C(net334),
    .Y(_16520_));
 INVx1_ASAP7_75t_R _21935_ (.A(_00959_),
    .Y(_16521_));
 NOR2x1_ASAP7_75t_R _21936_ (.A(net2371),
    .B(_00961_),
    .Y(_16522_));
 AO21x1_ASAP7_75t_R _21937_ (.A1(net2371),
    .A2(_16521_),
    .B(_16522_),
    .Y(_16523_));
 INVx1_ASAP7_75t_R _21938_ (.A(_00962_),
    .Y(_16524_));
 NAND2x1_ASAP7_75t_R _21939_ (.A(net2284),
    .B(_00960_),
    .Y(_16525_));
 OA211x2_ASAP7_75t_R _21940_ (.A1(net2294),
    .A2(_16524_),
    .B(_16525_),
    .C(net324),
    .Y(_16526_));
 AO21x1_ASAP7_75t_R _21941_ (.A1(net371),
    .A2(_16523_),
    .B(_16526_),
    .Y(_16527_));
 INVx1_ASAP7_75t_R _21942_ (.A(_00954_),
    .Y(_16528_));
 NAND2x1_ASAP7_75t_R _21943_ (.A(net2284),
    .B(_00952_),
    .Y(_16529_));
 OA211x2_ASAP7_75t_R _21944_ (.A1(net2294),
    .A2(_16528_),
    .B(_16529_),
    .C(net324),
    .Y(_16530_));
 INVx1_ASAP7_75t_R _21945_ (.A(_00953_),
    .Y(_16531_));
 NAND2x1_ASAP7_75t_R _21946_ (.A(net2284),
    .B(_00951_),
    .Y(_16532_));
 OA211x2_ASAP7_75t_R _21947_ (.A1(net2294),
    .A2(_16531_),
    .B(_16532_),
    .C(net371),
    .Y(_16533_));
 OR3x1_ASAP7_75t_R _21948_ (.A(_13373_),
    .B(_16530_),
    .C(_16533_),
    .Y(_16534_));
 OA211x2_ASAP7_75t_R _21949_ (.A1(net330),
    .A2(_16527_),
    .B(_16534_),
    .C(_13350_),
    .Y(_16535_));
 OR3x1_ASAP7_75t_R _21950_ (.A(_13355_),
    .B(_16520_),
    .C(_16535_),
    .Y(_16536_));
 INVx1_ASAP7_75t_R _21951_ (.A(_00974_),
    .Y(_16537_));
 NAND2x1_ASAP7_75t_R _21952_ (.A(net2282),
    .B(_00972_),
    .Y(_16538_));
 OA211x2_ASAP7_75t_R _21953_ (.A1(net2279),
    .A2(_16537_),
    .B(_16538_),
    .C(net324),
    .Y(_16539_));
 INVx1_ASAP7_75t_R _21954_ (.A(_00973_),
    .Y(_16540_));
 NAND2x1_ASAP7_75t_R _21955_ (.A(net2373),
    .B(_00971_),
    .Y(_16541_));
 OA211x2_ASAP7_75t_R _21956_ (.A1(net2279),
    .A2(_16540_),
    .B(_16541_),
    .C(net371),
    .Y(_16542_));
 OR3x1_ASAP7_75t_R _21957_ (.A(net330),
    .B(_16539_),
    .C(_16542_),
    .Y(_16543_));
 INVx1_ASAP7_75t_R _21958_ (.A(_00966_),
    .Y(_16544_));
 NAND2x1_ASAP7_75t_R _21959_ (.A(net2283),
    .B(_00964_),
    .Y(_16545_));
 OA211x2_ASAP7_75t_R _21960_ (.A1(net2279),
    .A2(_16544_),
    .B(_16545_),
    .C(net324),
    .Y(_16546_));
 INVx1_ASAP7_75t_R _21961_ (.A(_00965_),
    .Y(_16547_));
 NAND2x1_ASAP7_75t_R _21962_ (.A(net2283),
    .B(_00963_),
    .Y(_16548_));
 OA211x2_ASAP7_75t_R _21963_ (.A1(net2279),
    .A2(_16547_),
    .B(_16548_),
    .C(net371),
    .Y(_16549_));
 OR3x1_ASAP7_75t_R _21964_ (.A(_13373_),
    .B(_16546_),
    .C(_16549_),
    .Y(_16550_));
 AND3x1_ASAP7_75t_R _21965_ (.A(net334),
    .B(_16543_),
    .C(_16550_),
    .Y(_16551_));
 INVx1_ASAP7_75t_R _21966_ (.A(_00970_),
    .Y(_16552_));
 NAND2x1_ASAP7_75t_R _21967_ (.A(net2284),
    .B(_00968_),
    .Y(_16553_));
 OA211x2_ASAP7_75t_R _21968_ (.A1(net2371),
    .A2(_16552_),
    .B(_16553_),
    .C(net324),
    .Y(_16554_));
 INVx1_ASAP7_75t_R _21969_ (.A(_00969_),
    .Y(_16555_));
 NAND2x1_ASAP7_75t_R _21970_ (.A(net2284),
    .B(_00967_),
    .Y(_16556_));
 OA211x2_ASAP7_75t_R _21971_ (.A1(net2371),
    .A2(_16555_),
    .B(_16556_),
    .C(net371),
    .Y(_16557_));
 OR3x1_ASAP7_75t_R _21972_ (.A(_13373_),
    .B(_16554_),
    .C(_16557_),
    .Y(_16558_));
 INVx1_ASAP7_75t_R _21973_ (.A(_00978_),
    .Y(_16559_));
 NAND2x1_ASAP7_75t_R _21974_ (.A(net2373),
    .B(_00976_),
    .Y(_16560_));
 OA211x2_ASAP7_75t_R _21975_ (.A1(net2279),
    .A2(_16559_),
    .B(_16560_),
    .C(net324),
    .Y(_16561_));
 INVx1_ASAP7_75t_R _21976_ (.A(_00977_),
    .Y(_16562_));
 NAND2x1_ASAP7_75t_R _21977_ (.A(net2375),
    .B(_00975_),
    .Y(_16563_));
 OA211x2_ASAP7_75t_R _21978_ (.A1(net2279),
    .A2(_16562_),
    .B(_16563_),
    .C(net372),
    .Y(_16564_));
 OR3x1_ASAP7_75t_R _21979_ (.A(net330),
    .B(_16561_),
    .C(_16564_),
    .Y(_16565_));
 AND3x1_ASAP7_75t_R _21980_ (.A(_13350_),
    .B(_16558_),
    .C(_16565_),
    .Y(_16566_));
 OR3x1_ASAP7_75t_R _21981_ (.A(net327),
    .B(_16551_),
    .C(_16566_),
    .Y(_16567_));
 NAND2x2_ASAP7_75t_R _21982_ (.A(_16536_),
    .B(_16567_),
    .Y(_16568_));
 TAPCELL_ASAP7_75t_R TAP_1087 ();
 OA21x2_ASAP7_75t_R _21984_ (.A1(net2269),
    .A2(_15489_),
    .B(_16459_),
    .Y(_16570_));
 AO21x2_ASAP7_75t_R _21985_ (.A1(_13474_),
    .A2(net2181),
    .B(_16570_),
    .Y(_16571_));
 TAPCELL_ASAP7_75t_R TAP_1086 ();
 INVx1_ASAP7_75t_R _21987_ (.A(_16571_),
    .Y(_18430_));
 INVx1_ASAP7_75t_R _21988_ (.A(_00215_),
    .Y(\cs_registers_i.pc_id_i[21] ));
 NAND2x1_ASAP7_75t_R _21989_ (.A(net394),
    .B(_00968_),
    .Y(_16572_));
 OA211x2_ASAP7_75t_R _21990_ (.A1(net394),
    .A2(_16552_),
    .B(_16572_),
    .C(net317),
    .Y(_16573_));
 NAND2x1_ASAP7_75t_R _21991_ (.A(net394),
    .B(_00967_),
    .Y(_16574_));
 OA211x2_ASAP7_75t_R _21992_ (.A1(net394),
    .A2(_16555_),
    .B(_16574_),
    .C(net421),
    .Y(_16575_));
 OR3x1_ASAP7_75t_R _21993_ (.A(net383),
    .B(_16573_),
    .C(_16575_),
    .Y(_16576_));
 NAND2x1_ASAP7_75t_R _21994_ (.A(net394),
    .B(_00964_),
    .Y(_16577_));
 OA211x2_ASAP7_75t_R _21995_ (.A1(net394),
    .A2(_16544_),
    .B(_16577_),
    .C(net317),
    .Y(_16578_));
 NAND2x1_ASAP7_75t_R _21996_ (.A(net394),
    .B(_00963_),
    .Y(_16579_));
 OA211x2_ASAP7_75t_R _21997_ (.A1(net394),
    .A2(_16547_),
    .B(_16579_),
    .C(net421),
    .Y(_16580_));
 OR3x1_ASAP7_75t_R _21998_ (.A(net321),
    .B(_16578_),
    .C(_16580_),
    .Y(_16581_));
 NAND2x1_ASAP7_75t_R _21999_ (.A(net394),
    .B(_00952_),
    .Y(_16582_));
 OA211x2_ASAP7_75t_R _22000_ (.A1(net394),
    .A2(_16528_),
    .B(_16582_),
    .C(net317),
    .Y(_16583_));
 NAND2x1_ASAP7_75t_R _22001_ (.A(net394),
    .B(_00951_),
    .Y(_16584_));
 OA211x2_ASAP7_75t_R _22002_ (.A1(net394),
    .A2(_16531_),
    .B(_16584_),
    .C(net421),
    .Y(_16585_));
 OR3x1_ASAP7_75t_R _22003_ (.A(net312),
    .B(_16583_),
    .C(_16585_),
    .Y(_16586_));
 INVx1_ASAP7_75t_R _22004_ (.A(_00950_),
    .Y(_16587_));
 NAND2x1_ASAP7_75t_R _22005_ (.A(net399),
    .B(_01688_),
    .Y(_16588_));
 OA211x2_ASAP7_75t_R _22006_ (.A1(net399),
    .A2(_16587_),
    .B(_16588_),
    .C(net317),
    .Y(_16589_));
 NOR2x1_ASAP7_75t_R _22007_ (.A(net399),
    .B(_00949_),
    .Y(_16590_));
 AO21x1_ASAP7_75t_R _22008_ (.A1(net421),
    .A2(_16590_),
    .B(_14005_),
    .Y(_16591_));
 OA21x2_ASAP7_75t_R _22009_ (.A1(_16589_),
    .A2(_16591_),
    .B(net377),
    .Y(_16592_));
 AO32x1_ASAP7_75t_R _22010_ (.A1(_13626_),
    .A2(_16576_),
    .A3(_16581_),
    .B1(_16586_),
    .B2(_16592_),
    .Y(_16593_));
 NOR2x1_ASAP7_75t_R _22011_ (.A(net394),
    .B(_00961_),
    .Y(_16594_));
 AO21x1_ASAP7_75t_R _22012_ (.A1(net394),
    .A2(_16521_),
    .B(_16594_),
    .Y(_16595_));
 NAND2x1_ASAP7_75t_R _22013_ (.A(net394),
    .B(_00960_),
    .Y(_16596_));
 OA211x2_ASAP7_75t_R _22014_ (.A1(net394),
    .A2(_16524_),
    .B(_16596_),
    .C(net317),
    .Y(_16597_));
 AO21x1_ASAP7_75t_R _22015_ (.A1(net421),
    .A2(_16595_),
    .B(_16597_),
    .Y(_16598_));
 NAND2x1_ASAP7_75t_R _22016_ (.A(net394),
    .B(_00956_),
    .Y(_16599_));
 OA211x2_ASAP7_75t_R _22017_ (.A1(net394),
    .A2(_16513_),
    .B(_16599_),
    .C(net317),
    .Y(_16600_));
 NAND2x1_ASAP7_75t_R _22018_ (.A(net394),
    .B(_00955_),
    .Y(_16601_));
 OA211x2_ASAP7_75t_R _22019_ (.A1(net394),
    .A2(_16516_),
    .B(_16601_),
    .C(net421),
    .Y(_16602_));
 OA21x2_ASAP7_75t_R _22020_ (.A1(_16600_),
    .A2(_16602_),
    .B(net383),
    .Y(_16603_));
 AO21x1_ASAP7_75t_R _22021_ (.A1(net321),
    .A2(_16598_),
    .B(_16603_),
    .Y(_16604_));
 AND2x2_ASAP7_75t_R _22022_ (.A(_16586_),
    .B(_16592_),
    .Y(_16605_));
 NAND2x1_ASAP7_75t_R _22023_ (.A(net403),
    .B(_00972_),
    .Y(_16606_));
 OA211x2_ASAP7_75t_R _22024_ (.A1(net403),
    .A2(_16537_),
    .B(_16606_),
    .C(net317),
    .Y(_16607_));
 NAND2x1_ASAP7_75t_R _22025_ (.A(net403),
    .B(_00971_),
    .Y(_16608_));
 OA211x2_ASAP7_75t_R _22026_ (.A1(net403),
    .A2(_16540_),
    .B(_16608_),
    .C(net420),
    .Y(_16609_));
 OR3x1_ASAP7_75t_R _22027_ (.A(net321),
    .B(_16607_),
    .C(_16609_),
    .Y(_16610_));
 NAND2x1_ASAP7_75t_R _22028_ (.A(net394),
    .B(_00976_),
    .Y(_16611_));
 OA211x2_ASAP7_75t_R _22029_ (.A1(net394),
    .A2(_16559_),
    .B(_16611_),
    .C(net317),
    .Y(_16612_));
 NAND2x1_ASAP7_75t_R _22030_ (.A(net394),
    .B(_00975_),
    .Y(_16613_));
 OA211x2_ASAP7_75t_R _22031_ (.A1(net394),
    .A2(_16562_),
    .B(_16613_),
    .C(net420),
    .Y(_16614_));
 OR3x1_ASAP7_75t_R _22032_ (.A(net383),
    .B(_16612_),
    .C(_16614_),
    .Y(_16615_));
 AND3x1_ASAP7_75t_R _22033_ (.A(_14780_),
    .B(_16610_),
    .C(_16615_),
    .Y(_16616_));
 AO221x2_ASAP7_75t_R _22034_ (.A1(net380),
    .A2(_16593_),
    .B1(_16604_),
    .B2(_16605_),
    .C(_16616_),
    .Y(_16617_));
 OA211x2_ASAP7_75t_R _22035_ (.A1(_13788_),
    .A2(_13806_),
    .B(_00215_),
    .C(_13807_),
    .Y(_16618_));
 OAI22x1_ASAP7_75t_R _22036_ (.A1(_01620_),
    .A2(_13807_),
    .B1(_14988_),
    .B2(_16618_),
    .Y(_16619_));
 OA21x2_ASAP7_75t_R _22037_ (.A1(_15112_),
    .A2(_16617_),
    .B(_16619_),
    .Y(_16620_));
 TAPCELL_ASAP7_75t_R TAP_1085 ();
 INVx2_ASAP7_75t_R _22039_ (.A(_16620_),
    .Y(_18429_));
 AND2x2_ASAP7_75t_R _22040_ (.A(net342),
    .B(_01687_),
    .Y(_16621_));
 AO21x1_ASAP7_75t_R _22041_ (.A1(net326),
    .A2(_00982_),
    .B(_16621_),
    .Y(_16622_));
 OAI22x1_ASAP7_75t_R _22042_ (.A1(_00981_),
    .A2(net311),
    .B1(_16622_),
    .B2(net370),
    .Y(_16623_));
 INVx1_ASAP7_75t_R _22043_ (.A(_00990_),
    .Y(_16624_));
 NAND2x1_ASAP7_75t_R _22044_ (.A(net345),
    .B(_00988_),
    .Y(_16625_));
 OA211x2_ASAP7_75t_R _22045_ (.A1(net345),
    .A2(_16624_),
    .B(_16625_),
    .C(_13376_),
    .Y(_16626_));
 INVx1_ASAP7_75t_R _22046_ (.A(_00989_),
    .Y(_16627_));
 NAND2x1_ASAP7_75t_R _22047_ (.A(net345),
    .B(_00987_),
    .Y(_16628_));
 OA211x2_ASAP7_75t_R _22048_ (.A1(net345),
    .A2(_16627_),
    .B(_16628_),
    .C(net376),
    .Y(_16629_));
 OR3x1_ASAP7_75t_R _22049_ (.A(net332),
    .B(_16626_),
    .C(_16629_),
    .Y(_16630_));
 OA211x2_ASAP7_75t_R _22050_ (.A1(_13373_),
    .A2(_16623_),
    .B(_16630_),
    .C(net338),
    .Y(_16631_));
 INVx1_ASAP7_75t_R _22051_ (.A(_00986_),
    .Y(_16632_));
 NAND2x1_ASAP7_75t_R _22052_ (.A(net344),
    .B(_00984_),
    .Y(_16633_));
 OA211x2_ASAP7_75t_R _22053_ (.A1(net344),
    .A2(_16632_),
    .B(_16633_),
    .C(_13376_),
    .Y(_16634_));
 INVx1_ASAP7_75t_R _22054_ (.A(_00985_),
    .Y(_16635_));
 NAND2x1_ASAP7_75t_R _22055_ (.A(net344),
    .B(_00983_),
    .Y(_16636_));
 OA211x2_ASAP7_75t_R _22056_ (.A1(net344),
    .A2(_16635_),
    .B(_16636_),
    .C(net2314),
    .Y(_16637_));
 OR3x1_ASAP7_75t_R _22057_ (.A(_13373_),
    .B(_16634_),
    .C(_16637_),
    .Y(_16638_));
 INVx1_ASAP7_75t_R _22058_ (.A(_00994_),
    .Y(_16639_));
 NAND2x1_ASAP7_75t_R _22059_ (.A(net344),
    .B(_00992_),
    .Y(_16640_));
 OA211x2_ASAP7_75t_R _22060_ (.A1(net344),
    .A2(_16639_),
    .B(_16640_),
    .C(_13376_),
    .Y(_16641_));
 INVx1_ASAP7_75t_R _22061_ (.A(_00993_),
    .Y(_16642_));
 NAND2x1_ASAP7_75t_R _22062_ (.A(net344),
    .B(_00991_),
    .Y(_16643_));
 OA211x2_ASAP7_75t_R _22063_ (.A1(net344),
    .A2(_16642_),
    .B(_16643_),
    .C(net2315),
    .Y(_16644_));
 OR3x1_ASAP7_75t_R _22064_ (.A(_00245_),
    .B(_16641_),
    .C(_16644_),
    .Y(_16645_));
 AND3x1_ASAP7_75t_R _22065_ (.A(_13350_),
    .B(_16638_),
    .C(_16645_),
    .Y(_16646_));
 OR3x4_ASAP7_75t_R _22066_ (.A(_13355_),
    .B(_16631_),
    .C(_16646_),
    .Y(_16647_));
 INVx1_ASAP7_75t_R _22067_ (.A(_01002_),
    .Y(_16648_));
 NAND2x1_ASAP7_75t_R _22068_ (.A(net339),
    .B(_01000_),
    .Y(_16649_));
 OA211x2_ASAP7_75t_R _22069_ (.A1(net339),
    .A2(_16648_),
    .B(_16649_),
    .C(net323),
    .Y(_16650_));
 INVx1_ASAP7_75t_R _22070_ (.A(_01001_),
    .Y(_16651_));
 NAND2x1_ASAP7_75t_R _22071_ (.A(net339),
    .B(_00999_),
    .Y(_16652_));
 OA211x2_ASAP7_75t_R _22072_ (.A1(net339),
    .A2(_16651_),
    .B(_16652_),
    .C(net370),
    .Y(_16653_));
 OR3x1_ASAP7_75t_R _22073_ (.A(net337),
    .B(_16650_),
    .C(_16653_),
    .Y(_16654_));
 INVx1_ASAP7_75t_R _22074_ (.A(_00998_),
    .Y(_16655_));
 NAND2x1_ASAP7_75t_R _22075_ (.A(net340),
    .B(_00996_),
    .Y(_16656_));
 OA211x2_ASAP7_75t_R _22076_ (.A1(net340),
    .A2(_16655_),
    .B(_16656_),
    .C(_13376_),
    .Y(_16657_));
 INVx1_ASAP7_75t_R _22077_ (.A(_00997_),
    .Y(_16658_));
 NAND2x1_ASAP7_75t_R _22078_ (.A(net340),
    .B(_00995_),
    .Y(_16659_));
 OA211x2_ASAP7_75t_R _22079_ (.A1(net340),
    .A2(_16658_),
    .B(_16659_),
    .C(net370),
    .Y(_16660_));
 OR3x1_ASAP7_75t_R _22080_ (.A(_13350_),
    .B(_16657_),
    .C(_16660_),
    .Y(_16661_));
 AND3x1_ASAP7_75t_R _22081_ (.A(net332),
    .B(_16654_),
    .C(_16661_),
    .Y(_16662_));
 INVx1_ASAP7_75t_R _22082_ (.A(_01010_),
    .Y(_16663_));
 NAND2x1_ASAP7_75t_R _22083_ (.A(net343),
    .B(_01008_),
    .Y(_16664_));
 OA211x2_ASAP7_75t_R _22084_ (.A1(net343),
    .A2(_16663_),
    .B(_16664_),
    .C(_13376_),
    .Y(_16665_));
 INVx1_ASAP7_75t_R _22085_ (.A(_01009_),
    .Y(_16666_));
 NAND2x1_ASAP7_75t_R _22086_ (.A(net344),
    .B(_01007_),
    .Y(_16667_));
 OA211x2_ASAP7_75t_R _22087_ (.A1(net344),
    .A2(_16666_),
    .B(_16667_),
    .C(net2315),
    .Y(_16668_));
 OR3x1_ASAP7_75t_R _22088_ (.A(net338),
    .B(_16665_),
    .C(_16668_),
    .Y(_16669_));
 INVx1_ASAP7_75t_R _22089_ (.A(_01006_),
    .Y(_16670_));
 NAND2x1_ASAP7_75t_R _22090_ (.A(net343),
    .B(_01004_),
    .Y(_16671_));
 OA211x2_ASAP7_75t_R _22091_ (.A1(net343),
    .A2(_16670_),
    .B(_16671_),
    .C(_13376_),
    .Y(_16672_));
 INVx1_ASAP7_75t_R _22092_ (.A(_01005_),
    .Y(_16673_));
 NAND2x1_ASAP7_75t_R _22093_ (.A(net343),
    .B(_01003_),
    .Y(_16674_));
 OA211x2_ASAP7_75t_R _22094_ (.A1(net343),
    .A2(_16673_),
    .B(_16674_),
    .C(net2314),
    .Y(_16675_));
 OR3x1_ASAP7_75t_R _22095_ (.A(_13350_),
    .B(_16672_),
    .C(_16675_),
    .Y(_16676_));
 AND3x1_ASAP7_75t_R _22096_ (.A(_13373_),
    .B(_16669_),
    .C(_16676_),
    .Y(_16677_));
 OR3x4_ASAP7_75t_R _22097_ (.A(net328),
    .B(_16662_),
    .C(_16677_),
    .Y(_16678_));
 NAND2x2_ASAP7_75t_R _22098_ (.A(_16647_),
    .B(_16678_),
    .Y(_16679_));
 OA21x2_ASAP7_75t_R _22099_ (.A1(net336),
    .A2(_15489_),
    .B(_16459_),
    .Y(_16680_));
 AOI21x1_ASAP7_75t_R _22100_ (.A1(_13474_),
    .A2(_16679_),
    .B(_16680_),
    .Y(_18434_));
 NAND2x1_ASAP7_75t_R _22101_ (.A(_00217_),
    .B(_13993_),
    .Y(_16681_));
 NAND2x1_ASAP7_75t_R _22102_ (.A(net390),
    .B(_01004_),
    .Y(_16682_));
 OA211x2_ASAP7_75t_R _22103_ (.A1(net390),
    .A2(_16670_),
    .B(_16682_),
    .C(_13649_),
    .Y(_16683_));
 NAND2x1_ASAP7_75t_R _22104_ (.A(net390),
    .B(_01003_),
    .Y(_16684_));
 OA211x2_ASAP7_75t_R _22105_ (.A1(net390),
    .A2(_16673_),
    .B(_16684_),
    .C(net419),
    .Y(_16685_));
 OR3x1_ASAP7_75t_R _22106_ (.A(_13630_),
    .B(_16683_),
    .C(_16685_),
    .Y(_16686_));
 NAND2x1_ASAP7_75t_R _22107_ (.A(net390),
    .B(_01008_),
    .Y(_16687_));
 OA211x2_ASAP7_75t_R _22108_ (.A1(net390),
    .A2(_16663_),
    .B(_16687_),
    .C(_13649_),
    .Y(_16688_));
 NAND2x1_ASAP7_75t_R _22109_ (.A(net392),
    .B(_01007_),
    .Y(_16689_));
 OA211x2_ASAP7_75t_R _22110_ (.A1(net392),
    .A2(_16666_),
    .B(_16689_),
    .C(net419),
    .Y(_16690_));
 OR3x1_ASAP7_75t_R _22111_ (.A(net388),
    .B(_16688_),
    .C(_16690_),
    .Y(_16691_));
 AO21x1_ASAP7_75t_R _22112_ (.A1(_16686_),
    .A2(_16691_),
    .B(net381),
    .Y(_16692_));
 NAND2x1_ASAP7_75t_R _22113_ (.A(net415),
    .B(_00999_),
    .Y(_16693_));
 OA211x2_ASAP7_75t_R _22114_ (.A1(net415),
    .A2(_16651_),
    .B(_16693_),
    .C(net426),
    .Y(_16694_));
 NAND2x1_ASAP7_75t_R _22115_ (.A(net417),
    .B(_01000_),
    .Y(_16695_));
 OA211x2_ASAP7_75t_R _22116_ (.A1(net415),
    .A2(_16648_),
    .B(_16695_),
    .C(net319),
    .Y(_16696_));
 OR3x1_ASAP7_75t_R _22117_ (.A(_14015_),
    .B(_16694_),
    .C(_16696_),
    .Y(_16697_));
 NAND2x1_ASAP7_75t_R _22118_ (.A(net393),
    .B(_00995_),
    .Y(_16698_));
 OA211x2_ASAP7_75t_R _22119_ (.A1(net393),
    .A2(_16658_),
    .B(_16698_),
    .C(net427),
    .Y(_16699_));
 NAND2x1_ASAP7_75t_R _22120_ (.A(net393),
    .B(_00996_),
    .Y(_16700_));
 OA211x2_ASAP7_75t_R _22121_ (.A1(net393),
    .A2(_16655_),
    .B(_16700_),
    .C(net319),
    .Y(_16701_));
 OR3x1_ASAP7_75t_R _22122_ (.A(net315),
    .B(_16699_),
    .C(_16701_),
    .Y(_16702_));
 AND3x1_ASAP7_75t_R _22123_ (.A(_13626_),
    .B(_16697_),
    .C(_16702_),
    .Y(_16703_));
 NAND2x1_ASAP7_75t_R _22124_ (.A(net392),
    .B(_00984_),
    .Y(_16704_));
 OA211x2_ASAP7_75t_R _22125_ (.A1(net392),
    .A2(_16632_),
    .B(_16704_),
    .C(_13649_),
    .Y(_16705_));
 NAND2x1_ASAP7_75t_R _22126_ (.A(net392),
    .B(_00983_),
    .Y(_16706_));
 OA211x2_ASAP7_75t_R _22127_ (.A1(net392),
    .A2(_16635_),
    .B(_16706_),
    .C(net419),
    .Y(_16707_));
 OR3x1_ASAP7_75t_R _22128_ (.A(_13636_),
    .B(_16705_),
    .C(_16707_),
    .Y(_16708_));
 NAND2x1_ASAP7_75t_R _22129_ (.A(net392),
    .B(_00992_),
    .Y(_16709_));
 OA211x2_ASAP7_75t_R _22130_ (.A1(net392),
    .A2(_16639_),
    .B(_16709_),
    .C(_13649_),
    .Y(_16710_));
 NAND2x1_ASAP7_75t_R _22131_ (.A(net392),
    .B(_00991_),
    .Y(_16711_));
 OA211x2_ASAP7_75t_R _22132_ (.A1(net392),
    .A2(_16642_),
    .B(_16711_),
    .C(net419),
    .Y(_16712_));
 OR3x1_ASAP7_75t_R _22133_ (.A(net381),
    .B(_16710_),
    .C(_16712_),
    .Y(_16713_));
 AO21x1_ASAP7_75t_R _22134_ (.A1(_16708_),
    .A2(_16713_),
    .B(net388),
    .Y(_04504_));
 AND2x2_ASAP7_75t_R _22135_ (.A(net389),
    .B(_01687_),
    .Y(_04505_));
 AO21x1_ASAP7_75t_R _22136_ (.A1(_13675_),
    .A2(_00982_),
    .B(_04505_),
    .Y(_04506_));
 OAI22x1_ASAP7_75t_R _22137_ (.A1(_00981_),
    .A2(net2290),
    .B1(_04506_),
    .B2(net427),
    .Y(_04507_));
 NAND2x1_ASAP7_75t_R _22138_ (.A(net389),
    .B(_00988_),
    .Y(_04508_));
 OA211x2_ASAP7_75t_R _22139_ (.A1(net391),
    .A2(_16624_),
    .B(_04508_),
    .C(net319),
    .Y(_04509_));
 NAND2x1_ASAP7_75t_R _22140_ (.A(net391),
    .B(_00987_),
    .Y(_04510_));
 OA211x2_ASAP7_75t_R _22141_ (.A1(net391),
    .A2(_16627_),
    .B(_04510_),
    .C(net427),
    .Y(_04511_));
 OR3x1_ASAP7_75t_R _22142_ (.A(_14942_),
    .B(_04509_),
    .C(_04511_),
    .Y(_04512_));
 OA211x2_ASAP7_75t_R _22143_ (.A1(net315),
    .A2(_04507_),
    .B(_04512_),
    .C(_00286_),
    .Y(_04513_));
 AO221x2_ASAP7_75t_R _22144_ (.A1(_16692_),
    .A2(_16703_),
    .B1(_04504_),
    .B2(_04513_),
    .C(_13993_),
    .Y(_04514_));
 INVx1_ASAP7_75t_R _22145_ (.A(_01619_),
    .Y(_04515_));
 AO32x2_ASAP7_75t_R _22146_ (.A1(_13794_),
    .A2(_16681_),
    .A3(_04514_),
    .B1(_13450_),
    .B2(_04515_),
    .Y(_04516_));
 TAPCELL_ASAP7_75t_R TAP_1084 ();
 INVx3_ASAP7_75t_R _22148_ (.A(_04516_),
    .Y(_18435_));
 XNOR2x2_ASAP7_75t_R _22149_ (.A(_01014_),
    .B(_01012_),
    .Y(_04517_));
 INVx6_ASAP7_75t_R _22150_ (.A(_04517_),
    .Y(net163));
 AND2x2_ASAP7_75t_R _22151_ (.A(net348),
    .B(_01686_),
    .Y(_04518_));
 AO21x1_ASAP7_75t_R _22152_ (.A1(_13359_),
    .A2(_01016_),
    .B(_04518_),
    .Y(_04519_));
 OAI22x1_ASAP7_75t_R _22153_ (.A1(_01015_),
    .A2(net311),
    .B1(_04519_),
    .B2(net375),
    .Y(_04520_));
 INVx1_ASAP7_75t_R _22154_ (.A(_01024_),
    .Y(_04521_));
 NAND2x1_ASAP7_75t_R _22155_ (.A(net348),
    .B(_01022_),
    .Y(_04522_));
 OA211x2_ASAP7_75t_R _22156_ (.A1(net348),
    .A2(_04521_),
    .B(_04522_),
    .C(net325),
    .Y(_04523_));
 INVx1_ASAP7_75t_R _22157_ (.A(_01023_),
    .Y(_04524_));
 NAND2x1_ASAP7_75t_R _22158_ (.A(net348),
    .B(_01021_),
    .Y(_04525_));
 OA211x2_ASAP7_75t_R _22159_ (.A1(net348),
    .A2(_04524_),
    .B(_04525_),
    .C(net375),
    .Y(_04526_));
 OR3x1_ASAP7_75t_R _22160_ (.A(net331),
    .B(_04523_),
    .C(_04526_),
    .Y(_04527_));
 OA211x2_ASAP7_75t_R _22161_ (.A1(_13373_),
    .A2(_04520_),
    .B(_04527_),
    .C(net337),
    .Y(_04528_));
 INVx1_ASAP7_75t_R _22162_ (.A(_01020_),
    .Y(_04529_));
 NAND2x1_ASAP7_75t_R _22163_ (.A(net347),
    .B(_01018_),
    .Y(_04530_));
 OA211x2_ASAP7_75t_R _22164_ (.A1(net347),
    .A2(_04529_),
    .B(_04530_),
    .C(net325),
    .Y(_04531_));
 INVx1_ASAP7_75t_R _22165_ (.A(_01019_),
    .Y(_04532_));
 NAND2x1_ASAP7_75t_R _22166_ (.A(net347),
    .B(_01017_),
    .Y(_04533_));
 OA211x2_ASAP7_75t_R _22167_ (.A1(net347),
    .A2(_04532_),
    .B(_04533_),
    .C(net375),
    .Y(_04534_));
 OR3x1_ASAP7_75t_R _22168_ (.A(_13373_),
    .B(_04531_),
    .C(_04534_),
    .Y(_04535_));
 INVx1_ASAP7_75t_R _22169_ (.A(_01028_),
    .Y(_04536_));
 NAND2x1_ASAP7_75t_R _22170_ (.A(net347),
    .B(_01026_),
    .Y(_04537_));
 OA211x2_ASAP7_75t_R _22171_ (.A1(net347),
    .A2(_04536_),
    .B(_04537_),
    .C(net325),
    .Y(_04538_));
 INVx1_ASAP7_75t_R _22172_ (.A(_01027_),
    .Y(_04539_));
 NAND2x1_ASAP7_75t_R _22173_ (.A(net348),
    .B(_01025_),
    .Y(_04540_));
 OA211x2_ASAP7_75t_R _22174_ (.A1(net348),
    .A2(_04539_),
    .B(_04540_),
    .C(net369),
    .Y(_04541_));
 OR3x1_ASAP7_75t_R _22175_ (.A(net331),
    .B(_04538_),
    .C(_04541_),
    .Y(_04542_));
 AND3x1_ASAP7_75t_R _22176_ (.A(_13350_),
    .B(_04535_),
    .C(_04542_),
    .Y(_04543_));
 OR3x1_ASAP7_75t_R _22177_ (.A(_13355_),
    .B(_04528_),
    .C(_04543_),
    .Y(_04544_));
 INVx1_ASAP7_75t_R _22178_ (.A(_01036_),
    .Y(_04545_));
 NAND2x1_ASAP7_75t_R _22179_ (.A(net352),
    .B(_01034_),
    .Y(_04546_));
 OA211x2_ASAP7_75t_R _22180_ (.A1(net352),
    .A2(_04545_),
    .B(_04546_),
    .C(net325),
    .Y(_04547_));
 INVx1_ASAP7_75t_R _22181_ (.A(_01035_),
    .Y(_04548_));
 NAND2x1_ASAP7_75t_R _22182_ (.A(net352),
    .B(_01033_),
    .Y(_04549_));
 OA211x2_ASAP7_75t_R _22183_ (.A1(net352),
    .A2(_04548_),
    .B(_04549_),
    .C(net375),
    .Y(_04550_));
 OR3x1_ASAP7_75t_R _22184_ (.A(_13373_),
    .B(_04547_),
    .C(_04550_),
    .Y(_04551_));
 INVx1_ASAP7_75t_R _22185_ (.A(_01044_),
    .Y(_04552_));
 NAND2x1_ASAP7_75t_R _22186_ (.A(net352),
    .B(_01042_),
    .Y(_04553_));
 OA211x2_ASAP7_75t_R _22187_ (.A1(net352),
    .A2(_04552_),
    .B(_04553_),
    .C(net325),
    .Y(_04554_));
 INVx1_ASAP7_75t_R _22188_ (.A(_01043_),
    .Y(_04555_));
 NAND2x1_ASAP7_75t_R _22189_ (.A(net352),
    .B(_01041_),
    .Y(_04556_));
 OA211x2_ASAP7_75t_R _22190_ (.A1(net352),
    .A2(_04555_),
    .B(_04556_),
    .C(net375),
    .Y(_04557_));
 OR3x1_ASAP7_75t_R _22191_ (.A(net331),
    .B(_04554_),
    .C(_04557_),
    .Y(_04558_));
 AND3x1_ASAP7_75t_R _22192_ (.A(_13350_),
    .B(_04551_),
    .C(_04558_),
    .Y(_04559_));
 INVx1_ASAP7_75t_R _22193_ (.A(_01040_),
    .Y(_04560_));
 NAND2x1_ASAP7_75t_R _22194_ (.A(net351),
    .B(_01038_),
    .Y(_04561_));
 OA211x2_ASAP7_75t_R _22195_ (.A1(net351),
    .A2(_04560_),
    .B(_04561_),
    .C(net325),
    .Y(_04562_));
 INVx1_ASAP7_75t_R _22196_ (.A(_01039_),
    .Y(_04563_));
 NAND2x1_ASAP7_75t_R _22197_ (.A(net351),
    .B(_01037_),
    .Y(_04564_));
 OA211x2_ASAP7_75t_R _22198_ (.A1(net351),
    .A2(_04563_),
    .B(_04564_),
    .C(net375),
    .Y(_04565_));
 OR3x1_ASAP7_75t_R _22199_ (.A(net331),
    .B(_04562_),
    .C(_04565_),
    .Y(_04566_));
 INVx1_ASAP7_75t_R _22200_ (.A(_01032_),
    .Y(_04567_));
 NAND2x1_ASAP7_75t_R _22201_ (.A(net351),
    .B(_01030_),
    .Y(_04568_));
 OA211x2_ASAP7_75t_R _22202_ (.A1(net351),
    .A2(_04567_),
    .B(_04568_),
    .C(net325),
    .Y(_04569_));
 INVx1_ASAP7_75t_R _22203_ (.A(_01031_),
    .Y(_04570_));
 NAND2x1_ASAP7_75t_R _22204_ (.A(net351),
    .B(_01029_),
    .Y(_04571_));
 OA211x2_ASAP7_75t_R _22205_ (.A1(net351),
    .A2(_04570_),
    .B(_04571_),
    .C(net375),
    .Y(_04572_));
 OR3x1_ASAP7_75t_R _22206_ (.A(_13373_),
    .B(_04569_),
    .C(_04572_),
    .Y(_04573_));
 AND3x1_ASAP7_75t_R _22207_ (.A(net335),
    .B(_04566_),
    .C(_04573_),
    .Y(_04574_));
 OR3x1_ASAP7_75t_R _22208_ (.A(net327),
    .B(_04559_),
    .C(_04574_),
    .Y(_04575_));
 AND2x6_ASAP7_75t_R _22209_ (.A(_04544_),
    .B(_04575_),
    .Y(_04576_));
 INVx2_ASAP7_75t_R _22210_ (.A(_04576_),
    .Y(_04577_));
 OA21x2_ASAP7_75t_R _22211_ (.A1(net333),
    .A2(_15489_),
    .B(_16459_),
    .Y(_04578_));
 AOI21x1_ASAP7_75t_R _22212_ (.A1(_13474_),
    .A2(_04577_),
    .B(_04578_),
    .Y(_18439_));
 XOR2x1_ASAP7_75t_R _22213_ (.A(_13620_),
    .Y(_04579_),
    .B(_18439_));
 NAND2x1_ASAP7_75t_R _22214_ (.A(net396),
    .B(_01037_),
    .Y(_04580_));
 OA211x2_ASAP7_75t_R _22215_ (.A1(net396),
    .A2(_04563_),
    .B(_04580_),
    .C(net386),
    .Y(_04581_));
 NAND2x1_ASAP7_75t_R _22216_ (.A(net396),
    .B(_01041_),
    .Y(_04582_));
 OA211x2_ASAP7_75t_R _22217_ (.A1(net396),
    .A2(_04555_),
    .B(_04582_),
    .C(net321),
    .Y(_04583_));
 OR3x1_ASAP7_75t_R _22218_ (.A(_13649_),
    .B(_04581_),
    .C(_04583_),
    .Y(_04584_));
 NAND2x1_ASAP7_75t_R _22219_ (.A(net396),
    .B(_01038_),
    .Y(_04585_));
 OA211x2_ASAP7_75t_R _22220_ (.A1(net396),
    .A2(_04560_),
    .B(_04585_),
    .C(net386),
    .Y(_04586_));
 NAND2x1_ASAP7_75t_R _22221_ (.A(net396),
    .B(_01042_),
    .Y(_04587_));
 OA211x2_ASAP7_75t_R _22222_ (.A1(net396),
    .A2(_04552_),
    .B(_04587_),
    .C(net321),
    .Y(_04588_));
 OR3x1_ASAP7_75t_R _22223_ (.A(net424),
    .B(_04586_),
    .C(_04588_),
    .Y(_04589_));
 AND3x1_ASAP7_75t_R _22224_ (.A(_13636_),
    .B(_04584_),
    .C(_04589_),
    .Y(_04590_));
 NAND2x1_ASAP7_75t_R _22225_ (.A(net396),
    .B(_01029_),
    .Y(_04591_));
 OA211x2_ASAP7_75t_R _22226_ (.A1(net396),
    .A2(_04570_),
    .B(_04591_),
    .C(net386),
    .Y(_04592_));
 NAND2x1_ASAP7_75t_R _22227_ (.A(net398),
    .B(_01033_),
    .Y(_04593_));
 OA211x2_ASAP7_75t_R _22228_ (.A1(net398),
    .A2(_04548_),
    .B(_04593_),
    .C(net321),
    .Y(_04594_));
 OR3x1_ASAP7_75t_R _22229_ (.A(_13649_),
    .B(_04592_),
    .C(_04594_),
    .Y(_04595_));
 NAND2x1_ASAP7_75t_R _22230_ (.A(net396),
    .B(_01030_),
    .Y(_04596_));
 OA211x2_ASAP7_75t_R _22231_ (.A1(net396),
    .A2(_04567_),
    .B(_04596_),
    .C(net386),
    .Y(_04597_));
 NAND2x1_ASAP7_75t_R _22232_ (.A(net398),
    .B(_01034_),
    .Y(_04598_));
 OA211x2_ASAP7_75t_R _22233_ (.A1(net398),
    .A2(_04545_),
    .B(_04598_),
    .C(net321),
    .Y(_04599_));
 OR3x1_ASAP7_75t_R _22234_ (.A(net424),
    .B(_04597_),
    .C(_04599_),
    .Y(_04600_));
 AND3x1_ASAP7_75t_R _22235_ (.A(net382),
    .B(_04595_),
    .C(_04600_),
    .Y(_04601_));
 OR2x2_ASAP7_75t_R _22236_ (.A(_04590_),
    .B(_04601_),
    .Y(_04602_));
 NAND2x1_ASAP7_75t_R _22237_ (.A(net410),
    .B(_01018_),
    .Y(_04603_));
 OA211x2_ASAP7_75t_R _22238_ (.A1(net410),
    .A2(_04529_),
    .B(_04603_),
    .C(_13649_),
    .Y(_04604_));
 NAND2x1_ASAP7_75t_R _22239_ (.A(net412),
    .B(_01017_),
    .Y(_04605_));
 OA211x2_ASAP7_75t_R _22240_ (.A1(net412),
    .A2(_04532_),
    .B(_04605_),
    .C(net426),
    .Y(_04606_));
 INVx1_ASAP7_75t_R _22241_ (.A(_01016_),
    .Y(_04607_));
 NAND2x1_ASAP7_75t_R _22242_ (.A(net412),
    .B(_01686_),
    .Y(_04608_));
 OA211x2_ASAP7_75t_R _22243_ (.A1(net412),
    .A2(_04607_),
    .B(_04608_),
    .C(net319),
    .Y(_04609_));
 NOR2x1_ASAP7_75t_R _22244_ (.A(_01015_),
    .B(net2290),
    .Y(_04610_));
 OA33x2_ASAP7_75t_R _22245_ (.A1(_14015_),
    .A2(_04604_),
    .A3(_04606_),
    .B1(_04609_),
    .B2(_04610_),
    .B3(net315),
    .Y(_04611_));
 NAND2x1_ASAP7_75t_R _22246_ (.A(net412),
    .B(_01022_),
    .Y(_04612_));
 OA211x2_ASAP7_75t_R _22247_ (.A1(net412),
    .A2(_04521_),
    .B(_04612_),
    .C(net319),
    .Y(_04613_));
 NAND2x1_ASAP7_75t_R _22248_ (.A(net412),
    .B(_01021_),
    .Y(_04614_));
 OA211x2_ASAP7_75t_R _22249_ (.A1(net412),
    .A2(_04524_),
    .B(_04614_),
    .C(net426),
    .Y(_04615_));
 OR3x1_ASAP7_75t_R _22250_ (.A(net321),
    .B(_04613_),
    .C(_04615_),
    .Y(_04616_));
 NAND2x1_ASAP7_75t_R _22251_ (.A(net410),
    .B(_01026_),
    .Y(_04617_));
 OA211x2_ASAP7_75t_R _22252_ (.A1(net410),
    .A2(_04536_),
    .B(_04617_),
    .C(_13649_),
    .Y(_04618_));
 NAND2x1_ASAP7_75t_R _22253_ (.A(net412),
    .B(_01025_),
    .Y(_04619_));
 OA211x2_ASAP7_75t_R _22254_ (.A1(net412),
    .A2(_04539_),
    .B(_04619_),
    .C(net426),
    .Y(_04620_));
 OR3x1_ASAP7_75t_R _22255_ (.A(net387),
    .B(_04618_),
    .C(_04620_),
    .Y(_04621_));
 AO21x1_ASAP7_75t_R _22256_ (.A1(_04616_),
    .A2(_04621_),
    .B(net382),
    .Y(_04622_));
 AO21x2_ASAP7_75t_R _22257_ (.A1(_04611_),
    .A2(_04622_),
    .B(_13626_),
    .Y(_04623_));
 OA21x2_ASAP7_75t_R _22258_ (.A1(net377),
    .A2(_04602_),
    .B(_04623_),
    .Y(_04624_));
 TAPCELL_ASAP7_75t_R TAP_1083 ();
 AOI22x1_ASAP7_75t_R _22260_ (.A1(_13775_),
    .A2(_01045_),
    .B1(_02210_),
    .B2(_13778_),
    .Y(_04626_));
 OA211x2_ASAP7_75t_R _22261_ (.A1(_00284_),
    .A2(_04624_),
    .B(_04626_),
    .C(_13986_),
    .Y(_04627_));
 AO21x1_ASAP7_75t_R _22262_ (.A1(_13772_),
    .A2(_04576_),
    .B(_04627_),
    .Y(_04628_));
 AND2x2_ASAP7_75t_R _22263_ (.A(_13817_),
    .B(_04628_),
    .Y(_04629_));
 AOI21x1_ASAP7_75t_R _22264_ (.A1(net309),
    .A2(_04579_),
    .B(_04629_),
    .Y(_17795_));
 INVx1_ASAP7_75t_R _22265_ (.A(_17795_),
    .Y(_16754_));
 INVx1_ASAP7_75t_R _22266_ (.A(_00218_),
    .Y(\cs_registers_i.pc_id_i[23] ));
 OA211x2_ASAP7_75t_R _22267_ (.A1(net377),
    .A2(_04602_),
    .B(_04623_),
    .C(_13810_),
    .Y(_04630_));
 OAI22x1_ASAP7_75t_R _22268_ (.A1(_01618_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00218_),
    .Y(_04631_));
 OR2x2_ASAP7_75t_R _22269_ (.A(_04630_),
    .B(_04631_),
    .Y(_04632_));
 TAPCELL_ASAP7_75t_R TAP_1082 ();
 INVx2_ASAP7_75t_R _22271_ (.A(_04632_),
    .Y(_18440_));
 OA21x2_ASAP7_75t_R _22272_ (.A1(_01045_),
    .A2(_13815_),
    .B(_13817_),
    .Y(_04633_));
 AOI21x1_ASAP7_75t_R _22273_ (.A1(net309),
    .A2(_18440_),
    .B(_04633_),
    .Y(_17794_));
 INVx1_ASAP7_75t_R _22274_ (.A(_17794_),
    .Y(_16753_));
 OR4x1_ASAP7_75t_R _22275_ (.A(_00947_),
    .B(_00915_),
    .C(_01012_),
    .D(_00980_),
    .Y(_04634_));
 OA21x2_ASAP7_75t_R _22276_ (.A1(_00947_),
    .A2(_00948_),
    .B(_02277_),
    .Y(_04635_));
 OA21x2_ASAP7_75t_R _22277_ (.A1(_00980_),
    .A2(_04635_),
    .B(_01013_),
    .Y(_04636_));
 OA21x2_ASAP7_75t_R _22278_ (.A1(_01012_),
    .A2(_04636_),
    .B(_02278_),
    .Y(_04637_));
 OA21x2_ASAP7_75t_R _22279_ (.A1(_16747_),
    .A2(_04634_),
    .B(_04637_),
    .Y(_16752_));
 AND2x2_ASAP7_75t_R _22280_ (.A(net342),
    .B(_01685_),
    .Y(_04638_));
 AO21x1_ASAP7_75t_R _22281_ (.A1(net326),
    .A2(_01048_),
    .B(_04638_),
    .Y(_04639_));
 OAI22x1_ASAP7_75t_R _22282_ (.A1(_01047_),
    .A2(net311),
    .B1(_04639_),
    .B2(net376),
    .Y(_04640_));
 INVx1_ASAP7_75t_R _22283_ (.A(_01056_),
    .Y(_04641_));
 NAND2x1_ASAP7_75t_R _22284_ (.A(net345),
    .B(_01054_),
    .Y(_04642_));
 OA211x2_ASAP7_75t_R _22285_ (.A1(net345),
    .A2(_04641_),
    .B(_04642_),
    .C(_13376_),
    .Y(_04643_));
 INVx1_ASAP7_75t_R _22286_ (.A(_01055_),
    .Y(_04644_));
 NAND2x1_ASAP7_75t_R _22287_ (.A(net345),
    .B(_01053_),
    .Y(_04645_));
 OA211x2_ASAP7_75t_R _22288_ (.A1(net345),
    .A2(_04644_),
    .B(_04645_),
    .C(net376),
    .Y(_04646_));
 OR3x1_ASAP7_75t_R _22289_ (.A(net332),
    .B(_04643_),
    .C(_04646_),
    .Y(_04647_));
 OA211x2_ASAP7_75t_R _22290_ (.A1(_13373_),
    .A2(_04640_),
    .B(_04647_),
    .C(net338),
    .Y(_04648_));
 INVx1_ASAP7_75t_R _22291_ (.A(_01052_),
    .Y(_04649_));
 NAND2x1_ASAP7_75t_R _22292_ (.A(net345),
    .B(_01050_),
    .Y(_04650_));
 OA211x2_ASAP7_75t_R _22293_ (.A1(net345),
    .A2(_04649_),
    .B(_04650_),
    .C(_13376_),
    .Y(_04651_));
 INVx1_ASAP7_75t_R _22294_ (.A(_01051_),
    .Y(_04652_));
 NAND2x1_ASAP7_75t_R _22295_ (.A(net345),
    .B(_01049_),
    .Y(_04653_));
 OA211x2_ASAP7_75t_R _22296_ (.A1(net345),
    .A2(_04652_),
    .B(_04653_),
    .C(net376),
    .Y(_04654_));
 OR3x1_ASAP7_75t_R _22297_ (.A(_13373_),
    .B(_04651_),
    .C(_04654_),
    .Y(_04655_));
 INVx1_ASAP7_75t_R _22298_ (.A(_01060_),
    .Y(_04656_));
 NAND2x1_ASAP7_75t_R _22299_ (.A(net343),
    .B(_01058_),
    .Y(_04657_));
 OA211x2_ASAP7_75t_R _22300_ (.A1(net343),
    .A2(_04656_),
    .B(_04657_),
    .C(_13376_),
    .Y(_04658_));
 INVx1_ASAP7_75t_R _22301_ (.A(_01059_),
    .Y(_04659_));
 NAND2x1_ASAP7_75t_R _22302_ (.A(net343),
    .B(_01057_),
    .Y(_04660_));
 OA211x2_ASAP7_75t_R _22303_ (.A1(net343),
    .A2(_04659_),
    .B(_04660_),
    .C(net2314),
    .Y(_04661_));
 OR3x1_ASAP7_75t_R _22304_ (.A(_00245_),
    .B(_04658_),
    .C(_04661_),
    .Y(_04662_));
 AND3x1_ASAP7_75t_R _22305_ (.A(_13350_),
    .B(_04655_),
    .C(_04662_),
    .Y(_04663_));
 OR3x4_ASAP7_75t_R _22306_ (.A(_13355_),
    .B(_04648_),
    .C(_04663_),
    .Y(_04664_));
 TAPCELL_ASAP7_75t_R TAP_1081 ();
 INVx1_ASAP7_75t_R _22308_ (.A(_01068_),
    .Y(_04666_));
 NAND2x1_ASAP7_75t_R _22309_ (.A(net340),
    .B(_01066_),
    .Y(_04667_));
 OA211x2_ASAP7_75t_R _22310_ (.A1(net340),
    .A2(_04666_),
    .B(_04667_),
    .C(net323),
    .Y(_04668_));
 INVx1_ASAP7_75t_R _22311_ (.A(_01067_),
    .Y(_04669_));
 NAND2x1_ASAP7_75t_R _22312_ (.A(net340),
    .B(_01065_),
    .Y(_04670_));
 OA211x2_ASAP7_75t_R _22313_ (.A1(net340),
    .A2(_04669_),
    .B(_04670_),
    .C(net370),
    .Y(_04671_));
 OR3x1_ASAP7_75t_R _22314_ (.A(net338),
    .B(_04668_),
    .C(_04671_),
    .Y(_04672_));
 INVx1_ASAP7_75t_R _22315_ (.A(_01064_),
    .Y(_04673_));
 NAND2x1_ASAP7_75t_R _22316_ (.A(net340),
    .B(_01062_),
    .Y(_04674_));
 OA211x2_ASAP7_75t_R _22317_ (.A1(net340),
    .A2(_04673_),
    .B(_04674_),
    .C(net323),
    .Y(_04675_));
 INVx1_ASAP7_75t_R _22318_ (.A(_01063_),
    .Y(_04676_));
 NAND2x1_ASAP7_75t_R _22319_ (.A(net340),
    .B(_01061_),
    .Y(_04677_));
 OA211x2_ASAP7_75t_R _22320_ (.A1(net340),
    .A2(_04676_),
    .B(_04677_),
    .C(net370),
    .Y(_04678_));
 OR3x1_ASAP7_75t_R _22321_ (.A(_13350_),
    .B(_04675_),
    .C(_04678_),
    .Y(_04679_));
 AND3x1_ASAP7_75t_R _22322_ (.A(net332),
    .B(_04672_),
    .C(_04679_),
    .Y(_04680_));
 INVx1_ASAP7_75t_R _22323_ (.A(_01076_),
    .Y(_04681_));
 NAND2x1_ASAP7_75t_R _22324_ (.A(net343),
    .B(_01074_),
    .Y(_04682_));
 OA211x2_ASAP7_75t_R _22325_ (.A1(net343),
    .A2(_04681_),
    .B(_04682_),
    .C(_13376_),
    .Y(_04683_));
 INVx1_ASAP7_75t_R _22326_ (.A(_01075_),
    .Y(_04684_));
 NAND2x1_ASAP7_75t_R _22327_ (.A(net343),
    .B(_01073_),
    .Y(_04685_));
 OA211x2_ASAP7_75t_R _22328_ (.A1(net343),
    .A2(_04684_),
    .B(_04685_),
    .C(net2314),
    .Y(_04686_));
 OR3x1_ASAP7_75t_R _22329_ (.A(net338),
    .B(_04683_),
    .C(_04686_),
    .Y(_04687_));
 INVx1_ASAP7_75t_R _22330_ (.A(_01072_),
    .Y(_04688_));
 NAND2x1_ASAP7_75t_R _22331_ (.A(net343),
    .B(_01070_),
    .Y(_04689_));
 OA211x2_ASAP7_75t_R _22332_ (.A1(net343),
    .A2(_04688_),
    .B(_04689_),
    .C(_13376_),
    .Y(_04690_));
 INVx1_ASAP7_75t_R _22333_ (.A(_01071_),
    .Y(_04691_));
 NAND2x1_ASAP7_75t_R _22334_ (.A(net343),
    .B(_01069_),
    .Y(_04692_));
 OA211x2_ASAP7_75t_R _22335_ (.A1(net343),
    .A2(_04691_),
    .B(_04692_),
    .C(net2314),
    .Y(_04693_));
 OR3x1_ASAP7_75t_R _22336_ (.A(_13350_),
    .B(_04690_),
    .C(_04693_),
    .Y(_04694_));
 AND3x2_ASAP7_75t_R _22337_ (.A(_13373_),
    .B(_04687_),
    .C(_04694_),
    .Y(_04695_));
 OR3x4_ASAP7_75t_R _22338_ (.A(net328),
    .B(_04680_),
    .C(_04695_),
    .Y(_04696_));
 AND2x4_ASAP7_75t_R _22339_ (.A(_04664_),
    .B(_04696_),
    .Y(_04697_));
 INVx1_ASAP7_75t_R _22340_ (.A(_04697_),
    .Y(_04698_));
 OA21x2_ASAP7_75t_R _22341_ (.A1(_00244_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_04699_));
 AO21x2_ASAP7_75t_R _22342_ (.A1(_13474_),
    .A2(_04698_),
    .B(_04699_),
    .Y(_04700_));
 TAPCELL_ASAP7_75t_R TAP_1080 ();
 INVx1_ASAP7_75t_R _22344_ (.A(_04700_),
    .Y(_18445_));
 NAND2x1_ASAP7_75t_R _22345_ (.A(net393),
    .B(_01061_),
    .Y(_04701_));
 OA211x2_ASAP7_75t_R _22346_ (.A1(net393),
    .A2(_04676_),
    .B(_04701_),
    .C(net387),
    .Y(_04702_));
 NAND2x1_ASAP7_75t_R _22347_ (.A(net393),
    .B(_01065_),
    .Y(_04703_));
 OA211x2_ASAP7_75t_R _22348_ (.A1(net393),
    .A2(_04669_),
    .B(_04703_),
    .C(_13630_),
    .Y(_04704_));
 OR3x1_ASAP7_75t_R _22349_ (.A(_13649_),
    .B(_04702_),
    .C(_04704_),
    .Y(_04705_));
 NAND2x1_ASAP7_75t_R _22350_ (.A(net393),
    .B(_01062_),
    .Y(_04706_));
 OA211x2_ASAP7_75t_R _22351_ (.A1(net393),
    .A2(_04673_),
    .B(_04706_),
    .C(net387),
    .Y(_04707_));
 NAND2x1_ASAP7_75t_R _22352_ (.A(net393),
    .B(_01066_),
    .Y(_04708_));
 OA211x2_ASAP7_75t_R _22353_ (.A1(net393),
    .A2(_04666_),
    .B(_04708_),
    .C(net321),
    .Y(_04709_));
 OR3x1_ASAP7_75t_R _22354_ (.A(net426),
    .B(_04707_),
    .C(_04709_),
    .Y(_04710_));
 AND3x1_ASAP7_75t_R _22355_ (.A(net382),
    .B(_04705_),
    .C(_04710_),
    .Y(_04711_));
 NAND2x1_ASAP7_75t_R _22356_ (.A(net390),
    .B(_01069_),
    .Y(_04712_));
 OA211x2_ASAP7_75t_R _22357_ (.A1(net390),
    .A2(_04691_),
    .B(_04712_),
    .C(net388),
    .Y(_04713_));
 NAND2x1_ASAP7_75t_R _22358_ (.A(net390),
    .B(_01073_),
    .Y(_04714_));
 OA211x2_ASAP7_75t_R _22359_ (.A1(net390),
    .A2(_04684_),
    .B(_04714_),
    .C(_13630_),
    .Y(_04715_));
 OR3x1_ASAP7_75t_R _22360_ (.A(_13649_),
    .B(_04713_),
    .C(_04715_),
    .Y(_04716_));
 NAND2x1_ASAP7_75t_R _22361_ (.A(net391),
    .B(_01070_),
    .Y(_04717_));
 OA211x2_ASAP7_75t_R _22362_ (.A1(net391),
    .A2(_04688_),
    .B(_04717_),
    .C(net388),
    .Y(_04718_));
 NAND2x1_ASAP7_75t_R _22363_ (.A(net390),
    .B(_01074_),
    .Y(_04719_));
 OA211x2_ASAP7_75t_R _22364_ (.A1(net390),
    .A2(_04681_),
    .B(_04719_),
    .C(_13630_),
    .Y(_04720_));
 OR3x1_ASAP7_75t_R _22365_ (.A(net419),
    .B(_04718_),
    .C(_04720_),
    .Y(_04721_));
 AND3x2_ASAP7_75t_R _22366_ (.A(_13636_),
    .B(_04716_),
    .C(_04721_),
    .Y(_04722_));
 OR2x2_ASAP7_75t_R _22367_ (.A(_04711_),
    .B(_04722_),
    .Y(_04723_));
 NAND2x1_ASAP7_75t_R _22368_ (.A(net391),
    .B(_01050_),
    .Y(_04724_));
 OA211x2_ASAP7_75t_R _22369_ (.A1(net391),
    .A2(_04649_),
    .B(_04724_),
    .C(net319),
    .Y(_04725_));
 NAND2x1_ASAP7_75t_R _22370_ (.A(net391),
    .B(_01049_),
    .Y(_04726_));
 OA211x2_ASAP7_75t_R _22371_ (.A1(net391),
    .A2(_04652_),
    .B(_04726_),
    .C(net427),
    .Y(_04727_));
 INVx1_ASAP7_75t_R _22372_ (.A(_01048_),
    .Y(_04728_));
 NAND2x1_ASAP7_75t_R _22373_ (.A(net389),
    .B(_01685_),
    .Y(_04729_));
 OA211x2_ASAP7_75t_R _22374_ (.A1(net389),
    .A2(_04728_),
    .B(_04729_),
    .C(net319),
    .Y(_04730_));
 NOR2x1_ASAP7_75t_R _22375_ (.A(_01047_),
    .B(net2290),
    .Y(_04731_));
 OA33x2_ASAP7_75t_R _22376_ (.A1(_14015_),
    .A2(_04725_),
    .A3(_04727_),
    .B1(_04730_),
    .B2(_04731_),
    .B3(net315),
    .Y(_04732_));
 NAND2x1_ASAP7_75t_R _22377_ (.A(net391),
    .B(_01054_),
    .Y(_04733_));
 OA211x2_ASAP7_75t_R _22378_ (.A1(net391),
    .A2(_04641_),
    .B(_04733_),
    .C(_13649_),
    .Y(_04734_));
 NAND2x1_ASAP7_75t_R _22379_ (.A(net391),
    .B(_01053_),
    .Y(_04735_));
 OA211x2_ASAP7_75t_R _22380_ (.A1(net391),
    .A2(_04644_),
    .B(_04735_),
    .C(net427),
    .Y(_04736_));
 OR3x1_ASAP7_75t_R _22381_ (.A(_13630_),
    .B(_04734_),
    .C(_04736_),
    .Y(_04737_));
 NAND2x1_ASAP7_75t_R _22382_ (.A(net390),
    .B(_01058_),
    .Y(_04738_));
 OA211x2_ASAP7_75t_R _22383_ (.A1(net390),
    .A2(_04656_),
    .B(_04738_),
    .C(_13649_),
    .Y(_04739_));
 NAND2x1_ASAP7_75t_R _22384_ (.A(net390),
    .B(_01057_),
    .Y(_04740_));
 OA211x2_ASAP7_75t_R _22385_ (.A1(net390),
    .A2(_04659_),
    .B(_04740_),
    .C(net419),
    .Y(_04741_));
 OR3x1_ASAP7_75t_R _22386_ (.A(net388),
    .B(_04739_),
    .C(_04741_),
    .Y(_04742_));
 AO21x1_ASAP7_75t_R _22387_ (.A1(_04737_),
    .A2(_04742_),
    .B(net381),
    .Y(_04743_));
 AO21x2_ASAP7_75t_R _22388_ (.A1(_04732_),
    .A2(_04743_),
    .B(_13626_),
    .Y(_04744_));
 OA211x2_ASAP7_75t_R _22389_ (.A1(net378),
    .A2(_04723_),
    .B(_04744_),
    .C(_13810_),
    .Y(_04745_));
 OAI22x1_ASAP7_75t_R _22390_ (.A1(_01617_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00220_),
    .Y(_04746_));
 NOR2x2_ASAP7_75t_R _22391_ (.A(_04745_),
    .B(_04746_),
    .Y(_18444_));
 XOR2x2_ASAP7_75t_R _22392_ (.A(_01078_),
    .B(_02230_),
    .Y(_04747_));
 INVx5_ASAP7_75t_R _22393_ (.A(_04747_),
    .Y(net165));
 INVx1_ASAP7_75t_R _22394_ (.A(_01080_),
    .Y(_04748_));
 INVx1_ASAP7_75t_R _22395_ (.A(_01081_),
    .Y(_04749_));
 NAND2x1_ASAP7_75t_R _22396_ (.A(net357),
    .B(_01684_),
    .Y(_04750_));
 OA211x2_ASAP7_75t_R _22397_ (.A1(net357),
    .A2(_04749_),
    .B(_04750_),
    .C(net324),
    .Y(_04751_));
 AO21x1_ASAP7_75t_R _22398_ (.A1(_04748_),
    .A2(net2228),
    .B(_04751_),
    .Y(_04752_));
 INVx1_ASAP7_75t_R _22399_ (.A(_01089_),
    .Y(_04753_));
 NAND2x1_ASAP7_75t_R _22400_ (.A(net357),
    .B(_01087_),
    .Y(_04754_));
 OA211x2_ASAP7_75t_R _22401_ (.A1(net357),
    .A2(_04753_),
    .B(_04754_),
    .C(net324),
    .Y(_04755_));
 INVx1_ASAP7_75t_R _22402_ (.A(_01088_),
    .Y(_04756_));
 NAND2x1_ASAP7_75t_R _22403_ (.A(net357),
    .B(_01086_),
    .Y(_04757_));
 OA211x2_ASAP7_75t_R _22404_ (.A1(net357),
    .A2(_04756_),
    .B(_04757_),
    .C(net372),
    .Y(_04758_));
 OR3x1_ASAP7_75t_R _22405_ (.A(net330),
    .B(_04755_),
    .C(_04758_),
    .Y(_04759_));
 OA211x2_ASAP7_75t_R _22406_ (.A1(_13373_),
    .A2(_04752_),
    .B(_04759_),
    .C(net334),
    .Y(_04760_));
 INVx1_ASAP7_75t_R _22407_ (.A(_01085_),
    .Y(_04761_));
 NAND2x1_ASAP7_75t_R _22408_ (.A(net359),
    .B(_01083_),
    .Y(_04762_));
 OA211x2_ASAP7_75t_R _22409_ (.A1(net2332),
    .A2(_04761_),
    .B(_04762_),
    .C(net324),
    .Y(_04763_));
 INVx1_ASAP7_75t_R _22410_ (.A(_01084_),
    .Y(_04764_));
 NAND2x1_ASAP7_75t_R _22411_ (.A(net2332),
    .B(_01082_),
    .Y(_04765_));
 OA211x2_ASAP7_75t_R _22412_ (.A1(net2332),
    .A2(_04764_),
    .B(_04765_),
    .C(net372),
    .Y(_04766_));
 OR3x1_ASAP7_75t_R _22413_ (.A(_13373_),
    .B(_04763_),
    .C(_04766_),
    .Y(_04767_));
 INVx1_ASAP7_75t_R _22414_ (.A(_01093_),
    .Y(_04768_));
 NAND2x1_ASAP7_75t_R _22415_ (.A(net2280),
    .B(_01091_),
    .Y(_04769_));
 OA211x2_ASAP7_75t_R _22416_ (.A1(net2280),
    .A2(_04768_),
    .B(_04769_),
    .C(net324),
    .Y(_04770_));
 INVx1_ASAP7_75t_R _22417_ (.A(_01092_),
    .Y(_04771_));
 NAND2x1_ASAP7_75t_R _22418_ (.A(net357),
    .B(_01090_),
    .Y(_04772_));
 OA211x2_ASAP7_75t_R _22419_ (.A1(net357),
    .A2(_04771_),
    .B(_04772_),
    .C(net372),
    .Y(_04773_));
 OR3x1_ASAP7_75t_R _22420_ (.A(net330),
    .B(_04770_),
    .C(_04773_),
    .Y(_04774_));
 AND3x1_ASAP7_75t_R _22421_ (.A(_13350_),
    .B(_04767_),
    .C(_04774_),
    .Y(_04775_));
 OR3x1_ASAP7_75t_R _22422_ (.A(_13355_),
    .B(_04760_),
    .C(_04775_),
    .Y(_04776_));
 INVx1_ASAP7_75t_R _22423_ (.A(_01101_),
    .Y(_04777_));
 NAND2x1_ASAP7_75t_R _22424_ (.A(net2280),
    .B(_01099_),
    .Y(_04778_));
 OA211x2_ASAP7_75t_R _22425_ (.A1(net2280),
    .A2(_04777_),
    .B(_04778_),
    .C(net324),
    .Y(_04779_));
 INVx1_ASAP7_75t_R _22426_ (.A(_01100_),
    .Y(_04780_));
 NAND2x1_ASAP7_75t_R _22427_ (.A(net2280),
    .B(_01098_),
    .Y(_04781_));
 OA211x2_ASAP7_75t_R _22428_ (.A1(net2280),
    .A2(_04780_),
    .B(_04781_),
    .C(net371),
    .Y(_04782_));
 OR3x1_ASAP7_75t_R _22429_ (.A(net334),
    .B(_04779_),
    .C(_04782_),
    .Y(_04783_));
 INVx1_ASAP7_75t_R _22430_ (.A(_01097_),
    .Y(_04784_));
 NAND2x1_ASAP7_75t_R _22431_ (.A(net355),
    .B(_01095_),
    .Y(_04785_));
 OA211x2_ASAP7_75t_R _22432_ (.A1(net2331),
    .A2(_04784_),
    .B(_04785_),
    .C(net324),
    .Y(_04786_));
 INVx1_ASAP7_75t_R _22433_ (.A(_01096_),
    .Y(_04787_));
 NAND2x1_ASAP7_75t_R _22434_ (.A(net355),
    .B(_01094_),
    .Y(_04788_));
 OA211x2_ASAP7_75t_R _22435_ (.A1(net2331),
    .A2(_04787_),
    .B(_04788_),
    .C(net371),
    .Y(_04789_));
 OR3x1_ASAP7_75t_R _22436_ (.A(_13350_),
    .B(_04786_),
    .C(_04789_),
    .Y(_04790_));
 AND3x1_ASAP7_75t_R _22437_ (.A(net330),
    .B(_04783_),
    .C(_04790_),
    .Y(_04791_));
 INVx1_ASAP7_75t_R _22438_ (.A(_01105_),
    .Y(_04792_));
 NAND2x1_ASAP7_75t_R _22439_ (.A(net2284),
    .B(_01103_),
    .Y(_04793_));
 OA211x2_ASAP7_75t_R _22440_ (.A1(net2294),
    .A2(_04792_),
    .B(_04793_),
    .C(net324),
    .Y(_04794_));
 INVx1_ASAP7_75t_R _22441_ (.A(_01104_),
    .Y(_04795_));
 NAND2x1_ASAP7_75t_R _22442_ (.A(net355),
    .B(_01102_),
    .Y(_04796_));
 OA211x2_ASAP7_75t_R _22443_ (.A1(net2331),
    .A2(_04795_),
    .B(_04796_),
    .C(net371),
    .Y(_04797_));
 OR3x1_ASAP7_75t_R _22444_ (.A(_13350_),
    .B(_04794_),
    .C(_04797_),
    .Y(_04798_));
 INVx1_ASAP7_75t_R _22445_ (.A(_01109_),
    .Y(_04799_));
 NAND2x1_ASAP7_75t_R _22446_ (.A(net2373),
    .B(_01107_),
    .Y(_04800_));
 OA211x2_ASAP7_75t_R _22447_ (.A1(net2279),
    .A2(_04799_),
    .B(_04800_),
    .C(net324),
    .Y(_04801_));
 INVx1_ASAP7_75t_R _22448_ (.A(_01108_),
    .Y(_04802_));
 NAND2x1_ASAP7_75t_R _22449_ (.A(net2373),
    .B(_01106_),
    .Y(_04803_));
 OA211x2_ASAP7_75t_R _22450_ (.A1(net2279),
    .A2(_04802_),
    .B(_04803_),
    .C(net371),
    .Y(_04804_));
 OR3x1_ASAP7_75t_R _22451_ (.A(net334),
    .B(_04801_),
    .C(_04804_),
    .Y(_04805_));
 AND3x1_ASAP7_75t_R _22452_ (.A(_13373_),
    .B(_04798_),
    .C(_04805_),
    .Y(_04806_));
 OR3x2_ASAP7_75t_R _22453_ (.A(net327),
    .B(_04791_),
    .C(_04806_),
    .Y(_04807_));
 NAND2x2_ASAP7_75t_R _22454_ (.A(_04776_),
    .B(_04807_),
    .Y(_04808_));
 OA21x2_ASAP7_75t_R _22455_ (.A1(_01743_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_04809_));
 AO21x2_ASAP7_75t_R _22456_ (.A1(_13474_),
    .A2(_04808_),
    .B(_04809_),
    .Y(_04810_));
 TAPCELL_ASAP7_75t_R TAP_1079 ();
 INVx1_ASAP7_75t_R _22458_ (.A(_04810_),
    .Y(_18450_));
 INVx1_ASAP7_75t_R _22459_ (.A(_00221_),
    .Y(\cs_registers_i.pc_id_i[25] ));
 NAND2x1_ASAP7_75t_R _22460_ (.A(net400),
    .B(_01098_),
    .Y(_04811_));
 OA211x2_ASAP7_75t_R _22461_ (.A1(net400),
    .A2(_04780_),
    .B(_04811_),
    .C(net421),
    .Y(_04812_));
 NAND2x1_ASAP7_75t_R _22462_ (.A(net400),
    .B(_01099_),
    .Y(_04813_));
 OA211x2_ASAP7_75t_R _22463_ (.A1(net400),
    .A2(_04777_),
    .B(_04813_),
    .C(net317),
    .Y(_04814_));
 OR3x1_ASAP7_75t_R _22464_ (.A(net312),
    .B(_04812_),
    .C(_04814_),
    .Y(_04815_));
 NAND2x1_ASAP7_75t_R _22465_ (.A(net399),
    .B(_01094_),
    .Y(_04816_));
 OA211x2_ASAP7_75t_R _22466_ (.A1(net399),
    .A2(_04787_),
    .B(_04816_),
    .C(net421),
    .Y(_04817_));
 NAND2x1_ASAP7_75t_R _22467_ (.A(net399),
    .B(_01095_),
    .Y(_04818_));
 OA211x2_ASAP7_75t_R _22468_ (.A1(net399),
    .A2(_04784_),
    .B(_04818_),
    .C(net317),
    .Y(_04819_));
 OR3x1_ASAP7_75t_R _22469_ (.A(_14005_),
    .B(_04817_),
    .C(_04819_),
    .Y(_04820_));
 AND3x1_ASAP7_75t_R _22470_ (.A(_13626_),
    .B(_04815_),
    .C(_04820_),
    .Y(_04821_));
 NAND2x1_ASAP7_75t_R _22471_ (.A(net399),
    .B(_01103_),
    .Y(_04822_));
 OA211x2_ASAP7_75t_R _22472_ (.A1(net399),
    .A2(_04792_),
    .B(_04822_),
    .C(net317),
    .Y(_04823_));
 NAND2x1_ASAP7_75t_R _22473_ (.A(net399),
    .B(_01102_),
    .Y(_04824_));
 OA211x2_ASAP7_75t_R _22474_ (.A1(net399),
    .A2(_04795_),
    .B(_04824_),
    .C(net421),
    .Y(_04825_));
 OR3x1_ASAP7_75t_R _22475_ (.A(net321),
    .B(_04823_),
    .C(_04825_),
    .Y(_04826_));
 NAND2x1_ASAP7_75t_R _22476_ (.A(net399),
    .B(_01107_),
    .Y(_04827_));
 OA211x2_ASAP7_75t_R _22477_ (.A1(net399),
    .A2(_04799_),
    .B(_04827_),
    .C(net317),
    .Y(_04828_));
 NAND2x1_ASAP7_75t_R _22478_ (.A(net399),
    .B(_01106_),
    .Y(_04829_));
 OA211x2_ASAP7_75t_R _22479_ (.A1(net399),
    .A2(_04802_),
    .B(_04829_),
    .C(net421),
    .Y(_04830_));
 OR3x1_ASAP7_75t_R _22480_ (.A(net383),
    .B(_04828_),
    .C(_04830_),
    .Y(_04831_));
 AND2x2_ASAP7_75t_R _22481_ (.A(_04826_),
    .B(_04831_),
    .Y(_04832_));
 NAND2x1_ASAP7_75t_R _22482_ (.A(net400),
    .B(_01083_),
    .Y(_04833_));
 OA211x2_ASAP7_75t_R _22483_ (.A1(net400),
    .A2(_04761_),
    .B(_04833_),
    .C(net317),
    .Y(_04834_));
 NAND2x1_ASAP7_75t_R _22484_ (.A(net400),
    .B(_01082_),
    .Y(_04835_));
 OA211x2_ASAP7_75t_R _22485_ (.A1(net400),
    .A2(_04764_),
    .B(_04835_),
    .C(net422),
    .Y(_04836_));
 OR3x1_ASAP7_75t_R _22486_ (.A(net312),
    .B(_04834_),
    .C(_04836_),
    .Y(_04837_));
 NAND2x1_ASAP7_75t_R _22487_ (.A(net399),
    .B(_01684_),
    .Y(_04838_));
 OA211x2_ASAP7_75t_R _22488_ (.A1(net399),
    .A2(_04749_),
    .B(_04838_),
    .C(net317),
    .Y(_04839_));
 AND3x1_ASAP7_75t_R _22489_ (.A(net421),
    .B(net316),
    .C(_04748_),
    .Y(_04840_));
 OA31x2_ASAP7_75t_R _22490_ (.A1(_14005_),
    .A2(_04839_),
    .A3(_04840_),
    .B1(net377),
    .Y(_04841_));
 AO32x1_ASAP7_75t_R _22491_ (.A1(_13626_),
    .A2(_04815_),
    .A3(_04820_),
    .B1(_04837_),
    .B2(_04841_),
    .Y(_04842_));
 NAND2x1_ASAP7_75t_R _22492_ (.A(net400),
    .B(_01091_),
    .Y(_04843_));
 OA211x2_ASAP7_75t_R _22493_ (.A1(net400),
    .A2(_04768_),
    .B(_04843_),
    .C(net317),
    .Y(_04844_));
 NAND2x1_ASAP7_75t_R _22494_ (.A(net400),
    .B(_01090_),
    .Y(_04845_));
 OA211x2_ASAP7_75t_R _22495_ (.A1(net400),
    .A2(_04771_),
    .B(_04845_),
    .C(net421),
    .Y(_04846_));
 OR3x1_ASAP7_75t_R _22496_ (.A(net383),
    .B(_04844_),
    .C(_04846_),
    .Y(_04847_));
 NAND2x1_ASAP7_75t_R _22497_ (.A(net400),
    .B(_01087_),
    .Y(_04848_));
 OA211x2_ASAP7_75t_R _22498_ (.A1(net400),
    .A2(_04753_),
    .B(_04848_),
    .C(net317),
    .Y(_04849_));
 NAND2x1_ASAP7_75t_R _22499_ (.A(net400),
    .B(_01086_),
    .Y(_04850_));
 OA211x2_ASAP7_75t_R _22500_ (.A1(net400),
    .A2(_04756_),
    .B(_04850_),
    .C(net421),
    .Y(_04851_));
 OR3x1_ASAP7_75t_R _22501_ (.A(net320),
    .B(_04849_),
    .C(_04851_),
    .Y(_04852_));
 AND4x1_ASAP7_75t_R _22502_ (.A(_04837_),
    .B(_04841_),
    .C(_04847_),
    .D(_04852_),
    .Y(_04853_));
 AO221x2_ASAP7_75t_R _22503_ (.A1(_04821_),
    .A2(_04832_),
    .B1(_04842_),
    .B2(net379),
    .C(_04853_),
    .Y(_04854_));
 OA211x2_ASAP7_75t_R _22504_ (.A1(_13788_),
    .A2(_13806_),
    .B(_00221_),
    .C(_13807_),
    .Y(_04855_));
 OAI22x1_ASAP7_75t_R _22505_ (.A1(_01616_),
    .A2(_13807_),
    .B1(_14988_),
    .B2(_04855_),
    .Y(_04856_));
 OA21x2_ASAP7_75t_R _22506_ (.A1(_15112_),
    .A2(_04854_),
    .B(_04856_),
    .Y(_04857_));
 TAPCELL_ASAP7_75t_R TAP_1078 ();
 INVx2_ASAP7_75t_R _22508_ (.A(_04857_),
    .Y(_18449_));
 INVx1_ASAP7_75t_R _22509_ (.A(_01122_),
    .Y(_04858_));
 NOR2x1_ASAP7_75t_R _22510_ (.A(net349),
    .B(_01124_),
    .Y(_04859_));
 AO21x1_ASAP7_75t_R _22511_ (.A1(net349),
    .A2(_04858_),
    .B(_04859_),
    .Y(_04860_));
 INVx1_ASAP7_75t_R _22512_ (.A(_01125_),
    .Y(_04861_));
 NAND2x1_ASAP7_75t_R _22513_ (.A(net349),
    .B(_01123_),
    .Y(_04862_));
 OA211x2_ASAP7_75t_R _22514_ (.A1(net349),
    .A2(_04861_),
    .B(_04862_),
    .C(net325),
    .Y(_04863_));
 AO21x1_ASAP7_75t_R _22515_ (.A1(net369),
    .A2(_04860_),
    .B(_04863_),
    .Y(_04864_));
 INVx1_ASAP7_75t_R _22516_ (.A(_01117_),
    .Y(_04865_));
 NAND2x1_ASAP7_75t_R _22517_ (.A(net349),
    .B(_01115_),
    .Y(_04866_));
 OA211x2_ASAP7_75t_R _22518_ (.A1(net349),
    .A2(_04865_),
    .B(_04866_),
    .C(net325),
    .Y(_04867_));
 INVx1_ASAP7_75t_R _22519_ (.A(_01116_),
    .Y(_04868_));
 NAND2x1_ASAP7_75t_R _22520_ (.A(net349),
    .B(_01114_),
    .Y(_04869_));
 OA211x2_ASAP7_75t_R _22521_ (.A1(net349),
    .A2(_04868_),
    .B(_04869_),
    .C(net369),
    .Y(_04870_));
 OR3x1_ASAP7_75t_R _22522_ (.A(_13373_),
    .B(_04867_),
    .C(_04870_),
    .Y(_04871_));
 OA21x2_ASAP7_75t_R _22523_ (.A1(net331),
    .A2(_04864_),
    .B(_04871_),
    .Y(_04872_));
 AND2x2_ASAP7_75t_R _22524_ (.A(net351),
    .B(_01683_),
    .Y(_04873_));
 AO21x1_ASAP7_75t_R _22525_ (.A1(net2260),
    .A2(_01113_),
    .B(_04873_),
    .Y(_04874_));
 OAI22x1_ASAP7_75t_R _22526_ (.A1(_01112_),
    .A2(net311),
    .B1(_04874_),
    .B2(net369),
    .Y(_04875_));
 INVx1_ASAP7_75t_R _22527_ (.A(_01121_),
    .Y(_04876_));
 NAND2x1_ASAP7_75t_R _22528_ (.A(net351),
    .B(_01119_),
    .Y(_04877_));
 OA211x2_ASAP7_75t_R _22529_ (.A1(net351),
    .A2(_04876_),
    .B(_04877_),
    .C(net325),
    .Y(_04878_));
 INVx1_ASAP7_75t_R _22530_ (.A(_01120_),
    .Y(_04879_));
 NAND2x1_ASAP7_75t_R _22531_ (.A(net351),
    .B(_01118_),
    .Y(_04880_));
 OA211x2_ASAP7_75t_R _22532_ (.A1(net351),
    .A2(_04879_),
    .B(_04880_),
    .C(net369),
    .Y(_04881_));
 OR3x1_ASAP7_75t_R _22533_ (.A(net330),
    .B(_04878_),
    .C(_04881_),
    .Y(_04882_));
 OA211x2_ASAP7_75t_R _22534_ (.A1(_13373_),
    .A2(_04875_),
    .B(_04882_),
    .C(net335),
    .Y(_04883_));
 AO21x1_ASAP7_75t_R _22535_ (.A1(_13350_),
    .A2(_04872_),
    .B(_04883_),
    .Y(_04884_));
 INVx1_ASAP7_75t_R _22536_ (.A(_01129_),
    .Y(_04885_));
 NAND2x1_ASAP7_75t_R _22537_ (.A(net349),
    .B(_01127_),
    .Y(_04886_));
 OA211x2_ASAP7_75t_R _22538_ (.A1(net349),
    .A2(_04885_),
    .B(_04886_),
    .C(net325),
    .Y(_04887_));
 INVx1_ASAP7_75t_R _22539_ (.A(_01128_),
    .Y(_04888_));
 NAND2x1_ASAP7_75t_R _22540_ (.A(net349),
    .B(_01126_),
    .Y(_04889_));
 OA211x2_ASAP7_75t_R _22541_ (.A1(net349),
    .A2(_04888_),
    .B(_04889_),
    .C(net369),
    .Y(_04890_));
 OR3x1_ASAP7_75t_R _22542_ (.A(_13350_),
    .B(_04887_),
    .C(_04890_),
    .Y(_04891_));
 INVx1_ASAP7_75t_R _22543_ (.A(_01133_),
    .Y(_04892_));
 NAND2x1_ASAP7_75t_R _22544_ (.A(net349),
    .B(_01131_),
    .Y(_04893_));
 OA211x2_ASAP7_75t_R _22545_ (.A1(net349),
    .A2(_04892_),
    .B(_04893_),
    .C(net325),
    .Y(_04894_));
 INVx1_ASAP7_75t_R _22546_ (.A(_01132_),
    .Y(_04895_));
 NAND2x1_ASAP7_75t_R _22547_ (.A(net349),
    .B(_01130_),
    .Y(_04896_));
 OA211x2_ASAP7_75t_R _22548_ (.A1(net349),
    .A2(_04895_),
    .B(_04896_),
    .C(net369),
    .Y(_04897_));
 OR3x1_ASAP7_75t_R _22549_ (.A(net335),
    .B(_04894_),
    .C(_04897_),
    .Y(_04898_));
 AND3x1_ASAP7_75t_R _22550_ (.A(net331),
    .B(_04891_),
    .C(_04898_),
    .Y(_04899_));
 INVx1_ASAP7_75t_R _22551_ (.A(_01137_),
    .Y(_04900_));
 NAND2x1_ASAP7_75t_R _22552_ (.A(net351),
    .B(_01135_),
    .Y(_04901_));
 OA211x2_ASAP7_75t_R _22553_ (.A1(net351),
    .A2(_04900_),
    .B(_04901_),
    .C(net325),
    .Y(_04902_));
 INVx1_ASAP7_75t_R _22554_ (.A(_01136_),
    .Y(_04903_));
 NAND2x1_ASAP7_75t_R _22555_ (.A(net351),
    .B(_01134_),
    .Y(_04904_));
 OA211x2_ASAP7_75t_R _22556_ (.A1(net351),
    .A2(_04903_),
    .B(_04904_),
    .C(net369),
    .Y(_04905_));
 OR3x1_ASAP7_75t_R _22557_ (.A(_13350_),
    .B(_04902_),
    .C(_04905_),
    .Y(_04906_));
 INVx1_ASAP7_75t_R _22558_ (.A(_01141_),
    .Y(_04907_));
 NAND2x1_ASAP7_75t_R _22559_ (.A(net350),
    .B(_01139_),
    .Y(_04908_));
 OA211x2_ASAP7_75t_R _22560_ (.A1(net350),
    .A2(_04907_),
    .B(_04908_),
    .C(net325),
    .Y(_04909_));
 INVx1_ASAP7_75t_R _22561_ (.A(_01140_),
    .Y(_04910_));
 NAND2x1_ASAP7_75t_R _22562_ (.A(net350),
    .B(_01138_),
    .Y(_04911_));
 OA211x2_ASAP7_75t_R _22563_ (.A1(net350),
    .A2(_04910_),
    .B(_04911_),
    .C(net373),
    .Y(_04912_));
 OR3x1_ASAP7_75t_R _22564_ (.A(net335),
    .B(_04909_),
    .C(_04912_),
    .Y(_04913_));
 AND3x1_ASAP7_75t_R _22565_ (.A(_13373_),
    .B(_04906_),
    .C(_04913_),
    .Y(_04914_));
 OR3x1_ASAP7_75t_R _22566_ (.A(net327),
    .B(_04899_),
    .C(_04914_),
    .Y(_04915_));
 OA21x2_ASAP7_75t_R _22567_ (.A1(_13355_),
    .A2(_04884_),
    .B(_04915_),
    .Y(_04916_));
 TAPCELL_ASAP7_75t_R TAP_1077 ();
 OAI21x1_ASAP7_75t_R _22569_ (.A1(_00283_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_04918_));
 OA21x2_ASAP7_75t_R _22570_ (.A1(_13521_),
    .A2(_04916_),
    .B(_04918_),
    .Y(_04919_));
 TAPCELL_ASAP7_75t_R TAP_1076 ();
 AND2x2_ASAP7_75t_R _22572_ (.A(net396),
    .B(_01683_),
    .Y(_04920_));
 AO21x1_ASAP7_75t_R _22573_ (.A1(net316),
    .A2(_01113_),
    .B(_04920_),
    .Y(_04921_));
 OAI22x1_ASAP7_75t_R _22574_ (.A1(_01112_),
    .A2(net2289),
    .B1(_04921_),
    .B2(net423),
    .Y(_04922_));
 NAND2x1_ASAP7_75t_R _22575_ (.A(net396),
    .B(_01127_),
    .Y(_04923_));
 OA211x2_ASAP7_75t_R _22576_ (.A1(net396),
    .A2(_04885_),
    .B(_04923_),
    .C(_13649_),
    .Y(_04924_));
 NAND2x1_ASAP7_75t_R _22577_ (.A(net396),
    .B(_01126_),
    .Y(_04925_));
 OA211x2_ASAP7_75t_R _22578_ (.A1(net396),
    .A2(_04888_),
    .B(_04925_),
    .C(net423),
    .Y(_04926_));
 OR3x1_ASAP7_75t_R _22579_ (.A(net378),
    .B(_04924_),
    .C(_04926_),
    .Y(_04927_));
 OA211x2_ASAP7_75t_R _22580_ (.A1(_13626_),
    .A2(_04922_),
    .B(_04927_),
    .C(net386),
    .Y(_04928_));
 NAND2x1_ASAP7_75t_R _22581_ (.A(net396),
    .B(_01115_),
    .Y(_04929_));
 OA211x2_ASAP7_75t_R _22582_ (.A1(net396),
    .A2(_04865_),
    .B(_04929_),
    .C(_13649_),
    .Y(_04930_));
 NAND2x1_ASAP7_75t_R _22583_ (.A(net396),
    .B(_01114_),
    .Y(_04931_));
 OA211x2_ASAP7_75t_R _22584_ (.A1(net396),
    .A2(_04868_),
    .B(_04931_),
    .C(net423),
    .Y(_04932_));
 OR3x1_ASAP7_75t_R _22585_ (.A(_13626_),
    .B(_04930_),
    .C(_04932_),
    .Y(_04933_));
 NAND2x1_ASAP7_75t_R _22586_ (.A(net396),
    .B(_01131_),
    .Y(_04934_));
 OA211x2_ASAP7_75t_R _22587_ (.A1(net396),
    .A2(_04892_),
    .B(_04934_),
    .C(_13649_),
    .Y(_04935_));
 NAND2x1_ASAP7_75t_R _22588_ (.A(net395),
    .B(_01130_),
    .Y(_04936_));
 OA211x2_ASAP7_75t_R _22589_ (.A1(net396),
    .A2(_04895_),
    .B(_04936_),
    .C(net423),
    .Y(_04937_));
 OR3x1_ASAP7_75t_R _22590_ (.A(net378),
    .B(_04935_),
    .C(_04937_),
    .Y(_04938_));
 AND3x1_ASAP7_75t_R _22591_ (.A(net321),
    .B(_04933_),
    .C(_04938_),
    .Y(_04939_));
 OR3x1_ASAP7_75t_R _22592_ (.A(_13636_),
    .B(_04928_),
    .C(_04939_),
    .Y(_04940_));
 NAND2x1_ASAP7_75t_R _22593_ (.A(net397),
    .B(_01135_),
    .Y(_04941_));
 OA211x2_ASAP7_75t_R _22594_ (.A1(net397),
    .A2(_04900_),
    .B(_04941_),
    .C(net318),
    .Y(_04942_));
 NAND2x1_ASAP7_75t_R _22595_ (.A(net397),
    .B(_01134_),
    .Y(_04943_));
 OA211x2_ASAP7_75t_R _22596_ (.A1(net397),
    .A2(_04903_),
    .B(_04943_),
    .C(net423),
    .Y(_04944_));
 OR3x1_ASAP7_75t_R _22597_ (.A(net320),
    .B(_04942_),
    .C(_04944_),
    .Y(_04945_));
 NAND2x1_ASAP7_75t_R _22598_ (.A(net396),
    .B(_01139_),
    .Y(_04946_));
 OA211x2_ASAP7_75t_R _22599_ (.A1(net396),
    .A2(_04907_),
    .B(_04946_),
    .C(net317),
    .Y(_04947_));
 NAND2x1_ASAP7_75t_R _22600_ (.A(net396),
    .B(_01138_),
    .Y(_04948_));
 OA211x2_ASAP7_75t_R _22601_ (.A1(net396),
    .A2(_04910_),
    .B(_04948_),
    .C(net423),
    .Y(_04949_));
 OR3x1_ASAP7_75t_R _22602_ (.A(net386),
    .B(_04947_),
    .C(_04949_),
    .Y(_04950_));
 AND3x1_ASAP7_75t_R _22603_ (.A(_13626_),
    .B(_04945_),
    .C(_04950_),
    .Y(_04951_));
 INVx1_ASAP7_75t_R _22604_ (.A(_01123_),
    .Y(_04952_));
 NAND2x1_ASAP7_75t_R _22605_ (.A(net386),
    .B(_01119_),
    .Y(_04953_));
 OA211x2_ASAP7_75t_R _22606_ (.A1(net386),
    .A2(_04952_),
    .B(_04953_),
    .C(net317),
    .Y(_04954_));
 NAND2x1_ASAP7_75t_R _22607_ (.A(net386),
    .B(_01118_),
    .Y(_04955_));
 OA211x2_ASAP7_75t_R _22608_ (.A1(net386),
    .A2(_04858_),
    .B(_04955_),
    .C(net423),
    .Y(_04956_));
 OR3x1_ASAP7_75t_R _22609_ (.A(net316),
    .B(_04954_),
    .C(_04956_),
    .Y(_04957_));
 NAND2x1_ASAP7_75t_R _22610_ (.A(net423),
    .B(_01120_),
    .Y(_04958_));
 OA211x2_ASAP7_75t_R _22611_ (.A1(net423),
    .A2(_04876_),
    .B(_04958_),
    .C(net386),
    .Y(_04959_));
 NAND2x1_ASAP7_75t_R _22612_ (.A(net423),
    .B(_01124_),
    .Y(_04960_));
 OA211x2_ASAP7_75t_R _22613_ (.A1(net423),
    .A2(_04861_),
    .B(_04960_),
    .C(net320),
    .Y(_04961_));
 OR3x1_ASAP7_75t_R _22614_ (.A(net396),
    .B(_04959_),
    .C(_04961_),
    .Y(_04962_));
 AND3x1_ASAP7_75t_R _22615_ (.A(net378),
    .B(_04957_),
    .C(_04962_),
    .Y(_04963_));
 OR3x1_ASAP7_75t_R _22616_ (.A(net379),
    .B(_04951_),
    .C(_04963_),
    .Y(_04964_));
 AND2x6_ASAP7_75t_R _22617_ (.A(_04940_),
    .B(_04964_),
    .Y(_04965_));
 OAI22x1_ASAP7_75t_R _22618_ (.A1(_01615_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00223_),
    .Y(_04966_));
 AO21x2_ASAP7_75t_R _22619_ (.A1(_13810_),
    .A2(_04965_),
    .B(_04966_),
    .Y(_04967_));
 TAPCELL_ASAP7_75t_R TAP_1075 ();
 INVx2_ASAP7_75t_R _22621_ (.A(_04967_),
    .Y(_18455_));
 XNOR2x2_ASAP7_75t_R _22622_ (.A(_01145_),
    .B(_01143_),
    .Y(_04968_));
 INVx2_ASAP7_75t_R _22623_ (.A(_04968_),
    .Y(net167));
 AND2x2_ASAP7_75t_R _22624_ (.A(net352),
    .B(_01682_),
    .Y(_04969_));
 AO21x1_ASAP7_75t_R _22625_ (.A1(net2260),
    .A2(_01147_),
    .B(_04969_),
    .Y(_04970_));
 OAI22x1_ASAP7_75t_R _22626_ (.A1(_01146_),
    .A2(net311),
    .B1(_04970_),
    .B2(net375),
    .Y(_04971_));
 INVx1_ASAP7_75t_R _22627_ (.A(_01155_),
    .Y(_04972_));
 NAND2x1_ASAP7_75t_R _22628_ (.A(net348),
    .B(_01153_),
    .Y(_04973_));
 OA211x2_ASAP7_75t_R _22629_ (.A1(net348),
    .A2(_04972_),
    .B(_04973_),
    .C(net325),
    .Y(_04974_));
 INVx1_ASAP7_75t_R _22630_ (.A(_01154_),
    .Y(_04975_));
 NAND2x1_ASAP7_75t_R _22631_ (.A(net348),
    .B(_01152_),
    .Y(_04976_));
 OA211x2_ASAP7_75t_R _22632_ (.A1(net348),
    .A2(_04975_),
    .B(_04976_),
    .C(net375),
    .Y(_04977_));
 OR3x1_ASAP7_75t_R _22633_ (.A(net331),
    .B(_04974_),
    .C(_04977_),
    .Y(_04978_));
 OA211x2_ASAP7_75t_R _22634_ (.A1(_13373_),
    .A2(_04971_),
    .B(_04978_),
    .C(net335),
    .Y(_04979_));
 INVx1_ASAP7_75t_R _22635_ (.A(_01151_),
    .Y(_04980_));
 NAND2x1_ASAP7_75t_R _22636_ (.A(net348),
    .B(_01149_),
    .Y(_04981_));
 OA211x2_ASAP7_75t_R _22637_ (.A1(net348),
    .A2(_04980_),
    .B(_04981_),
    .C(net325),
    .Y(_04982_));
 INVx1_ASAP7_75t_R _22638_ (.A(_01150_),
    .Y(_04983_));
 NAND2x1_ASAP7_75t_R _22639_ (.A(net348),
    .B(_01148_),
    .Y(_04984_));
 OA211x2_ASAP7_75t_R _22640_ (.A1(net348),
    .A2(_04983_),
    .B(_04984_),
    .C(net369),
    .Y(_04985_));
 OR3x1_ASAP7_75t_R _22641_ (.A(_13373_),
    .B(_04982_),
    .C(_04985_),
    .Y(_04986_));
 INVx1_ASAP7_75t_R _22642_ (.A(_01159_),
    .Y(_04987_));
 NAND2x1_ASAP7_75t_R _22643_ (.A(net348),
    .B(_01157_),
    .Y(_04988_));
 OA211x2_ASAP7_75t_R _22644_ (.A1(net348),
    .A2(_04987_),
    .B(_04988_),
    .C(net325),
    .Y(_04989_));
 INVx1_ASAP7_75t_R _22645_ (.A(_01158_),
    .Y(_04990_));
 NAND2x1_ASAP7_75t_R _22646_ (.A(net348),
    .B(_01156_),
    .Y(_04991_));
 OA211x2_ASAP7_75t_R _22647_ (.A1(net348),
    .A2(_04990_),
    .B(_04991_),
    .C(net369),
    .Y(_04992_));
 OR3x1_ASAP7_75t_R _22648_ (.A(net331),
    .B(_04989_),
    .C(_04992_),
    .Y(_04993_));
 AND3x1_ASAP7_75t_R _22649_ (.A(_13350_),
    .B(_04986_),
    .C(_04993_),
    .Y(_04994_));
 OR3x4_ASAP7_75t_R _22650_ (.A(_13355_),
    .B(_04979_),
    .C(_04994_),
    .Y(_04995_));
 INVx1_ASAP7_75t_R _22651_ (.A(_01167_),
    .Y(_04996_));
 NAND2x1_ASAP7_75t_R _22652_ (.A(net347),
    .B(_01165_),
    .Y(_04997_));
 OA211x2_ASAP7_75t_R _22653_ (.A1(net347),
    .A2(_04996_),
    .B(_04997_),
    .C(net325),
    .Y(_04998_));
 INVx1_ASAP7_75t_R _22654_ (.A(_01166_),
    .Y(_04999_));
 NAND2x1_ASAP7_75t_R _22655_ (.A(net347),
    .B(_01164_),
    .Y(_05000_));
 OA211x2_ASAP7_75t_R _22656_ (.A1(net347),
    .A2(_04999_),
    .B(_05000_),
    .C(net369),
    .Y(_05001_));
 OR3x1_ASAP7_75t_R _22657_ (.A(_13373_),
    .B(_04998_),
    .C(_05001_),
    .Y(_05002_));
 INVx1_ASAP7_75t_R _22658_ (.A(_01175_),
    .Y(_05003_));
 NAND2x1_ASAP7_75t_R _22659_ (.A(net347),
    .B(_01173_),
    .Y(_05004_));
 OA211x2_ASAP7_75t_R _22660_ (.A1(net347),
    .A2(_05003_),
    .B(_05004_),
    .C(net325),
    .Y(_05005_));
 INVx1_ASAP7_75t_R _22661_ (.A(_01174_),
    .Y(_05006_));
 NAND2x1_ASAP7_75t_R _22662_ (.A(net347),
    .B(_01172_),
    .Y(_05007_));
 OA211x2_ASAP7_75t_R _22663_ (.A1(net347),
    .A2(_05006_),
    .B(_05007_),
    .C(net369),
    .Y(_05008_));
 OR3x1_ASAP7_75t_R _22664_ (.A(net331),
    .B(_05005_),
    .C(_05008_),
    .Y(_05009_));
 AND3x1_ASAP7_75t_R _22665_ (.A(_13350_),
    .B(_05002_),
    .C(_05009_),
    .Y(_05010_));
 INVx1_ASAP7_75t_R _22666_ (.A(_01168_),
    .Y(_05011_));
 NOR2x1_ASAP7_75t_R _22667_ (.A(net347),
    .B(_01170_),
    .Y(_05012_));
 AO21x1_ASAP7_75t_R _22668_ (.A1(net347),
    .A2(_05011_),
    .B(_05012_),
    .Y(_05013_));
 INVx1_ASAP7_75t_R _22669_ (.A(_01171_),
    .Y(_05014_));
 NAND2x1_ASAP7_75t_R _22670_ (.A(net347),
    .B(_01169_),
    .Y(_05015_));
 OA211x2_ASAP7_75t_R _22671_ (.A1(net347),
    .A2(_05014_),
    .B(_05015_),
    .C(net325),
    .Y(_05016_));
 AO21x1_ASAP7_75t_R _22672_ (.A1(net369),
    .A2(_05013_),
    .B(_05016_),
    .Y(_05017_));
 TAPCELL_ASAP7_75t_R TAP_1074 ();
 INVx1_ASAP7_75t_R _22674_ (.A(_01163_),
    .Y(_05019_));
 NAND2x1_ASAP7_75t_R _22675_ (.A(net347),
    .B(_01161_),
    .Y(_05020_));
 OA211x2_ASAP7_75t_R _22676_ (.A1(net347),
    .A2(_05019_),
    .B(_05020_),
    .C(net325),
    .Y(_05021_));
 INVx1_ASAP7_75t_R _22677_ (.A(_01162_),
    .Y(_05022_));
 NAND2x1_ASAP7_75t_R _22678_ (.A(net347),
    .B(_01160_),
    .Y(_05023_));
 OA211x2_ASAP7_75t_R _22679_ (.A1(net347),
    .A2(_05022_),
    .B(_05023_),
    .C(net369),
    .Y(_05024_));
 OR3x1_ASAP7_75t_R _22680_ (.A(_13373_),
    .B(_05021_),
    .C(_05024_),
    .Y(_05025_));
 OA211x2_ASAP7_75t_R _22681_ (.A1(net331),
    .A2(_05017_),
    .B(_05025_),
    .C(net335),
    .Y(_05026_));
 OR3x4_ASAP7_75t_R _22682_ (.A(net327),
    .B(_05010_),
    .C(_05026_),
    .Y(_05027_));
 NAND2x2_ASAP7_75t_R _22683_ (.A(_04995_),
    .B(_05027_),
    .Y(_05028_));
 OA21x2_ASAP7_75t_R _22684_ (.A1(_01742_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_05029_));
 AO21x2_ASAP7_75t_R _22685_ (.A1(_13474_),
    .A2(_05028_),
    .B(_05029_),
    .Y(_05030_));
 TAPCELL_ASAP7_75t_R TAP_1073 ();
 INVx1_ASAP7_75t_R _22687_ (.A(_05030_),
    .Y(_18459_));
 INVx1_ASAP7_75t_R _22688_ (.A(_00224_),
    .Y(\cs_registers_i.pc_id_i[27] ));
 AND2x2_ASAP7_75t_R _22689_ (.A(net398),
    .B(_01682_),
    .Y(_05031_));
 AO21x1_ASAP7_75t_R _22690_ (.A1(net316),
    .A2(_01147_),
    .B(_05031_),
    .Y(_05032_));
 OAI22x1_ASAP7_75t_R _22691_ (.A1(_01146_),
    .A2(net2290),
    .B1(_05032_),
    .B2(net424),
    .Y(_05033_));
 NAND2x1_ASAP7_75t_R _22692_ (.A(net412),
    .B(_01149_),
    .Y(_05034_));
 OA211x2_ASAP7_75t_R _22693_ (.A1(net412),
    .A2(_04980_),
    .B(_05034_),
    .C(_13649_),
    .Y(_05035_));
 NAND2x1_ASAP7_75t_R _22694_ (.A(net412),
    .B(_01148_),
    .Y(_05036_));
 OA211x2_ASAP7_75t_R _22695_ (.A1(net412),
    .A2(_04983_),
    .B(_05036_),
    .C(net426),
    .Y(_05037_));
 OR3x1_ASAP7_75t_R _22696_ (.A(_13636_),
    .B(_05035_),
    .C(_05037_),
    .Y(_05038_));
 NAND2x1_ASAP7_75t_R _22697_ (.A(net412),
    .B(_01157_),
    .Y(_05039_));
 OA211x2_ASAP7_75t_R _22698_ (.A1(net412),
    .A2(_04987_),
    .B(_05039_),
    .C(_13649_),
    .Y(_05040_));
 NAND2x1_ASAP7_75t_R _22699_ (.A(net412),
    .B(_01156_),
    .Y(_05041_));
 OA211x2_ASAP7_75t_R _22700_ (.A1(net412),
    .A2(_04990_),
    .B(_05041_),
    .C(net426),
    .Y(_05042_));
 OR3x1_ASAP7_75t_R _22701_ (.A(net382),
    .B(_05040_),
    .C(_05042_),
    .Y(_05043_));
 AO21x1_ASAP7_75t_R _22702_ (.A1(_05038_),
    .A2(_05043_),
    .B(net387),
    .Y(_05044_));
 NAND2x1_ASAP7_75t_R _22703_ (.A(net410),
    .B(_01153_),
    .Y(_05045_));
 OA211x2_ASAP7_75t_R _22704_ (.A1(net410),
    .A2(_04972_),
    .B(_05045_),
    .C(_13649_),
    .Y(_05046_));
 NAND2x1_ASAP7_75t_R _22705_ (.A(net410),
    .B(_01152_),
    .Y(_05047_));
 OA211x2_ASAP7_75t_R _22706_ (.A1(net410),
    .A2(_04975_),
    .B(_05047_),
    .C(net424),
    .Y(_05048_));
 OR3x1_ASAP7_75t_R _22707_ (.A(_14942_),
    .B(_05046_),
    .C(_05048_),
    .Y(_05049_));
 OA211x2_ASAP7_75t_R _22708_ (.A1(net315),
    .A2(_05033_),
    .B(_05044_),
    .C(_05049_),
    .Y(_05050_));
 NOR2x1_ASAP7_75t_R _22709_ (.A(net424),
    .B(_01169_),
    .Y(_05051_));
 AO21x1_ASAP7_75t_R _22710_ (.A1(net424),
    .A2(_05011_),
    .B(_05051_),
    .Y(_05052_));
 INVx1_ASAP7_75t_R _22711_ (.A(_01173_),
    .Y(_05053_));
 NAND2x1_ASAP7_75t_R _22712_ (.A(net424),
    .B(_01172_),
    .Y(_05054_));
 OA211x2_ASAP7_75t_R _22713_ (.A1(net424),
    .A2(_05053_),
    .B(_05054_),
    .C(net321),
    .Y(_05055_));
 AO21x1_ASAP7_75t_R _22714_ (.A1(net386),
    .A2(_05052_),
    .B(_05055_),
    .Y(_05056_));
 NAND2x1_ASAP7_75t_R _22715_ (.A(net423),
    .B(_01170_),
    .Y(_05057_));
 OA211x2_ASAP7_75t_R _22716_ (.A1(net423),
    .A2(_05014_),
    .B(_05057_),
    .C(net386),
    .Y(_05058_));
 NAND2x1_ASAP7_75t_R _22717_ (.A(net424),
    .B(_01174_),
    .Y(_05059_));
 OA211x2_ASAP7_75t_R _22718_ (.A1(net424),
    .A2(_05003_),
    .B(_05059_),
    .C(net321),
    .Y(_05060_));
 OR3x1_ASAP7_75t_R _22719_ (.A(net410),
    .B(_05058_),
    .C(_05060_),
    .Y(_05061_));
 OA211x2_ASAP7_75t_R _22720_ (.A1(net316),
    .A2(_05056_),
    .B(_05061_),
    .C(_13636_),
    .Y(_05062_));
 NAND2x1_ASAP7_75t_R _22721_ (.A(net410),
    .B(_01164_),
    .Y(_05063_));
 OA211x2_ASAP7_75t_R _22722_ (.A1(net410),
    .A2(_04999_),
    .B(_05063_),
    .C(net321),
    .Y(_05064_));
 NAND2x1_ASAP7_75t_R _22723_ (.A(net410),
    .B(_01160_),
    .Y(_05065_));
 OA211x2_ASAP7_75t_R _22724_ (.A1(net410),
    .A2(_05022_),
    .B(_05065_),
    .C(net386),
    .Y(_05066_));
 OR3x1_ASAP7_75t_R _22725_ (.A(_13649_),
    .B(_05064_),
    .C(_05066_),
    .Y(_05067_));
 NAND2x1_ASAP7_75t_R _22726_ (.A(net410),
    .B(_01165_),
    .Y(_05068_));
 OA211x2_ASAP7_75t_R _22727_ (.A1(net410),
    .A2(_04996_),
    .B(_05068_),
    .C(net321),
    .Y(_05069_));
 NAND2x1_ASAP7_75t_R _22728_ (.A(net410),
    .B(_01161_),
    .Y(_05070_));
 OA211x2_ASAP7_75t_R _22729_ (.A1(net410),
    .A2(_05019_),
    .B(_05070_),
    .C(net386),
    .Y(_05071_));
 OR3x1_ASAP7_75t_R _22730_ (.A(net423),
    .B(_05069_),
    .C(_05071_),
    .Y(_05072_));
 AND3x1_ASAP7_75t_R _22731_ (.A(net382),
    .B(_05067_),
    .C(_05072_),
    .Y(_05073_));
 OR3x1_ASAP7_75t_R _22732_ (.A(net378),
    .B(_05062_),
    .C(_05073_),
    .Y(_05074_));
 OA21x2_ASAP7_75t_R _22733_ (.A1(_13626_),
    .A2(_05050_),
    .B(_05074_),
    .Y(_05075_));
 OAI22x1_ASAP7_75t_R _22734_ (.A1(_01614_),
    .A2(_13807_),
    .B1(_14103_),
    .B2(_00224_),
    .Y(_05076_));
 AO21x2_ASAP7_75t_R _22735_ (.A1(_13810_),
    .A2(_05075_),
    .B(_05076_),
    .Y(_05077_));
 TAPCELL_ASAP7_75t_R TAP_1072 ();
 INVx3_ASAP7_75t_R _22737_ (.A(_05077_),
    .Y(_18460_));
 AND2x2_ASAP7_75t_R _22738_ (.A(net346),
    .B(_01681_),
    .Y(_05078_));
 AO21x1_ASAP7_75t_R _22739_ (.A1(net2278),
    .A2(_01179_),
    .B(_05078_),
    .Y(_05079_));
 OAI22x1_ASAP7_75t_R _22740_ (.A1(_01178_),
    .A2(net311),
    .B1(_05079_),
    .B2(net369),
    .Y(_05080_));
 INVx1_ASAP7_75t_R _22741_ (.A(_01187_),
    .Y(_05081_));
 NAND2x1_ASAP7_75t_R _22742_ (.A(net2248),
    .B(_01185_),
    .Y(_05082_));
 OA211x2_ASAP7_75t_R _22743_ (.A1(net2248),
    .A2(_05081_),
    .B(_05082_),
    .C(net323),
    .Y(_05083_));
 INVx1_ASAP7_75t_R _22744_ (.A(_01186_),
    .Y(_05084_));
 NAND2x1_ASAP7_75t_R _22745_ (.A(net2248),
    .B(_01184_),
    .Y(_05085_));
 OA211x2_ASAP7_75t_R _22746_ (.A1(net2249),
    .A2(_05084_),
    .B(_05085_),
    .C(net375),
    .Y(_05086_));
 OR3x1_ASAP7_75t_R _22747_ (.A(net331),
    .B(_05083_),
    .C(_05086_),
    .Y(_05087_));
 OA211x2_ASAP7_75t_R _22748_ (.A1(_13373_),
    .A2(_05080_),
    .B(_05087_),
    .C(net336),
    .Y(_05088_));
 INVx1_ASAP7_75t_R _22749_ (.A(_01183_),
    .Y(_05089_));
 NAND2x1_ASAP7_75t_R _22750_ (.A(net2248),
    .B(_01181_),
    .Y(_05090_));
 OA211x2_ASAP7_75t_R _22751_ (.A1(net2248),
    .A2(_05089_),
    .B(_05090_),
    .C(net323),
    .Y(_05091_));
 INVx1_ASAP7_75t_R _22752_ (.A(_01182_),
    .Y(_05092_));
 NAND2x1_ASAP7_75t_R _22753_ (.A(net348),
    .B(_01180_),
    .Y(_05093_));
 OA211x2_ASAP7_75t_R _22754_ (.A1(net348),
    .A2(_05092_),
    .B(_05093_),
    .C(net375),
    .Y(_05094_));
 OR3x1_ASAP7_75t_R _22755_ (.A(_13373_),
    .B(_05091_),
    .C(_05094_),
    .Y(_05095_));
 INVx1_ASAP7_75t_R _22756_ (.A(_01191_),
    .Y(_05096_));
 NAND2x1_ASAP7_75t_R _22757_ (.A(net346),
    .B(_01189_),
    .Y(_05097_));
 OA211x2_ASAP7_75t_R _22758_ (.A1(net346),
    .A2(_05096_),
    .B(_05097_),
    .C(net323),
    .Y(_05098_));
 INVx1_ASAP7_75t_R _22759_ (.A(_01190_),
    .Y(_05099_));
 NAND2x1_ASAP7_75t_R _22760_ (.A(net346),
    .B(_01188_),
    .Y(_05100_));
 OA211x2_ASAP7_75t_R _22761_ (.A1(net346),
    .A2(_05099_),
    .B(_05100_),
    .C(net369),
    .Y(_05101_));
 OR3x1_ASAP7_75t_R _22762_ (.A(net331),
    .B(_05098_),
    .C(_05101_),
    .Y(_05102_));
 AND3x1_ASAP7_75t_R _22763_ (.A(_13350_),
    .B(_05095_),
    .C(_05102_),
    .Y(_05103_));
 OR3x4_ASAP7_75t_R _22764_ (.A(_13355_),
    .B(_05088_),
    .C(_05103_),
    .Y(_05104_));
 INVx1_ASAP7_75t_R _22765_ (.A(_01199_),
    .Y(_05105_));
 NAND2x1_ASAP7_75t_R _22766_ (.A(net348),
    .B(_01197_),
    .Y(_05106_));
 OA211x2_ASAP7_75t_R _22767_ (.A1(net348),
    .A2(_05105_),
    .B(_05106_),
    .C(net323),
    .Y(_05107_));
 INVx1_ASAP7_75t_R _22768_ (.A(_01198_),
    .Y(_05108_));
 NAND2x1_ASAP7_75t_R _22769_ (.A(net348),
    .B(_01196_),
    .Y(_05109_));
 OA211x2_ASAP7_75t_R _22770_ (.A1(net348),
    .A2(_05108_),
    .B(_05109_),
    .C(net375),
    .Y(_05110_));
 OR3x1_ASAP7_75t_R _22771_ (.A(_13373_),
    .B(_05107_),
    .C(_05110_),
    .Y(_05111_));
 INVx1_ASAP7_75t_R _22772_ (.A(_01207_),
    .Y(_05112_));
 NAND2x1_ASAP7_75t_R _22773_ (.A(net348),
    .B(_01205_),
    .Y(_05113_));
 OA211x2_ASAP7_75t_R _22774_ (.A1(net348),
    .A2(_05112_),
    .B(_05113_),
    .C(net323),
    .Y(_05114_));
 INVx1_ASAP7_75t_R _22775_ (.A(_01206_),
    .Y(_05115_));
 NAND2x1_ASAP7_75t_R _22776_ (.A(net348),
    .B(_01204_),
    .Y(_05116_));
 OA211x2_ASAP7_75t_R _22777_ (.A1(net348),
    .A2(_05115_),
    .B(_05116_),
    .C(net375),
    .Y(_05117_));
 OR3x1_ASAP7_75t_R _22778_ (.A(net331),
    .B(_05114_),
    .C(_05117_),
    .Y(_05118_));
 AND3x1_ASAP7_75t_R _22779_ (.A(_13350_),
    .B(_05111_),
    .C(_05118_),
    .Y(_05119_));
 INVx1_ASAP7_75t_R _22780_ (.A(_01195_),
    .Y(_05120_));
 NAND2x1_ASAP7_75t_R _22781_ (.A(net352),
    .B(_01193_),
    .Y(_05121_));
 OA211x2_ASAP7_75t_R _22782_ (.A1(net352),
    .A2(_05120_),
    .B(_05121_),
    .C(net323),
    .Y(_05122_));
 INVx1_ASAP7_75t_R _22783_ (.A(_01194_),
    .Y(_05123_));
 NAND2x1_ASAP7_75t_R _22784_ (.A(net352),
    .B(_01192_),
    .Y(_05124_));
 OA211x2_ASAP7_75t_R _22785_ (.A1(net352),
    .A2(_05123_),
    .B(_05124_),
    .C(net375),
    .Y(_05125_));
 OR3x1_ASAP7_75t_R _22786_ (.A(_13373_),
    .B(_05122_),
    .C(_05125_),
    .Y(_05126_));
 INVx1_ASAP7_75t_R _22787_ (.A(_01203_),
    .Y(_05127_));
 NAND2x1_ASAP7_75t_R _22788_ (.A(net352),
    .B(_01201_),
    .Y(_05128_));
 OA211x2_ASAP7_75t_R _22789_ (.A1(net352),
    .A2(_05127_),
    .B(_05128_),
    .C(net323),
    .Y(_05129_));
 INVx1_ASAP7_75t_R _22790_ (.A(_01202_),
    .Y(_05130_));
 NAND2x1_ASAP7_75t_R _22791_ (.A(net352),
    .B(_01200_),
    .Y(_05131_));
 OA211x2_ASAP7_75t_R _22792_ (.A1(net352),
    .A2(_05130_),
    .B(_05131_),
    .C(net374),
    .Y(_05132_));
 OR3x1_ASAP7_75t_R _22793_ (.A(net331),
    .B(_05129_),
    .C(_05132_),
    .Y(_05133_));
 AND3x1_ASAP7_75t_R _22794_ (.A(net335),
    .B(_05126_),
    .C(_05133_),
    .Y(_05134_));
 OR3x4_ASAP7_75t_R _22795_ (.A(net327),
    .B(_05119_),
    .C(_05134_),
    .Y(_05135_));
 NAND2x2_ASAP7_75t_R _22796_ (.A(_05104_),
    .B(_05135_),
    .Y(_05136_));
 OA21x2_ASAP7_75t_R _22797_ (.A1(_01741_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_05137_));
 AO21x2_ASAP7_75t_R _22798_ (.A1(_13474_),
    .A2(_05136_),
    .B(_05137_),
    .Y(_05138_));
 TAPCELL_ASAP7_75t_R TAP_1071 ();
 INVx1_ASAP7_75t_R _22800_ (.A(_05138_),
    .Y(_18465_));
 AND2x2_ASAP7_75t_R _22801_ (.A(_00226_),
    .B(_13993_),
    .Y(_05139_));
 NAND2x1_ASAP7_75t_R _22802_ (.A(net398),
    .B(_01201_),
    .Y(_05140_));
 OA211x2_ASAP7_75t_R _22803_ (.A1(net398),
    .A2(_05127_),
    .B(_05140_),
    .C(net318),
    .Y(_05141_));
 NAND2x1_ASAP7_75t_R _22804_ (.A(net398),
    .B(_01200_),
    .Y(_05142_));
 OA211x2_ASAP7_75t_R _22805_ (.A1(net398),
    .A2(_05130_),
    .B(_05142_),
    .C(net424),
    .Y(_05143_));
 OR3x1_ASAP7_75t_R _22806_ (.A(net320),
    .B(_05141_),
    .C(_05143_),
    .Y(_05144_));
 NAND2x1_ASAP7_75t_R _22807_ (.A(net410),
    .B(_01205_),
    .Y(_05145_));
 OA211x2_ASAP7_75t_R _22808_ (.A1(net410),
    .A2(_05112_),
    .B(_05145_),
    .C(net318),
    .Y(_05146_));
 NAND2x1_ASAP7_75t_R _22809_ (.A(net410),
    .B(_01204_),
    .Y(_05147_));
 OA211x2_ASAP7_75t_R _22810_ (.A1(net410),
    .A2(_05115_),
    .B(_05147_),
    .C(net424),
    .Y(_05148_));
 OR3x1_ASAP7_75t_R _22811_ (.A(net386),
    .B(_05146_),
    .C(_05148_),
    .Y(_05149_));
 AO21x1_ASAP7_75t_R _22812_ (.A1(_05144_),
    .A2(_05149_),
    .B(net380),
    .Y(_05150_));
 NAND2x1_ASAP7_75t_R _22813_ (.A(net410),
    .B(_01197_),
    .Y(_05151_));
 OA211x2_ASAP7_75t_R _22814_ (.A1(net410),
    .A2(_05105_),
    .B(_05151_),
    .C(net318),
    .Y(_05152_));
 NAND2x1_ASAP7_75t_R _22815_ (.A(net410),
    .B(_01196_),
    .Y(_05153_));
 OA211x2_ASAP7_75t_R _22816_ (.A1(net410),
    .A2(_05108_),
    .B(_05153_),
    .C(net424),
    .Y(_05154_));
 OR3x1_ASAP7_75t_R _22817_ (.A(_14015_),
    .B(_05152_),
    .C(_05154_),
    .Y(_05155_));
 NAND2x1_ASAP7_75t_R _22818_ (.A(net398),
    .B(_01193_),
    .Y(_05156_));
 OA211x2_ASAP7_75t_R _22819_ (.A1(net398),
    .A2(_05120_),
    .B(_05156_),
    .C(net318),
    .Y(_05157_));
 NAND2x1_ASAP7_75t_R _22820_ (.A(net398),
    .B(_01192_),
    .Y(_05158_));
 OA211x2_ASAP7_75t_R _22821_ (.A1(net398),
    .A2(_05123_),
    .B(_05158_),
    .C(net424),
    .Y(_05159_));
 OR3x1_ASAP7_75t_R _22822_ (.A(net315),
    .B(_05157_),
    .C(_05159_),
    .Y(_05160_));
 AND3x1_ASAP7_75t_R _22823_ (.A(_13626_),
    .B(_05155_),
    .C(_05160_),
    .Y(_05161_));
 NAND2x1_ASAP7_75t_R _22824_ (.A(net412),
    .B(_01181_),
    .Y(_05162_));
 OA211x2_ASAP7_75t_R _22825_ (.A1(net412),
    .A2(_05089_),
    .B(_05162_),
    .C(net318),
    .Y(_05163_));
 NAND2x1_ASAP7_75t_R _22826_ (.A(net412),
    .B(_01180_),
    .Y(_05164_));
 OA211x2_ASAP7_75t_R _22827_ (.A1(net412),
    .A2(_05092_),
    .B(_05164_),
    .C(net424),
    .Y(_05165_));
 OR3x1_ASAP7_75t_R _22828_ (.A(_13636_),
    .B(_05163_),
    .C(_05165_),
    .Y(_05166_));
 NAND2x1_ASAP7_75t_R _22829_ (.A(net413),
    .B(_01189_),
    .Y(_05167_));
 OA211x2_ASAP7_75t_R _22830_ (.A1(net413),
    .A2(_05096_),
    .B(_05167_),
    .C(net318),
    .Y(_05168_));
 NAND2x1_ASAP7_75t_R _22831_ (.A(net416),
    .B(_01188_),
    .Y(_05169_));
 OA211x2_ASAP7_75t_R _22832_ (.A1(net416),
    .A2(_05099_),
    .B(_05169_),
    .C(net426),
    .Y(_05170_));
 OR3x1_ASAP7_75t_R _22833_ (.A(net382),
    .B(_05168_),
    .C(_05170_),
    .Y(_05171_));
 AO21x1_ASAP7_75t_R _22834_ (.A1(_05166_),
    .A2(_05171_),
    .B(net386),
    .Y(_05172_));
 AND2x2_ASAP7_75t_R _22835_ (.A(net416),
    .B(_01681_),
    .Y(_05173_));
 AO21x1_ASAP7_75t_R _22836_ (.A1(net316),
    .A2(_01179_),
    .B(_05173_),
    .Y(_05174_));
 OAI22x1_ASAP7_75t_R _22837_ (.A1(_01178_),
    .A2(net2290),
    .B1(_05174_),
    .B2(net426),
    .Y(_05175_));
 NAND2x1_ASAP7_75t_R _22838_ (.A(net413),
    .B(_01185_),
    .Y(_05176_));
 OA211x2_ASAP7_75t_R _22839_ (.A1(net413),
    .A2(_05081_),
    .B(_05176_),
    .C(net318),
    .Y(_05177_));
 NAND2x1_ASAP7_75t_R _22840_ (.A(net413),
    .B(_01184_),
    .Y(_05178_));
 OA211x2_ASAP7_75t_R _22841_ (.A1(net413),
    .A2(_05084_),
    .B(_05178_),
    .C(net426),
    .Y(_05179_));
 OR3x1_ASAP7_75t_R _22842_ (.A(_14942_),
    .B(_05177_),
    .C(_05179_),
    .Y(_05180_));
 OA211x2_ASAP7_75t_R _22843_ (.A1(net315),
    .A2(_05175_),
    .B(_05180_),
    .C(net378),
    .Y(_05181_));
 AOI221x1_ASAP7_75t_R _22844_ (.A1(_05150_),
    .A2(_05161_),
    .B1(_05172_),
    .B2(_05181_),
    .C(_13993_),
    .Y(_05182_));
 OR3x2_ASAP7_75t_R _22845_ (.A(_14988_),
    .B(_05139_),
    .C(_05182_),
    .Y(_05183_));
 OA21x2_ASAP7_75t_R _22846_ (.A1(_01613_),
    .A2(_13807_),
    .B(_05183_),
    .Y(_05184_));
 TAPCELL_ASAP7_75t_R TAP_1070 ();
 XNOR2x2_ASAP7_75t_R _22848_ (.A(_01211_),
    .B(_01209_),
    .Y(_05185_));
 INVx6_ASAP7_75t_R _22849_ (.A(_05185_),
    .Y(net169));
 AND2x2_ASAP7_75t_R _22850_ (.A(net357),
    .B(_01680_),
    .Y(_05186_));
 AO21x1_ASAP7_75t_R _22851_ (.A1(net2260),
    .A2(_01213_),
    .B(_05186_),
    .Y(_05187_));
 OAI22x1_ASAP7_75t_R _22852_ (.A1(_01212_),
    .A2(_14184_),
    .B1(_05187_),
    .B2(net372),
    .Y(_05188_));
 INVx1_ASAP7_75t_R _22853_ (.A(_01221_),
    .Y(_05189_));
 NAND2x1_ASAP7_75t_R _22854_ (.A(net356),
    .B(_01219_),
    .Y(_05190_));
 OA211x2_ASAP7_75t_R _22855_ (.A1(net356),
    .A2(_05189_),
    .B(_05190_),
    .C(net324),
    .Y(_05191_));
 INVx1_ASAP7_75t_R _22856_ (.A(_01220_),
    .Y(_05192_));
 NAND2x1_ASAP7_75t_R _22857_ (.A(net356),
    .B(_01218_),
    .Y(_05193_));
 OA211x2_ASAP7_75t_R _22858_ (.A1(net356),
    .A2(_05192_),
    .B(_05193_),
    .C(net373),
    .Y(_05194_));
 OR3x1_ASAP7_75t_R _22859_ (.A(net330),
    .B(_05191_),
    .C(_05194_),
    .Y(_05195_));
 OA21x2_ASAP7_75t_R _22860_ (.A1(_13373_),
    .A2(_05188_),
    .B(_05195_),
    .Y(_05196_));
 INVx1_ASAP7_75t_R _22861_ (.A(_01217_),
    .Y(_05197_));
 NAND2x1_ASAP7_75t_R _22862_ (.A(net357),
    .B(_01215_),
    .Y(_05198_));
 OA211x2_ASAP7_75t_R _22863_ (.A1(net357),
    .A2(_05197_),
    .B(_05198_),
    .C(net324),
    .Y(_05199_));
 INVx1_ASAP7_75t_R _22864_ (.A(_01216_),
    .Y(_05200_));
 NAND2x1_ASAP7_75t_R _22865_ (.A(net357),
    .B(_01214_),
    .Y(_05201_));
 OA211x2_ASAP7_75t_R _22866_ (.A1(net357),
    .A2(_05200_),
    .B(_05201_),
    .C(net372),
    .Y(_05202_));
 OR3x1_ASAP7_75t_R _22867_ (.A(_13373_),
    .B(_05199_),
    .C(_05202_),
    .Y(_05203_));
 INVx1_ASAP7_75t_R _22868_ (.A(_01225_),
    .Y(_05204_));
 NAND2x1_ASAP7_75t_R _22869_ (.A(net356),
    .B(_01223_),
    .Y(_05205_));
 OA211x2_ASAP7_75t_R _22870_ (.A1(net356),
    .A2(_05204_),
    .B(_05205_),
    .C(net324),
    .Y(_05206_));
 INVx1_ASAP7_75t_R _22871_ (.A(_01224_),
    .Y(_05207_));
 NAND2x1_ASAP7_75t_R _22872_ (.A(net356),
    .B(_01222_),
    .Y(_05208_));
 OA211x2_ASAP7_75t_R _22873_ (.A1(net356),
    .A2(_05207_),
    .B(_05208_),
    .C(net373),
    .Y(_05209_));
 OR3x1_ASAP7_75t_R _22874_ (.A(net330),
    .B(_05206_),
    .C(_05209_),
    .Y(_05210_));
 AND3x1_ASAP7_75t_R _22875_ (.A(_13350_),
    .B(_05203_),
    .C(_05210_),
    .Y(_05211_));
 AO21x1_ASAP7_75t_R _22876_ (.A1(net334),
    .A2(_05196_),
    .B(_05211_),
    .Y(_05212_));
 INVx1_ASAP7_75t_R _22877_ (.A(_01234_),
    .Y(_05213_));
 NOR2x1_ASAP7_75t_R _22878_ (.A(net356),
    .B(_01236_),
    .Y(_05214_));
 AO21x1_ASAP7_75t_R _22879_ (.A1(net356),
    .A2(_05213_),
    .B(_05214_),
    .Y(_05215_));
 INVx1_ASAP7_75t_R _22880_ (.A(_01237_),
    .Y(_05216_));
 NAND2x1_ASAP7_75t_R _22881_ (.A(net356),
    .B(_01235_),
    .Y(_05217_));
 OA211x2_ASAP7_75t_R _22882_ (.A1(net356),
    .A2(_05216_),
    .B(_05217_),
    .C(net324),
    .Y(_05218_));
 AO21x1_ASAP7_75t_R _22883_ (.A1(net372),
    .A2(_05215_),
    .B(_05218_),
    .Y(_05219_));
 INVx1_ASAP7_75t_R _22884_ (.A(_01241_),
    .Y(_05220_));
 NAND2x1_ASAP7_75t_R _22885_ (.A(net356),
    .B(_01239_),
    .Y(_05221_));
 OA211x2_ASAP7_75t_R _22886_ (.A1(net356),
    .A2(_05220_),
    .B(_05221_),
    .C(net324),
    .Y(_05222_));
 INVx1_ASAP7_75t_R _22887_ (.A(_01240_),
    .Y(_05223_));
 NAND2x1_ASAP7_75t_R _22888_ (.A(net356),
    .B(_01238_),
    .Y(_05224_));
 OA211x2_ASAP7_75t_R _22889_ (.A1(net356),
    .A2(_05223_),
    .B(_05224_),
    .C(net372),
    .Y(_05225_));
 OR3x1_ASAP7_75t_R _22890_ (.A(net334),
    .B(_05222_),
    .C(_05225_),
    .Y(_05226_));
 OA211x2_ASAP7_75t_R _22891_ (.A1(_13350_),
    .A2(_05219_),
    .B(_05226_),
    .C(_13373_),
    .Y(_05227_));
 INVx1_ASAP7_75t_R _22892_ (.A(_01229_),
    .Y(_05228_));
 NAND2x1_ASAP7_75t_R _22893_ (.A(net357),
    .B(_01227_),
    .Y(_05229_));
 OA211x2_ASAP7_75t_R _22894_ (.A1(net357),
    .A2(_05228_),
    .B(_05229_),
    .C(net324),
    .Y(_05230_));
 INVx1_ASAP7_75t_R _22895_ (.A(_01228_),
    .Y(_05231_));
 NAND2x1_ASAP7_75t_R _22896_ (.A(net357),
    .B(_01226_),
    .Y(_05232_));
 OA211x2_ASAP7_75t_R _22897_ (.A1(net357),
    .A2(_05231_),
    .B(_05232_),
    .C(net372),
    .Y(_05233_));
 OR3x1_ASAP7_75t_R _22898_ (.A(_13350_),
    .B(_05230_),
    .C(_05233_),
    .Y(_05234_));
 INVx1_ASAP7_75t_R _22899_ (.A(_01233_),
    .Y(_05235_));
 NAND2x1_ASAP7_75t_R _22900_ (.A(net357),
    .B(_01231_),
    .Y(_05236_));
 OA211x2_ASAP7_75t_R _22901_ (.A1(net357),
    .A2(_05235_),
    .B(_05236_),
    .C(net324),
    .Y(_05237_));
 INVx1_ASAP7_75t_R _22902_ (.A(_01232_),
    .Y(_05238_));
 NAND2x1_ASAP7_75t_R _22903_ (.A(net356),
    .B(_01230_),
    .Y(_05239_));
 OA211x2_ASAP7_75t_R _22904_ (.A1(net356),
    .A2(_05238_),
    .B(_05239_),
    .C(net372),
    .Y(_05240_));
 OR3x1_ASAP7_75t_R _22905_ (.A(net334),
    .B(_05237_),
    .C(_05240_),
    .Y(_05241_));
 AND3x1_ASAP7_75t_R _22906_ (.A(net329),
    .B(_05234_),
    .C(_05241_),
    .Y(_05242_));
 OR3x1_ASAP7_75t_R _22907_ (.A(net327),
    .B(_05227_),
    .C(_05242_),
    .Y(_05243_));
 OA21x2_ASAP7_75t_R _22908_ (.A1(_13355_),
    .A2(_05212_),
    .B(_05243_),
    .Y(_05244_));
 INVx3_ASAP7_75t_R _22909_ (.A(_05244_),
    .Y(_05245_));
 OA21x2_ASAP7_75t_R _22910_ (.A1(_01740_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_05246_));
 AO21x2_ASAP7_75t_R _22911_ (.A1(_13474_),
    .A2(_05245_),
    .B(_05246_),
    .Y(_05247_));
 TAPCELL_ASAP7_75t_R TAP_1069 ();
 INVx1_ASAP7_75t_R _22913_ (.A(_05247_),
    .Y(_18470_));
 INVx1_ASAP7_75t_R _22914_ (.A(_00227_),
    .Y(\cs_registers_i.pc_id_i[29] ));
 NAND2x1_ASAP7_75t_R _22915_ (.A(net402),
    .B(_01223_),
    .Y(_05248_));
 OA21x2_ASAP7_75t_R _22916_ (.A1(net2376),
    .A2(_05204_),
    .B(_05248_),
    .Y(_05249_));
 NAND2x1_ASAP7_75t_R _22917_ (.A(net402),
    .B(_01219_),
    .Y(_05250_));
 OA211x2_ASAP7_75t_R _22918_ (.A1(net402),
    .A2(_05189_),
    .B(_05250_),
    .C(net384),
    .Y(_05251_));
 AO21x1_ASAP7_75t_R _22919_ (.A1(net320),
    .A2(_05249_),
    .B(_05251_),
    .Y(_05252_));
 NAND2x1_ASAP7_75t_R _22920_ (.A(net403),
    .B(_01222_),
    .Y(_05253_));
 OA211x2_ASAP7_75t_R _22921_ (.A1(net403),
    .A2(_05207_),
    .B(_05253_),
    .C(net320),
    .Y(_05254_));
 NAND2x1_ASAP7_75t_R _22922_ (.A(net403),
    .B(_01218_),
    .Y(_05255_));
 OA211x2_ASAP7_75t_R _22923_ (.A1(net403),
    .A2(_05192_),
    .B(_05255_),
    .C(net384),
    .Y(_05256_));
 OR3x1_ASAP7_75t_R _22924_ (.A(net317),
    .B(_05254_),
    .C(_05256_),
    .Y(_05257_));
 OA21x2_ASAP7_75t_R _22925_ (.A1(net420),
    .A2(_05252_),
    .B(_05257_),
    .Y(_05258_));
 NAND2x1_ASAP7_75t_R _22926_ (.A(net317),
    .B(_01235_),
    .Y(_05259_));
 OA211x2_ASAP7_75t_R _22927_ (.A1(net317),
    .A2(_05213_),
    .B(_05259_),
    .C(net384),
    .Y(_05260_));
 AND2x2_ASAP7_75t_R _22928_ (.A(net420),
    .B(_01238_),
    .Y(_05261_));
 AO21x1_ASAP7_75t_R _22929_ (.A1(net317),
    .A2(_01239_),
    .B(_05261_),
    .Y(_05262_));
 OAI21x1_ASAP7_75t_R _22930_ (.A1(net384),
    .A2(_05262_),
    .B(net403),
    .Y(_05263_));
 NAND2x1_ASAP7_75t_R _22931_ (.A(net420),
    .B(_01236_),
    .Y(_05264_));
 OA211x2_ASAP7_75t_R _22932_ (.A1(net420),
    .A2(_05216_),
    .B(_05264_),
    .C(net384),
    .Y(_05265_));
 NAND2x1_ASAP7_75t_R _22933_ (.A(net420),
    .B(_01240_),
    .Y(_05266_));
 OA211x2_ASAP7_75t_R _22934_ (.A1(net420),
    .A2(_05220_),
    .B(_05266_),
    .C(net320),
    .Y(_05267_));
 OR3x1_ASAP7_75t_R _22935_ (.A(net403),
    .B(_05265_),
    .C(_05267_),
    .Y(_05268_));
 OA211x2_ASAP7_75t_R _22936_ (.A1(_05260_),
    .A2(_05263_),
    .B(_05268_),
    .C(_13626_),
    .Y(_05269_));
 AOI211x1_ASAP7_75t_R _22937_ (.A1(net377),
    .A2(_05258_),
    .B(_05269_),
    .C(net380),
    .Y(_05270_));
 NAND2x1_ASAP7_75t_R _22938_ (.A(net2352),
    .B(_01215_),
    .Y(_05271_));
 OA211x2_ASAP7_75t_R _22939_ (.A1(net2352),
    .A2(_05197_),
    .B(_05271_),
    .C(net317),
    .Y(_05272_));
 NAND2x1_ASAP7_75t_R _22940_ (.A(net2352),
    .B(_01214_),
    .Y(_05273_));
 OA211x2_ASAP7_75t_R _22941_ (.A1(net2352),
    .A2(_05200_),
    .B(_05273_),
    .C(net420),
    .Y(_05274_));
 INVx1_ASAP7_75t_R _22942_ (.A(_01213_),
    .Y(_05275_));
 NAND2x1_ASAP7_75t_R _22943_ (.A(net2352),
    .B(_01680_),
    .Y(_05276_));
 OA211x2_ASAP7_75t_R _22944_ (.A1(net2352),
    .A2(_05275_),
    .B(_05276_),
    .C(net317),
    .Y(_05277_));
 NOR2x1_ASAP7_75t_R _22945_ (.A(_01212_),
    .B(net2292),
    .Y(_05278_));
 OA33x2_ASAP7_75t_R _22946_ (.A1(net312),
    .A2(_05272_),
    .A3(_05274_),
    .B1(_05277_),
    .B2(_05278_),
    .B3(_14005_),
    .Y(_05279_));
 NAND2x1_ASAP7_75t_R _22947_ (.A(net404),
    .B(_01227_),
    .Y(_05280_));
 OA211x2_ASAP7_75t_R _22948_ (.A1(net404),
    .A2(_05228_),
    .B(_05280_),
    .C(net317),
    .Y(_05281_));
 NAND2x1_ASAP7_75t_R _22949_ (.A(net404),
    .B(_01226_),
    .Y(_05282_));
 OA211x2_ASAP7_75t_R _22950_ (.A1(net404),
    .A2(_05231_),
    .B(_05282_),
    .C(net420),
    .Y(_05283_));
 OR3x1_ASAP7_75t_R _22951_ (.A(net321),
    .B(_05281_),
    .C(_05283_),
    .Y(_05284_));
 NAND2x1_ASAP7_75t_R _22952_ (.A(net404),
    .B(_01231_),
    .Y(_05285_));
 OA211x2_ASAP7_75t_R _22953_ (.A1(net404),
    .A2(_05235_),
    .B(_05285_),
    .C(net317),
    .Y(_05286_));
 NAND2x1_ASAP7_75t_R _22954_ (.A(net404),
    .B(_01230_),
    .Y(_05287_));
 OA211x2_ASAP7_75t_R _22955_ (.A1(net404),
    .A2(_05238_),
    .B(_05287_),
    .C(net420),
    .Y(_05288_));
 OR3x1_ASAP7_75t_R _22956_ (.A(net383),
    .B(_05286_),
    .C(_05288_),
    .Y(_05289_));
 AO21x1_ASAP7_75t_R _22957_ (.A1(_05284_),
    .A2(_05289_),
    .B(_14049_),
    .Y(_05290_));
 OAI21x1_ASAP7_75t_R _22958_ (.A1(_13626_),
    .A2(_05279_),
    .B(_05290_),
    .Y(_05291_));
 OR4x2_ASAP7_75t_R _22959_ (.A(_13993_),
    .B(_14988_),
    .C(_05270_),
    .D(_05291_),
    .Y(_05292_));
 OR3x1_ASAP7_75t_R _22960_ (.A(_00227_),
    .B(_13808_),
    .C(_14988_),
    .Y(_05293_));
 OA21x2_ASAP7_75t_R _22961_ (.A1(_01612_),
    .A2(_13807_),
    .B(_05293_),
    .Y(_05294_));
 NAND2x2_ASAP7_75t_R _22962_ (.A(_05292_),
    .B(_05294_),
    .Y(_18471_));
 INVx3_ASAP7_75t_R _22963_ (.A(_18471_),
    .Y(_18469_));
 INVx1_ASAP7_75t_R _22964_ (.A(_01253_),
    .Y(_05295_));
 NAND2x1_ASAP7_75t_R _22965_ (.A(net341),
    .B(_01251_),
    .Y(_05296_));
 OA211x2_ASAP7_75t_R _22966_ (.A1(net341),
    .A2(_05295_),
    .B(_05296_),
    .C(net323),
    .Y(_05297_));
 INVx1_ASAP7_75t_R _22967_ (.A(_01252_),
    .Y(_05298_));
 NAND2x1_ASAP7_75t_R _22968_ (.A(net341),
    .B(_01250_),
    .Y(_05299_));
 OA211x2_ASAP7_75t_R _22969_ (.A1(net341),
    .A2(_05298_),
    .B(_05299_),
    .C(net370),
    .Y(_05300_));
 OR3x1_ASAP7_75t_R _22970_ (.A(net331),
    .B(_05297_),
    .C(_05300_),
    .Y(_05301_));
 INVx1_ASAP7_75t_R _22971_ (.A(_01244_),
    .Y(_05302_));
 INVx1_ASAP7_75t_R _22972_ (.A(_01245_),
    .Y(_05303_));
 NAND2x1_ASAP7_75t_R _22973_ (.A(net341),
    .B(_01679_),
    .Y(_05304_));
 OA21x2_ASAP7_75t_R _22974_ (.A1(net341),
    .A2(_05303_),
    .B(_05304_),
    .Y(_05305_));
 AO221x1_ASAP7_75t_R _22975_ (.A1(_05302_),
    .A2(net2215),
    .B1(_05305_),
    .B2(net323),
    .C(_13373_),
    .Y(_05306_));
 AO21x1_ASAP7_75t_R _22976_ (.A1(_05301_),
    .A2(_05306_),
    .B(_13350_),
    .Y(_05307_));
 INVx1_ASAP7_75t_R _22977_ (.A(_01249_),
    .Y(_05308_));
 NAND2x1_ASAP7_75t_R _22978_ (.A(net339),
    .B(_01247_),
    .Y(_05309_));
 OA211x2_ASAP7_75t_R _22979_ (.A1(net339),
    .A2(_05308_),
    .B(_05309_),
    .C(net323),
    .Y(_05310_));
 INVx1_ASAP7_75t_R _22980_ (.A(_01248_),
    .Y(_05311_));
 NAND2x1_ASAP7_75t_R _22981_ (.A(net339),
    .B(_01246_),
    .Y(_05312_));
 OA211x2_ASAP7_75t_R _22982_ (.A1(net339),
    .A2(_05311_),
    .B(_05312_),
    .C(net369),
    .Y(_05313_));
 OR3x1_ASAP7_75t_R _22983_ (.A(_13373_),
    .B(_05310_),
    .C(_05313_),
    .Y(_05314_));
 INVx1_ASAP7_75t_R _22984_ (.A(_01257_),
    .Y(_05315_));
 NAND2x1_ASAP7_75t_R _22985_ (.A(net339),
    .B(_01255_),
    .Y(_05316_));
 OA211x2_ASAP7_75t_R _22986_ (.A1(net339),
    .A2(_05315_),
    .B(_05316_),
    .C(net323),
    .Y(_05317_));
 INVx1_ASAP7_75t_R _22987_ (.A(_01256_),
    .Y(_05318_));
 NAND2x1_ASAP7_75t_R _22988_ (.A(net339),
    .B(_01254_),
    .Y(_05319_));
 OA211x2_ASAP7_75t_R _22989_ (.A1(net339),
    .A2(_05318_),
    .B(_05319_),
    .C(net369),
    .Y(_05320_));
 OR3x1_ASAP7_75t_R _22990_ (.A(net331),
    .B(_05317_),
    .C(_05320_),
    .Y(_05321_));
 AO21x1_ASAP7_75t_R _22991_ (.A1(_05314_),
    .A2(_05321_),
    .B(net337),
    .Y(_05322_));
 AO21x2_ASAP7_75t_R _22992_ (.A1(_05307_),
    .A2(_05322_),
    .B(_13355_),
    .Y(_05323_));
 INVx1_ASAP7_75t_R _22993_ (.A(_01265_),
    .Y(_05324_));
 NAND2x1_ASAP7_75t_R _22994_ (.A(net346),
    .B(_01263_),
    .Y(_05325_));
 OA211x2_ASAP7_75t_R _22995_ (.A1(net346),
    .A2(_05324_),
    .B(_05325_),
    .C(net323),
    .Y(_05326_));
 INVx1_ASAP7_75t_R _22996_ (.A(_01264_),
    .Y(_05327_));
 NAND2x1_ASAP7_75t_R _22997_ (.A(net346),
    .B(_01262_),
    .Y(_05328_));
 OA211x2_ASAP7_75t_R _22998_ (.A1(net346),
    .A2(_05327_),
    .B(_05328_),
    .C(net369),
    .Y(_05329_));
 OR3x1_ASAP7_75t_R _22999_ (.A(net337),
    .B(_05326_),
    .C(_05329_),
    .Y(_05330_));
 INVx1_ASAP7_75t_R _23000_ (.A(_01261_),
    .Y(_05331_));
 NAND2x1_ASAP7_75t_R _23001_ (.A(net2248),
    .B(_01259_),
    .Y(_05332_));
 OA211x2_ASAP7_75t_R _23002_ (.A1(net2249),
    .A2(_05331_),
    .B(_05332_),
    .C(net323),
    .Y(_05333_));
 INVx1_ASAP7_75t_R _23003_ (.A(_01260_),
    .Y(_05334_));
 NAND2x1_ASAP7_75t_R _23004_ (.A(net2248),
    .B(_01258_),
    .Y(_05335_));
 OA211x2_ASAP7_75t_R _23005_ (.A1(net2249),
    .A2(_05334_),
    .B(_05335_),
    .C(net369),
    .Y(_05336_));
 OR3x1_ASAP7_75t_R _23006_ (.A(_13350_),
    .B(_05333_),
    .C(_05336_),
    .Y(_05337_));
 AND3x1_ASAP7_75t_R _23007_ (.A(net331),
    .B(_05330_),
    .C(_05337_),
    .Y(_05338_));
 INVx1_ASAP7_75t_R _23008_ (.A(_01269_),
    .Y(_05339_));
 NAND2x1_ASAP7_75t_R _23009_ (.A(net348),
    .B(_01267_),
    .Y(_05340_));
 OA211x2_ASAP7_75t_R _23010_ (.A1(net347),
    .A2(_05339_),
    .B(_05340_),
    .C(net323),
    .Y(_05341_));
 INVx1_ASAP7_75t_R _23011_ (.A(_01268_),
    .Y(_05342_));
 NAND2x1_ASAP7_75t_R _23012_ (.A(net347),
    .B(_01266_),
    .Y(_05343_));
 OA211x2_ASAP7_75t_R _23013_ (.A1(net347),
    .A2(_05342_),
    .B(_05343_),
    .C(net375),
    .Y(_05344_));
 OR3x1_ASAP7_75t_R _23014_ (.A(_13350_),
    .B(_05341_),
    .C(_05344_),
    .Y(_05345_));
 INVx1_ASAP7_75t_R _23015_ (.A(_01273_),
    .Y(_05346_));
 NAND2x1_ASAP7_75t_R _23016_ (.A(net339),
    .B(_01271_),
    .Y(_05347_));
 OA211x2_ASAP7_75t_R _23017_ (.A1(net339),
    .A2(_05346_),
    .B(_05347_),
    .C(net323),
    .Y(_05348_));
 INVx1_ASAP7_75t_R _23018_ (.A(_01272_),
    .Y(_05349_));
 NAND2x1_ASAP7_75t_R _23019_ (.A(net346),
    .B(_01270_),
    .Y(_05350_));
 OA211x2_ASAP7_75t_R _23020_ (.A1(net346),
    .A2(_05349_),
    .B(_05350_),
    .C(net369),
    .Y(_05351_));
 OR3x1_ASAP7_75t_R _23021_ (.A(net337),
    .B(_05348_),
    .C(_05351_),
    .Y(_05352_));
 AND3x1_ASAP7_75t_R _23022_ (.A(_13373_),
    .B(_05345_),
    .C(_05352_),
    .Y(_05353_));
 OR3x4_ASAP7_75t_R _23023_ (.A(net328),
    .B(_05338_),
    .C(_05353_),
    .Y(_05354_));
 NAND2x2_ASAP7_75t_R _23024_ (.A(_05323_),
    .B(_05354_),
    .Y(_05355_));
 OA21x2_ASAP7_75t_R _23025_ (.A1(_01739_),
    .A2(_15489_),
    .B(_16459_),
    .Y(_05356_));
 AO21x2_ASAP7_75t_R _23026_ (.A1(_13474_),
    .A2(_05355_),
    .B(_05356_),
    .Y(_05357_));
 TAPCELL_ASAP7_75t_R TAP_1068 ();
 INVx1_ASAP7_75t_R _23028_ (.A(_05357_),
    .Y(_18475_));
 NAND2x1_ASAP7_75t_R _23029_ (.A(net413),
    .B(_01263_),
    .Y(_05358_));
 OA211x2_ASAP7_75t_R _23030_ (.A1(net413),
    .A2(_05324_),
    .B(_05358_),
    .C(net319),
    .Y(_05359_));
 NAND2x1_ASAP7_75t_R _23031_ (.A(net413),
    .B(_01262_),
    .Y(_05360_));
 OA211x2_ASAP7_75t_R _23032_ (.A1(net413),
    .A2(_05327_),
    .B(_05360_),
    .C(net426),
    .Y(_05361_));
 OR3x1_ASAP7_75t_R _23033_ (.A(_14015_),
    .B(_05359_),
    .C(_05361_),
    .Y(_05362_));
 NAND2x1_ASAP7_75t_R _23034_ (.A(net413),
    .B(_01259_),
    .Y(_05363_));
 OA211x2_ASAP7_75t_R _23035_ (.A1(net413),
    .A2(_05331_),
    .B(_05363_),
    .C(net319),
    .Y(_05364_));
 NAND2x1_ASAP7_75t_R _23036_ (.A(net413),
    .B(_01258_),
    .Y(_05365_));
 OA211x2_ASAP7_75t_R _23037_ (.A1(net413),
    .A2(_05334_),
    .B(_05365_),
    .C(net426),
    .Y(_05366_));
 OR3x1_ASAP7_75t_R _23038_ (.A(net315),
    .B(_05364_),
    .C(_05366_),
    .Y(_05367_));
 NAND2x1_ASAP7_75t_R _23039_ (.A(net415),
    .B(_01246_),
    .Y(_05368_));
 OA211x2_ASAP7_75t_R _23040_ (.A1(net415),
    .A2(_05311_),
    .B(_05368_),
    .C(net426),
    .Y(_05369_));
 NAND2x1_ASAP7_75t_R _23041_ (.A(net415),
    .B(_01247_),
    .Y(_05370_));
 OA211x2_ASAP7_75t_R _23042_ (.A1(net415),
    .A2(_05308_),
    .B(_05370_),
    .C(net319),
    .Y(_05371_));
 OR3x1_ASAP7_75t_R _23043_ (.A(_14015_),
    .B(_05369_),
    .C(_05371_),
    .Y(_05372_));
 NAND2x1_ASAP7_75t_R _23044_ (.A(net415),
    .B(_01679_),
    .Y(_05373_));
 OA211x2_ASAP7_75t_R _23045_ (.A1(net415),
    .A2(_05303_),
    .B(_05373_),
    .C(net318),
    .Y(_05374_));
 AND3x1_ASAP7_75t_R _23046_ (.A(net426),
    .B(net316),
    .C(_05302_),
    .Y(_05375_));
 OA31x2_ASAP7_75t_R _23047_ (.A1(net315),
    .A2(_05374_),
    .A3(_05375_),
    .B1(net378),
    .Y(_05376_));
 AO32x1_ASAP7_75t_R _23048_ (.A1(_13626_),
    .A2(_05362_),
    .A3(_05367_),
    .B1(_05372_),
    .B2(_05376_),
    .Y(_05377_));
 NAND2x1_ASAP7_75t_R _23049_ (.A(net412),
    .B(_01267_),
    .Y(_05378_));
 OA211x2_ASAP7_75t_R _23050_ (.A1(net412),
    .A2(_05339_),
    .B(_05378_),
    .C(net319),
    .Y(_05379_));
 NAND2x1_ASAP7_75t_R _23051_ (.A(net412),
    .B(_01266_),
    .Y(_05380_));
 OA211x2_ASAP7_75t_R _23052_ (.A1(net412),
    .A2(_05342_),
    .B(_05380_),
    .C(net426),
    .Y(_05381_));
 OR3x1_ASAP7_75t_R _23053_ (.A(net321),
    .B(_05379_),
    .C(_05381_),
    .Y(_05382_));
 NAND2x1_ASAP7_75t_R _23054_ (.A(net415),
    .B(_01271_),
    .Y(_05383_));
 OA211x2_ASAP7_75t_R _23055_ (.A1(net415),
    .A2(_05346_),
    .B(_05383_),
    .C(net319),
    .Y(_05384_));
 NAND2x1_ASAP7_75t_R _23056_ (.A(net415),
    .B(_01270_),
    .Y(_05385_));
 OA211x2_ASAP7_75t_R _23057_ (.A1(net415),
    .A2(_05349_),
    .B(_05385_),
    .C(net426),
    .Y(_05386_));
 OR3x1_ASAP7_75t_R _23058_ (.A(net387),
    .B(_05384_),
    .C(_05386_),
    .Y(_05387_));
 AND5x1_ASAP7_75t_R _23059_ (.A(_13626_),
    .B(_05362_),
    .C(_05367_),
    .D(_05382_),
    .E(_05387_),
    .Y(_05388_));
 NAND2x1_ASAP7_75t_R _23060_ (.A(net415),
    .B(_01251_),
    .Y(_05389_));
 OA211x2_ASAP7_75t_R _23061_ (.A1(net415),
    .A2(_05295_),
    .B(_05389_),
    .C(net319),
    .Y(_05390_));
 NAND2x1_ASAP7_75t_R _23062_ (.A(net415),
    .B(_01250_),
    .Y(_05391_));
 OA211x2_ASAP7_75t_R _23063_ (.A1(net415),
    .A2(_05298_),
    .B(_05391_),
    .C(net426),
    .Y(_05392_));
 OR3x1_ASAP7_75t_R _23064_ (.A(net321),
    .B(_05390_),
    .C(_05392_),
    .Y(_05393_));
 NAND2x1_ASAP7_75t_R _23065_ (.A(net415),
    .B(_01255_),
    .Y(_05394_));
 OA211x2_ASAP7_75t_R _23066_ (.A1(net415),
    .A2(_05315_),
    .B(_05394_),
    .C(net319),
    .Y(_05395_));
 NAND2x1_ASAP7_75t_R _23067_ (.A(net415),
    .B(_01254_),
    .Y(_05396_));
 OA211x2_ASAP7_75t_R _23068_ (.A1(net415),
    .A2(_05318_),
    .B(_05396_),
    .C(net426),
    .Y(_05397_));
 OR3x1_ASAP7_75t_R _23069_ (.A(net387),
    .B(_05395_),
    .C(_05397_),
    .Y(_05398_));
 AND4x1_ASAP7_75t_R _23070_ (.A(_05372_),
    .B(_05376_),
    .C(_05393_),
    .D(_05398_),
    .Y(_05399_));
 AO211x2_ASAP7_75t_R _23071_ (.A1(net382),
    .A2(_05377_),
    .B(_05388_),
    .C(_05399_),
    .Y(_05400_));
 INVx2_ASAP7_75t_R _23072_ (.A(_00229_),
    .Y(_05401_));
 INVx1_ASAP7_75t_R _23073_ (.A(_01611_),
    .Y(_05402_));
 AO32x2_ASAP7_75t_R _23074_ (.A1(_05401_),
    .A2(_13993_),
    .A3(_13794_),
    .B1(_05402_),
    .B2(_13450_),
    .Y(_05403_));
 AOI21x1_ASAP7_75t_R _23075_ (.A1(_13810_),
    .A2(_05400_),
    .B(_05403_),
    .Y(_18474_));
 XNOR2x2_ASAP7_75t_R _23076_ (.A(_01277_),
    .B(_01275_),
    .Y(_05404_));
 INVx4_ASAP7_75t_R _23077_ (.A(_05404_),
    .Y(net172));
 INVx1_ASAP7_75t_R _23078_ (.A(_01295_),
    .Y(_05405_));
 NAND2x1_ASAP7_75t_R _23079_ (.A(net2248),
    .B(_01293_),
    .Y(_05406_));
 OA211x2_ASAP7_75t_R _23080_ (.A1(net2249),
    .A2(_05405_),
    .B(_05406_),
    .C(net323),
    .Y(_05407_));
 INVx1_ASAP7_75t_R _23081_ (.A(_01294_),
    .Y(_05408_));
 NAND2x1_ASAP7_75t_R _23082_ (.A(net2276),
    .B(_01292_),
    .Y(_05409_));
 OA211x2_ASAP7_75t_R _23083_ (.A1(net2277),
    .A2(_05408_),
    .B(_05409_),
    .C(net375),
    .Y(_05410_));
 OR3x1_ASAP7_75t_R _23084_ (.A(_13350_),
    .B(_05407_),
    .C(_05410_),
    .Y(_05411_));
 AND2x2_ASAP7_75t_R _23085_ (.A(net2276),
    .B(_01297_),
    .Y(_05412_));
 AO21x1_ASAP7_75t_R _23086_ (.A1(net326),
    .A2(_01299_),
    .B(_05412_),
    .Y(_05413_));
 AND2x2_ASAP7_75t_R _23087_ (.A(net2269),
    .B(_01296_),
    .Y(_05414_));
 AO21x1_ASAP7_75t_R _23088_ (.A1(net2278),
    .A2(_01298_),
    .B(_05414_),
    .Y(_05415_));
 AOI221x1_ASAP7_75t_R _23089_ (.A1(_13402_),
    .A2(_05413_),
    .B1(_05415_),
    .B2(_13366_),
    .C(_14275_),
    .Y(_05416_));
 INVx1_ASAP7_75t_R _23090_ (.A(_01291_),
    .Y(_05417_));
 NAND2x1_ASAP7_75t_R _23091_ (.A(net366),
    .B(_01289_),
    .Y(_05418_));
 OA211x2_ASAP7_75t_R _23092_ (.A1(net2277),
    .A2(_05417_),
    .B(_13402_),
    .C(_05418_),
    .Y(_05419_));
 INVx1_ASAP7_75t_R _23093_ (.A(_01288_),
    .Y(_05420_));
 NAND2x1_ASAP7_75t_R _23094_ (.A(net326),
    .B(_01290_),
    .Y(_05421_));
 OA211x2_ASAP7_75t_R _23095_ (.A1(net326),
    .A2(_05420_),
    .B(_13366_),
    .C(_05421_),
    .Y(_05422_));
 INVx1_ASAP7_75t_R _23096_ (.A(_01287_),
    .Y(_05423_));
 NAND2x1_ASAP7_75t_R _23097_ (.A(net366),
    .B(_01285_),
    .Y(_05424_));
 OA211x2_ASAP7_75t_R _23098_ (.A1(net2336),
    .A2(_05423_),
    .B(_13377_),
    .C(_05424_),
    .Y(_05425_));
 INVx1_ASAP7_75t_R _23099_ (.A(_01286_),
    .Y(_05426_));
 NAND2x1_ASAP7_75t_R _23100_ (.A(net366),
    .B(_01284_),
    .Y(_05427_));
 OA211x2_ASAP7_75t_R _23101_ (.A1(net2336),
    .A2(_05426_),
    .B(_13357_),
    .C(_05427_),
    .Y(_05428_));
 OR5x1_ASAP7_75t_R _23102_ (.A(net329),
    .B(_05419_),
    .C(_05422_),
    .D(_05425_),
    .E(_05428_),
    .Y(_05429_));
 AND2x2_ASAP7_75t_R _23103_ (.A(net367),
    .B(_01678_),
    .Y(_05430_));
 AO21x1_ASAP7_75t_R _23104_ (.A1(net326),
    .A2(_01279_),
    .B(_05430_),
    .Y(_05431_));
 OAI22x1_ASAP7_75t_R _23105_ (.A1(_01278_),
    .A2(net311),
    .B1(_05431_),
    .B2(net375),
    .Y(_05432_));
 INVx1_ASAP7_75t_R _23106_ (.A(_01282_),
    .Y(_05433_));
 NAND2x1_ASAP7_75t_R _23107_ (.A(net365),
    .B(_01280_),
    .Y(_05434_));
 OA211x2_ASAP7_75t_R _23108_ (.A1(net2269),
    .A2(_05433_),
    .B(_05434_),
    .C(net374),
    .Y(_05435_));
 INVx1_ASAP7_75t_R _23109_ (.A(_01283_),
    .Y(_05436_));
 NAND2x1_ASAP7_75t_R _23110_ (.A(net366),
    .B(_01281_),
    .Y(_05437_));
 OA211x2_ASAP7_75t_R _23111_ (.A1(net2336),
    .A2(_05436_),
    .B(_05437_),
    .C(net323),
    .Y(_05438_));
 OR3x1_ASAP7_75t_R _23112_ (.A(_14383_),
    .B(_05435_),
    .C(_05438_),
    .Y(_05439_));
 OA211x2_ASAP7_75t_R _23113_ (.A1(_13851_),
    .A2(_05432_),
    .B(_05439_),
    .C(net328),
    .Y(_05440_));
 INVx1_ASAP7_75t_R _23114_ (.A(_01307_),
    .Y(_05441_));
 NAND2x1_ASAP7_75t_R _23115_ (.A(net2249),
    .B(_01305_),
    .Y(_05442_));
 OA211x2_ASAP7_75t_R _23116_ (.A1(net367),
    .A2(_05441_),
    .B(_05442_),
    .C(net323),
    .Y(_05443_));
 INVx1_ASAP7_75t_R _23117_ (.A(_01306_),
    .Y(_05444_));
 NAND2x1_ASAP7_75t_R _23118_ (.A(net366),
    .B(_01304_),
    .Y(_05445_));
 OA211x2_ASAP7_75t_R _23119_ (.A1(net2336),
    .A2(_05444_),
    .B(_05445_),
    .C(net375),
    .Y(_05446_));
 OR3x1_ASAP7_75t_R _23120_ (.A(net2360),
    .B(_05443_),
    .C(_05446_),
    .Y(_05447_));
 AND2x2_ASAP7_75t_R _23121_ (.A(net2249),
    .B(_01301_),
    .Y(_05448_));
 AO21x1_ASAP7_75t_R _23122_ (.A1(net326),
    .A2(_01303_),
    .B(_05448_),
    .Y(_05449_));
 AND2x2_ASAP7_75t_R _23123_ (.A(net2249),
    .B(_01300_),
    .Y(_05450_));
 AO21x1_ASAP7_75t_R _23124_ (.A1(net326),
    .A2(_01302_),
    .B(_05450_),
    .Y(_05451_));
 AOI22x1_ASAP7_75t_R _23125_ (.A1(_13377_),
    .A2(_05449_),
    .B1(_05451_),
    .B2(_13357_),
    .Y(_05452_));
 AND3x1_ASAP7_75t_R _23126_ (.A(_13439_),
    .B(_05447_),
    .C(_05452_),
    .Y(_05453_));
 AO221x2_ASAP7_75t_R _23127_ (.A1(_05411_),
    .A2(_05416_),
    .B1(_05429_),
    .B2(_05440_),
    .C(_05453_),
    .Y(_05454_));
 OA211x2_ASAP7_75t_R _23128_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14704_),
    .C(_13521_),
    .Y(_05455_));
 AOI21x1_ASAP7_75t_R _23129_ (.A1(_13474_),
    .A2(_05454_),
    .B(_05455_),
    .Y(_17804_));
 INVx1_ASAP7_75t_R _23130_ (.A(_17804_),
    .Y(_17806_));
 AO21x2_ASAP7_75t_R _23131_ (.A1(_13445_),
    .A2(_13449_),
    .B(_01610_),
    .Y(_05456_));
 AOI22x1_ASAP7_75t_R _23132_ (.A1(_00230_),
    .A2(_13993_),
    .B1(_14988_),
    .B2(_05456_),
    .Y(_05457_));
 NAND2x1_ASAP7_75t_R _23133_ (.A(net386),
    .B(_01287_),
    .Y(_05458_));
 OA211x2_ASAP7_75t_R _23134_ (.A1(net386),
    .A2(_05417_),
    .B(_05458_),
    .C(net316),
    .Y(_05459_));
 INVx1_ASAP7_75t_R _23135_ (.A(_01289_),
    .Y(_05460_));
 NAND2x1_ASAP7_75t_R _23136_ (.A(net2301),
    .B(_01285_),
    .Y(_05461_));
 OA211x2_ASAP7_75t_R _23137_ (.A1(net386),
    .A2(_05460_),
    .B(_05461_),
    .C(net414),
    .Y(_05462_));
 OA21x2_ASAP7_75t_R _23138_ (.A1(_05459_),
    .A2(_05462_),
    .B(net319),
    .Y(_05463_));
 INVx1_ASAP7_75t_R _23139_ (.A(_01284_),
    .Y(_05464_));
 NOR2x1_ASAP7_75t_R _23140_ (.A(net2379),
    .B(_01286_),
    .Y(_05465_));
 AO21x1_ASAP7_75t_R _23141_ (.A1(net411),
    .A2(_05464_),
    .B(_05465_),
    .Y(_05466_));
 AND2x2_ASAP7_75t_R _23142_ (.A(net425),
    .B(net386),
    .Y(_05467_));
 AND2x2_ASAP7_75t_R _23143_ (.A(net425),
    .B(net321),
    .Y(_05468_));
 INVx1_ASAP7_75t_R _23144_ (.A(_01290_),
    .Y(_05469_));
 NAND2x1_ASAP7_75t_R _23145_ (.A(net2379),
    .B(_01288_),
    .Y(_05470_));
 OA21x2_ASAP7_75t_R _23146_ (.A1(net411),
    .A2(_05469_),
    .B(_05470_),
    .Y(_05471_));
 AO221x1_ASAP7_75t_R _23147_ (.A1(_05466_),
    .A2(_05467_),
    .B1(_05468_),
    .B2(_05471_),
    .C(net380),
    .Y(_05472_));
 NAND2x1_ASAP7_75t_R _23148_ (.A(net2379),
    .B(_01280_),
    .Y(_05473_));
 OA211x2_ASAP7_75t_R _23149_ (.A1(net411),
    .A2(_05433_),
    .B(_05473_),
    .C(net425),
    .Y(_05474_));
 NAND2x1_ASAP7_75t_R _23150_ (.A(net414),
    .B(_01281_),
    .Y(_05475_));
 OA211x2_ASAP7_75t_R _23151_ (.A1(net414),
    .A2(_05436_),
    .B(_05475_),
    .C(net319),
    .Y(_05476_));
 OR3x1_ASAP7_75t_R _23152_ (.A(_14015_),
    .B(_05474_),
    .C(_05476_),
    .Y(_05477_));
 INVx1_ASAP7_75t_R _23153_ (.A(_01279_),
    .Y(_05478_));
 NAND2x1_ASAP7_75t_R _23154_ (.A(net425),
    .B(_01278_),
    .Y(_05479_));
 OA211x2_ASAP7_75t_R _23155_ (.A1(net425),
    .A2(_05478_),
    .B(_05479_),
    .C(net316),
    .Y(_05480_));
 INVx1_ASAP7_75t_R _23156_ (.A(_01678_),
    .Y(_05481_));
 AND3x1_ASAP7_75t_R _23157_ (.A(net319),
    .B(net414),
    .C(_05481_),
    .Y(_05482_));
 OA31x2_ASAP7_75t_R _23158_ (.A1(net315),
    .A2(_05480_),
    .A3(_05482_),
    .B1(net378),
    .Y(_05483_));
 OA211x2_ASAP7_75t_R _23159_ (.A1(_05463_),
    .A2(_05472_),
    .B(_05477_),
    .C(_05483_),
    .Y(_05484_));
 AND2x2_ASAP7_75t_R _23160_ (.A(net410),
    .B(_01296_),
    .Y(_05485_));
 AO21x1_ASAP7_75t_R _23161_ (.A1(net316),
    .A2(_01298_),
    .B(_05485_),
    .Y(_05486_));
 AND2x2_ASAP7_75t_R _23162_ (.A(net410),
    .B(_01297_),
    .Y(_05487_));
 AO21x1_ASAP7_75t_R _23163_ (.A1(net316),
    .A2(_01299_),
    .B(_05487_),
    .Y(_05488_));
 NOR2x1_ASAP7_75t_R _23164_ (.A(net425),
    .B(net386),
    .Y(_05489_));
 AOI22x1_ASAP7_75t_R _23165_ (.A1(_05468_),
    .A2(_05486_),
    .B1(_05488_),
    .B2(_05489_),
    .Y(_05490_));
 NAND2x1_ASAP7_75t_R _23166_ (.A(net414),
    .B(_01293_),
    .Y(_05491_));
 OA21x2_ASAP7_75t_R _23167_ (.A1(net414),
    .A2(_05405_),
    .B(_05491_),
    .Y(_05492_));
 OR3x1_ASAP7_75t_R _23168_ (.A(net425),
    .B(net321),
    .C(_05492_),
    .Y(_05493_));
 AND2x2_ASAP7_75t_R _23169_ (.A(net414),
    .B(_01292_),
    .Y(_05494_));
 AO21x1_ASAP7_75t_R _23170_ (.A1(net316),
    .A2(_01294_),
    .B(_05494_),
    .Y(_05495_));
 NAND2x1_ASAP7_75t_R _23171_ (.A(_05467_),
    .B(_05495_),
    .Y(_05496_));
 AND5x1_ASAP7_75t_R _23172_ (.A(net380),
    .B(_13626_),
    .C(_05490_),
    .D(_05493_),
    .E(_05496_),
    .Y(_05497_));
 INVx1_ASAP7_75t_R _23173_ (.A(_01303_),
    .Y(_05498_));
 NAND2x1_ASAP7_75t_R _23174_ (.A(net414),
    .B(_01301_),
    .Y(_05499_));
 OA211x2_ASAP7_75t_R _23175_ (.A1(net414),
    .A2(_05498_),
    .B(_05499_),
    .C(net319),
    .Y(_05500_));
 INVx1_ASAP7_75t_R _23176_ (.A(_01302_),
    .Y(_05501_));
 NAND2x1_ASAP7_75t_R _23177_ (.A(net414),
    .B(_01300_),
    .Y(_05502_));
 OA211x2_ASAP7_75t_R _23178_ (.A1(net414),
    .A2(_05501_),
    .B(_05502_),
    .C(net425),
    .Y(_05503_));
 OR3x1_ASAP7_75t_R _23179_ (.A(net321),
    .B(_05500_),
    .C(_05503_),
    .Y(_05504_));
 NAND2x1_ASAP7_75t_R _23180_ (.A(net414),
    .B(_01305_),
    .Y(_05505_));
 OA211x2_ASAP7_75t_R _23181_ (.A1(net414),
    .A2(_05441_),
    .B(_05505_),
    .C(net319),
    .Y(_05506_));
 NAND2x1_ASAP7_75t_R _23182_ (.A(net414),
    .B(_01304_),
    .Y(_05507_));
 OA211x2_ASAP7_75t_R _23183_ (.A1(net414),
    .A2(_05444_),
    .B(_05507_),
    .C(net425),
    .Y(_05508_));
 OR3x1_ASAP7_75t_R _23184_ (.A(net2304),
    .B(_05506_),
    .C(_05508_),
    .Y(_05509_));
 AND3x1_ASAP7_75t_R _23185_ (.A(_14780_),
    .B(_05504_),
    .C(_05509_),
    .Y(_05510_));
 OR5x2_ASAP7_75t_R _23186_ (.A(_13993_),
    .B(_14988_),
    .C(_05484_),
    .D(_05497_),
    .E(_05510_),
    .Y(_05511_));
 AND2x6_ASAP7_75t_R _23187_ (.A(_05457_),
    .B(_05511_),
    .Y(_17807_));
 INVx2_ASAP7_75t_R _23188_ (.A(_17807_),
    .Y(_17805_));
 NOR2x2_ASAP7_75t_R _23189_ (.A(_13620_),
    .B(_17804_),
    .Y(_05512_));
 OR3x4_ASAP7_75t_R _23190_ (.A(_05484_),
    .B(_05497_),
    .C(_05510_),
    .Y(_05513_));
 OR2x2_ASAP7_75t_R _23191_ (.A(_00284_),
    .B(_05513_),
    .Y(_05514_));
 AO221x1_ASAP7_75t_R _23192_ (.A1(_13775_),
    .A2(_01308_),
    .B1(_02202_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_05515_));
 NOR2x1_ASAP7_75t_R _23193_ (.A(_13538_),
    .B(_05515_),
    .Y(_05516_));
 TAPCELL_ASAP7_75t_R TAP_1067 ();
 AND3x1_ASAP7_75t_R _23195_ (.A(_13817_),
    .B(_13772_),
    .C(_05454_),
    .Y(_05518_));
 AO221x2_ASAP7_75t_R _23196_ (.A1(_14002_),
    .A2(_17804_),
    .B1(_05514_),
    .B2(_05516_),
    .C(_05518_),
    .Y(_05519_));
 OA21x2_ASAP7_75t_R _23197_ (.A1(_01078_),
    .A2(_01079_),
    .B(_02279_),
    .Y(_05520_));
 OA21x2_ASAP7_75t_R _23198_ (.A1(_01111_),
    .A2(_05520_),
    .B(_01144_),
    .Y(_05521_));
 OA21x2_ASAP7_75t_R _23199_ (.A1(_01143_),
    .A2(_05521_),
    .B(_02280_),
    .Y(_05522_));
 OR4x1_ASAP7_75t_R _23200_ (.A(_01078_),
    .B(_01046_),
    .C(_01143_),
    .D(_01111_),
    .Y(_05523_));
 OR4x1_ASAP7_75t_R _23201_ (.A(_01209_),
    .B(_01177_),
    .C(_01275_),
    .D(_01243_),
    .Y(_05524_));
 AND3x1_ASAP7_75t_R _23202_ (.A(_04634_),
    .B(_04637_),
    .C(_05522_),
    .Y(_05525_));
 AOI211x1_ASAP7_75t_R _23203_ (.A1(_05522_),
    .A2(_05523_),
    .B(_05524_),
    .C(_05525_),
    .Y(_05526_));
 OR3x1_ASAP7_75t_R _23204_ (.A(_00719_),
    .B(_15656_),
    .C(_16388_),
    .Y(_05527_));
 OR4x1_ASAP7_75t_R _23205_ (.A(_00719_),
    .B(_15343_),
    .C(_15652_),
    .D(_16388_),
    .Y(_05528_));
 AO21x1_ASAP7_75t_R _23206_ (.A1(_16727_),
    .A2(_15227_),
    .B(_05528_),
    .Y(_05529_));
 AND3x1_ASAP7_75t_R _23207_ (.A(_16392_),
    .B(_04637_),
    .C(_05522_),
    .Y(_05530_));
 NAND3x1_ASAP7_75t_R _23208_ (.A(_05527_),
    .B(_05529_),
    .C(_05530_),
    .Y(_05531_));
 OA21x2_ASAP7_75t_R _23209_ (.A1(_01209_),
    .A2(_01210_),
    .B(_02281_),
    .Y(_05532_));
 OA21x2_ASAP7_75t_R _23210_ (.A1(_01243_),
    .A2(_05532_),
    .B(_01276_),
    .Y(_05533_));
 OAI21x1_ASAP7_75t_R _23211_ (.A1(_01275_),
    .A2(_05533_),
    .B(_01309_),
    .Y(_05534_));
 AO21x1_ASAP7_75t_R _23212_ (.A1(_05526_),
    .A2(_05531_),
    .B(_05534_),
    .Y(_05535_));
 INVx3_ASAP7_75t_R _23213_ (.A(_01308_),
    .Y(_05536_));
 AOI221x1_ASAP7_75t_R _23214_ (.A1(_00230_),
    .A2(_13993_),
    .B1(_14988_),
    .B2(_05456_),
    .C(_13817_),
    .Y(_05537_));
 AO32x1_ASAP7_75t_R _23215_ (.A1(_05536_),
    .A2(_13817_),
    .A3(_13778_),
    .B1(_05511_),
    .B2(_05537_),
    .Y(_05538_));
 XNOR2x2_ASAP7_75t_R _23216_ (.A(_05535_),
    .B(_05538_),
    .Y(_05539_));
 OA21x2_ASAP7_75t_R _23217_ (.A1(_05512_),
    .A2(_05519_),
    .B(_05539_),
    .Y(_05540_));
 NOR3x2_ASAP7_75t_R _23218_ (.B(_05519_),
    .C(_05539_),
    .Y(_05541_),
    .A(_05512_));
 OR2x6_ASAP7_75t_R _23219_ (.A(_05540_),
    .B(_05541_),
    .Y(_05542_));
 TAPCELL_ASAP7_75t_R TAP_1066 ();
 CKINVDCx5p33_ASAP7_75t_R _23221_ (.A(_05542_),
    .Y(net173));
 TAPCELL_ASAP7_75t_R TAP_1065 ();
 INVx1_ASAP7_75t_R _23223_ (.A(_02140_),
    .Y(\cs_registers_i.priv_lvl_q[0] ));
 INVx2_ASAP7_75t_R _23224_ (.A(_13534_),
    .Y(_05545_));
 AND3x4_ASAP7_75t_R _23225_ (.A(_00279_),
    .B(_00281_),
    .C(_00282_),
    .Y(_05546_));
 AO21x2_ASAP7_75t_R _23226_ (.A1(_14362_),
    .A2(_13574_),
    .B(_13612_),
    .Y(_05547_));
 OR4x2_ASAP7_75t_R _23227_ (.A(_01874_),
    .B(_05545_),
    .C(_05546_),
    .D(_05547_),
    .Y(_05548_));
 TAPCELL_ASAP7_75t_R TAP_1064 ();
 AND3x1_ASAP7_75t_R _23229_ (.A(_00279_),
    .B(_14843_),
    .C(_05548_),
    .Y(_05550_));
 AOI21x1_ASAP7_75t_R _23230_ (.A1(_01314_),
    .A2(_14845_),
    .B(_05550_),
    .Y(_00001_));
 INVx1_ASAP7_75t_R _23231_ (.A(net3036),
    .Y(_05551_));
 AND3x4_ASAP7_75t_R _23232_ (.A(_00277_),
    .B(_01608_),
    .C(_01609_),
    .Y(_05552_));
 NAND2x2_ASAP7_75t_R _23233_ (.A(net3055),
    .B(_05552_),
    .Y(_05553_));
 AO21x2_ASAP7_75t_R _23234_ (.A1(net3037),
    .A2(_01607_),
    .B(net3056),
    .Y(_05554_));
 NOR2x1_ASAP7_75t_R _23235_ (.A(_01316_),
    .B(net3058),
    .Y(\id_stage_i.controller_i.store_err_d ));
 INVx1_ASAP7_75t_R _23236_ (.A(_01316_),
    .Y(_05555_));
 NOR2x1_ASAP7_75t_R _23237_ (.A(_05555_),
    .B(net3058),
    .Y(\id_stage_i.controller_i.load_err_d ));
 INVx2_ASAP7_75t_R _23238_ (.A(_01716_),
    .Y(_05556_));
 AND4x2_ASAP7_75t_R _23239_ (.A(_01714_),
    .B(_14793_),
    .C(_05556_),
    .D(_01717_),
    .Y(_05557_));
 TAPCELL_ASAP7_75t_R TAP_1063 ();
 TAPCELL_ASAP7_75t_R TAP_1062 ();
 TAPCELL_ASAP7_75t_R TAP_1061 ();
 TAPCELL_ASAP7_75t_R TAP_1060 ();
 OR5x2_ASAP7_75t_R _23244_ (.A(_00172_),
    .B(_14837_),
    .C(_13470_),
    .D(_13463_),
    .E(_05546_),
    .Y(_05562_));
 AO21x2_ASAP7_75t_R _23245_ (.A1(_14812_),
    .A2(_14836_),
    .B(_05562_),
    .Y(_05563_));
 AOI21x1_ASAP7_75t_R _23246_ (.A1(_13495_),
    .A2(_14236_),
    .B(_05563_),
    .Y(_05564_));
 TAPCELL_ASAP7_75t_R TAP_1059 ();
 AND2x2_ASAP7_75t_R _23248_ (.A(_14297_),
    .B(_05564_),
    .Y(_05566_));
 NOR2x2_ASAP7_75t_R _23249_ (.A(_14394_),
    .B(_14419_),
    .Y(_05567_));
 AO33x2_ASAP7_75t_R _23250_ (.A1(_00283_),
    .A2(_14423_),
    .A3(_14424_),
    .B1(_05567_),
    .B2(_14479_),
    .B3(_13474_),
    .Y(_05568_));
 TAPCELL_ASAP7_75t_R TAP_1058 ();
 AOI21x1_ASAP7_75t_R _23252_ (.A1(_14812_),
    .A2(_14836_),
    .B(_05562_),
    .Y(_05570_));
 NOR2x2_ASAP7_75t_R _23253_ (.A(_01740_),
    .B(_01741_),
    .Y(_05571_));
 AND2x4_ASAP7_75t_R _23254_ (.A(_01739_),
    .B(_05571_),
    .Y(_05572_));
 AND2x2_ASAP7_75t_R _23255_ (.A(_05570_),
    .B(_05572_),
    .Y(_05573_));
 AND4x1_ASAP7_75t_R _23256_ (.A(_13528_),
    .B(_14424_),
    .C(_14710_),
    .D(_05573_),
    .Y(_05574_));
 AND3x1_ASAP7_75t_R _23257_ (.A(_05566_),
    .B(_05568_),
    .C(_05574_),
    .Y(_05575_));
 OR3x1_ASAP7_75t_R _23258_ (.A(_01317_),
    .B(_13804_),
    .C(_05575_),
    .Y(_05576_));
 TAPCELL_ASAP7_75t_R TAP_1057 ();
 TAPCELL_ASAP7_75t_R TAP_1056 ();
 TAPCELL_ASAP7_75t_R TAP_1055 ();
 TAPCELL_ASAP7_75t_R TAP_1054 ();
 OA21x2_ASAP7_75t_R _23263_ (.A1(_14179_),
    .A2(_14239_),
    .B(_05570_),
    .Y(_05581_));
 AND2x2_ASAP7_75t_R _23264_ (.A(_13528_),
    .B(_05570_),
    .Y(_05582_));
 OA211x2_ASAP7_75t_R _23265_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14356_),
    .C(_05582_),
    .Y(_05583_));
 OA21x2_ASAP7_75t_R _23266_ (.A1(_14295_),
    .A2(_14294_),
    .B(_05583_),
    .Y(_05584_));
 AND3x1_ASAP7_75t_R _23267_ (.A(_13595_),
    .B(_05571_),
    .C(_05570_),
    .Y(_05585_));
 OA211x2_ASAP7_75t_R _23268_ (.A1(_13495_),
    .A2(_13888_),
    .B(_05585_),
    .C(_13481_),
    .Y(_05586_));
 TAPCELL_ASAP7_75t_R TAP_1053 ();
 OA211x2_ASAP7_75t_R _23270_ (.A1(_13521_),
    .A2(_14703_),
    .B(_05586_),
    .C(_14709_),
    .Y(_05588_));
 NAND3x2_ASAP7_75t_R _23271_ (.B(_05584_),
    .C(_05588_),
    .Y(_05589_),
    .A(_05568_));
 OR3x1_ASAP7_75t_R _23272_ (.A(_01311_),
    .B(_05581_),
    .C(_05589_),
    .Y(_05590_));
 INVx1_ASAP7_75t_R _23273_ (.A(_05590_),
    .Y(_05591_));
 TAPCELL_ASAP7_75t_R TAP_1052 ();
 AND2x2_ASAP7_75t_R _23275_ (.A(_14239_),
    .B(net310),
    .Y(_05593_));
 NAND2x2_ASAP7_75t_R _23276_ (.A(_00283_),
    .B(_01742_),
    .Y(_05594_));
 OR4x2_ASAP7_75t_R _23277_ (.A(_14394_),
    .B(_14419_),
    .C(_14452_),
    .D(_14478_),
    .Y(_05595_));
 AOI22x1_ASAP7_75t_R _23278_ (.A1(_05594_),
    .A2(_14424_),
    .B1(_05595_),
    .B2(_13474_),
    .Y(_05596_));
 TAPCELL_ASAP7_75t_R TAP_1051 ();
 AO32x2_ASAP7_75t_R _23280_ (.A1(net323),
    .A2(_13495_),
    .A3(_13505_),
    .B1(_14706_),
    .B2(_14707_),
    .Y(_05598_));
 TAPCELL_ASAP7_75t_R TAP_1050 ();
 NAND2x2_ASAP7_75t_R _23282_ (.A(_05570_),
    .B(_05572_),
    .Y(_05600_));
 NOR3x2_ASAP7_75t_R _23283_ (.B(_05598_),
    .C(_05600_),
    .Y(_05601_),
    .A(_14543_));
 AND2x4_ASAP7_75t_R _23284_ (.A(_05596_),
    .B(_05601_),
    .Y(_05602_));
 AND3x1_ASAP7_75t_R _23285_ (.A(_05593_),
    .B(_05584_),
    .C(_05602_),
    .Y(_05603_));
 AND3x2_ASAP7_75t_R _23286_ (.A(_14358_),
    .B(_05596_),
    .C(_05601_),
    .Y(_05604_));
 OR3x1_ASAP7_75t_R _23287_ (.A(_00323_),
    .B(_14542_),
    .C(_13512_),
    .Y(_05605_));
 OR3x1_ASAP7_75t_R _23288_ (.A(net375),
    .B(_13450_),
    .C(_13505_),
    .Y(_05606_));
 AO21x1_ASAP7_75t_R _23289_ (.A1(net2277),
    .A2(_05606_),
    .B(_13520_),
    .Y(_05607_));
 AND4x2_ASAP7_75t_R _23290_ (.A(_13521_),
    .B(_13514_),
    .C(_05605_),
    .D(_05607_),
    .Y(_05608_));
 TAPCELL_ASAP7_75t_R TAP_1049 ();
 AND2x2_ASAP7_75t_R _23292_ (.A(_14180_),
    .B(_05608_),
    .Y(_05610_));
 AO33x2_ASAP7_75t_R _23293_ (.A1(net305),
    .A2(_14179_),
    .A3(_05603_),
    .B1(_05604_),
    .B2(_05610_),
    .B3(_05566_),
    .Y(_05611_));
 AND2x2_ASAP7_75t_R _23294_ (.A(_13523_),
    .B(_13894_),
    .Y(_05612_));
 AND3x1_ASAP7_75t_R _23295_ (.A(_14296_),
    .B(_14359_),
    .C(_05596_),
    .Y(_05613_));
 AND3x1_ASAP7_75t_R _23296_ (.A(net310),
    .B(_05612_),
    .C(_05613_),
    .Y(_05614_));
 AND3x1_ASAP7_75t_R _23297_ (.A(_14179_),
    .B(_05564_),
    .C(_05601_),
    .Y(_05615_));
 AND3x4_ASAP7_75t_R _23298_ (.A(_14424_),
    .B(_05598_),
    .C(_05573_),
    .Y(_05616_));
 TAPCELL_ASAP7_75t_R TAP_1048 ();
 AND4x1_ASAP7_75t_R _23300_ (.A(_14180_),
    .B(_14239_),
    .C(net310),
    .D(_05616_),
    .Y(_05618_));
 OR2x2_ASAP7_75t_R _23301_ (.A(_05615_),
    .B(_05618_),
    .Y(_05619_));
 OR3x1_ASAP7_75t_R _23302_ (.A(_14180_),
    .B(_14238_),
    .C(_05563_),
    .Y(_05620_));
 NAND2x1_ASAP7_75t_R _23303_ (.A(_14359_),
    .B(_05568_),
    .Y(_05621_));
 OAI21x1_ASAP7_75t_R _23304_ (.A1(_13495_),
    .A2(_13888_),
    .B(_14356_),
    .Y(_05622_));
 OR3x4_ASAP7_75t_R _23305_ (.A(_05622_),
    .B(_14709_),
    .C(_05600_),
    .Y(_05623_));
 AOI211x1_ASAP7_75t_R _23306_ (.A1(net302),
    .A2(_05620_),
    .B(_05621_),
    .C(_05623_),
    .Y(_05624_));
 AND2x2_ASAP7_75t_R _23307_ (.A(_14238_),
    .B(_05608_),
    .Y(_05625_));
 OR3x1_ASAP7_75t_R _23308_ (.A(_00244_),
    .B(_13474_),
    .C(_13520_),
    .Y(_05626_));
 OA211x2_ASAP7_75t_R _23309_ (.A1(_01743_),
    .A2(_05622_),
    .B(_05570_),
    .C(_05626_),
    .Y(_05627_));
 TAPCELL_ASAP7_75t_R TAP_1047 ();
 NOR2x2_ASAP7_75t_R _23311_ (.A(_14452_),
    .B(_14478_),
    .Y(_05629_));
 AO33x2_ASAP7_75t_R _23312_ (.A1(_14362_),
    .A2(_01742_),
    .A3(_14424_),
    .B1(_14420_),
    .B2(_05629_),
    .B3(_13474_),
    .Y(_05630_));
 TAPCELL_ASAP7_75t_R TAP_1046 ();
 AND3x2_ASAP7_75t_R _23314_ (.A(_05601_),
    .B(_05627_),
    .C(_05630_),
    .Y(_05632_));
 AND4x1_ASAP7_75t_R _23315_ (.A(_14296_),
    .B(_05568_),
    .C(_05583_),
    .D(_05601_),
    .Y(_05633_));
 AND2x4_ASAP7_75t_R _23316_ (.A(_14180_),
    .B(_14238_),
    .Y(_05634_));
 AO32x1_ASAP7_75t_R _23317_ (.A1(_14179_),
    .A2(_05625_),
    .A3(_05632_),
    .B1(_05633_),
    .B2(_05634_),
    .Y(_05635_));
 AO211x2_ASAP7_75t_R _23318_ (.A1(_05614_),
    .A2(_05619_),
    .B(_05624_),
    .C(_05635_),
    .Y(_05636_));
 OR4x1_ASAP7_75t_R _23319_ (.A(_05576_),
    .B(_05591_),
    .C(_05611_),
    .D(_05636_),
    .Y(_05637_));
 TAPCELL_ASAP7_75t_R TAP_1045 ();
 OA21x2_ASAP7_75t_R _23321_ (.A1(_05608_),
    .A2(_05612_),
    .B(_14179_),
    .Y(_05638_));
 XNOR2x1_ASAP7_75t_R _23322_ (.B(_14179_),
    .Y(_05639_),
    .A(net305));
 AND2x2_ASAP7_75t_R _23323_ (.A(_13525_),
    .B(_05639_),
    .Y(_05640_));
 AND2x2_ASAP7_75t_R _23324_ (.A(net302),
    .B(_05604_),
    .Y(_05641_));
 OA211x2_ASAP7_75t_R _23325_ (.A1(_05638_),
    .A2(_05640_),
    .B(_05641_),
    .C(_05564_),
    .Y(_05642_));
 NAND2x2_ASAP7_75t_R _23326_ (.A(_13528_),
    .B(_14424_),
    .Y(_05643_));
 AND4x2_ASAP7_75t_R _23327_ (.A(_14297_),
    .B(_05643_),
    .C(net310),
    .D(_05596_),
    .Y(_05644_));
 XNOR2x2_ASAP7_75t_R _23328_ (.A(_13525_),
    .B(net305),
    .Y(_05645_));
 AND3x1_ASAP7_75t_R _23329_ (.A(_14180_),
    .B(_14239_),
    .C(_05616_),
    .Y(_05646_));
 AND2x4_ASAP7_75t_R _23330_ (.A(_14179_),
    .B(_05564_),
    .Y(_05647_));
 AND4x1_ASAP7_75t_R _23331_ (.A(_18380_),
    .B(_05586_),
    .C(_05608_),
    .D(_05647_),
    .Y(_05648_));
 AO21x1_ASAP7_75t_R _23332_ (.A1(_05645_),
    .A2(_05646_),
    .B(_05648_),
    .Y(_05649_));
 AND2x2_ASAP7_75t_R _23333_ (.A(_05644_),
    .B(_05649_),
    .Y(_05650_));
 NAND2x1_ASAP7_75t_R _23334_ (.A(_13525_),
    .B(_13894_),
    .Y(_05651_));
 OR3x1_ASAP7_75t_R _23335_ (.A(_13525_),
    .B(_13894_),
    .C(_14179_),
    .Y(_05652_));
 OA21x2_ASAP7_75t_R _23336_ (.A1(_14180_),
    .A2(_05651_),
    .B(_05652_),
    .Y(_05653_));
 AND2x2_ASAP7_75t_R _23337_ (.A(_14424_),
    .B(_05572_),
    .Y(_05654_));
 AND4x1_ASAP7_75t_R _23338_ (.A(_13474_),
    .B(_14539_),
    .C(_14597_),
    .D(_14651_),
    .Y(_05655_));
 OA21x2_ASAP7_75t_R _23339_ (.A1(_05654_),
    .A2(_05655_),
    .B(_18380_),
    .Y(_05656_));
 AND3x2_ASAP7_75t_R _23340_ (.A(_05568_),
    .B(_05627_),
    .C(_05656_),
    .Y(_05657_));
 INVx3_ASAP7_75t_R _23341_ (.A(_00184_),
    .Y(_05658_));
 CKINVDCx8_ASAP7_75t_R _23342_ (.A(_00385_),
    .Y(_05659_));
 AO33x2_ASAP7_75t_R _23343_ (.A1(_05658_),
    .A2(_13520_),
    .A3(_14177_),
    .B1(_13891_),
    .B2(_13505_),
    .B3(_05659_),
    .Y(_05660_));
 AOI21x1_ASAP7_75t_R _23344_ (.A1(net2277),
    .A2(_05606_),
    .B(_13520_),
    .Y(_05661_));
 OR4x2_ASAP7_75t_R _23345_ (.A(_13474_),
    .B(_05660_),
    .C(_13892_),
    .D(_05661_),
    .Y(_05662_));
 AND3x4_ASAP7_75t_R _23346_ (.A(_13523_),
    .B(_14180_),
    .C(_05564_),
    .Y(_05663_));
 NAND2x1_ASAP7_75t_R _23347_ (.A(_05662_),
    .B(_05663_),
    .Y(_05664_));
 AO33x2_ASAP7_75t_R _23348_ (.A1(_05593_),
    .A2(_05641_),
    .A3(_05653_),
    .B1(_05657_),
    .B2(_05664_),
    .B3(_05620_),
    .Y(_05665_));
 AND2x2_ASAP7_75t_R _23349_ (.A(_05616_),
    .B(_05644_),
    .Y(_05666_));
 AND2x6_ASAP7_75t_R _23350_ (.A(_13525_),
    .B(_13894_),
    .Y(_05667_));
 TAPCELL_ASAP7_75t_R TAP_1044 ();
 AND3x1_ASAP7_75t_R _23352_ (.A(_14179_),
    .B(_14239_),
    .C(net310),
    .Y(_05669_));
 OA211x2_ASAP7_75t_R _23353_ (.A1(_05604_),
    .A2(_05666_),
    .B(_05667_),
    .C(_05669_),
    .Y(_05670_));
 OR2x2_ASAP7_75t_R _23354_ (.A(_05665_),
    .B(_05670_),
    .Y(_05671_));
 TAPCELL_ASAP7_75t_R TAP_1043 ();
 AND3x1_ASAP7_75t_R _23356_ (.A(_14179_),
    .B(_05566_),
    .C(_05604_),
    .Y(_05673_));
 AND4x1_ASAP7_75t_R _23357_ (.A(_13523_),
    .B(_05593_),
    .C(_05584_),
    .D(_05602_),
    .Y(_05674_));
 AO21x1_ASAP7_75t_R _23358_ (.A1(_13525_),
    .A2(_05673_),
    .B(_05674_),
    .Y(_05675_));
 AND2x2_ASAP7_75t_R _23359_ (.A(_05596_),
    .B(_05616_),
    .Y(_05676_));
 AND2x2_ASAP7_75t_R _23360_ (.A(_14423_),
    .B(_13521_),
    .Y(_05677_));
 AO32x2_ASAP7_75t_R _23361_ (.A1(_13474_),
    .A2(_14420_),
    .A3(_14479_),
    .B1(_05677_),
    .B2(_14363_),
    .Y(_05678_));
 AND2x2_ASAP7_75t_R _23362_ (.A(_05588_),
    .B(_05678_),
    .Y(_05679_));
 AO32x1_ASAP7_75t_R _23363_ (.A1(_05669_),
    .A2(_05667_),
    .A3(_05676_),
    .B1(_05679_),
    .B2(_05663_),
    .Y(_05680_));
 AND2x2_ASAP7_75t_R _23364_ (.A(net302),
    .B(_14359_),
    .Y(_05681_));
 AND3x1_ASAP7_75t_R _23365_ (.A(_14180_),
    .B(_14239_),
    .C(net310),
    .Y(_05682_));
 AO32x1_ASAP7_75t_R _23366_ (.A1(net310),
    .A2(_05647_),
    .A3(_05667_),
    .B1(_05682_),
    .B2(_05608_),
    .Y(_05683_));
 AND4x1_ASAP7_75t_R _23367_ (.A(_14297_),
    .B(_05643_),
    .C(net310),
    .D(_05676_),
    .Y(_05684_));
 TAPCELL_ASAP7_75t_R TAP_1042 ();
 AO21x1_ASAP7_75t_R _23369_ (.A1(_14238_),
    .A2(_05608_),
    .B(_05563_),
    .Y(_05686_));
 AO21x1_ASAP7_75t_R _23370_ (.A1(_05634_),
    .A2(_05667_),
    .B(_05686_),
    .Y(_05687_));
 AO32x1_ASAP7_75t_R _23371_ (.A1(net302),
    .A2(_05604_),
    .A3(_05683_),
    .B1(_05684_),
    .B2(_05687_),
    .Y(_05688_));
 AO221x1_ASAP7_75t_R _23372_ (.A1(_13894_),
    .A2(_05675_),
    .B1(_05680_),
    .B2(_05681_),
    .C(_05688_),
    .Y(_05689_));
 OR5x1_ASAP7_75t_R _23373_ (.A(_05637_),
    .B(_05642_),
    .C(_05650_),
    .D(_05671_),
    .E(_05689_),
    .Y(_05690_));
 AO21x1_ASAP7_75t_R _23374_ (.A1(_05627_),
    .A2(_05630_),
    .B(_05614_),
    .Y(_05691_));
 AO32x1_ASAP7_75t_R _23375_ (.A1(_05568_),
    .A2(_05593_),
    .A3(_05584_),
    .B1(_05691_),
    .B2(_05634_),
    .Y(_05692_));
 AO31x2_ASAP7_75t_R _23376_ (.A1(_14180_),
    .A2(_14238_),
    .A3(_05608_),
    .B(_05563_),
    .Y(_05693_));
 TAPCELL_ASAP7_75t_R TAP_1041 ();
 AO21x1_ASAP7_75t_R _23378_ (.A1(_14238_),
    .A2(_05608_),
    .B(_14358_),
    .Y(_05694_));
 OA211x2_ASAP7_75t_R _23379_ (.A1(_14359_),
    .A2(_05693_),
    .B(_05694_),
    .C(_14296_),
    .Y(_05695_));
 OA21x2_ASAP7_75t_R _23380_ (.A1(_05563_),
    .A2(_05695_),
    .B(_05602_),
    .Y(_05696_));
 AO21x1_ASAP7_75t_R _23381_ (.A1(_05601_),
    .A2(_05692_),
    .B(_05696_),
    .Y(_05697_));
 AND4x2_ASAP7_75t_R _23382_ (.A(net302),
    .B(_14359_),
    .C(_05596_),
    .D(_05616_),
    .Y(_05698_));
 AND2x2_ASAP7_75t_R _23383_ (.A(_13525_),
    .B(net305),
    .Y(_05699_));
 AND3x1_ASAP7_75t_R _23384_ (.A(_05566_),
    .B(_05583_),
    .C(_05602_),
    .Y(_05700_));
 AO32x1_ASAP7_75t_R _23385_ (.A1(_05564_),
    .A2(_05667_),
    .A3(_05698_),
    .B1(_05699_),
    .B2(_05700_),
    .Y(_05701_));
 AND2x2_ASAP7_75t_R _23386_ (.A(net305),
    .B(_14180_),
    .Y(_05702_));
 XNOR2x1_ASAP7_75t_R _23387_ (.B(_05667_),
    .Y(_05703_),
    .A(_14180_));
 OA211x2_ASAP7_75t_R _23388_ (.A1(_05702_),
    .A2(_05703_),
    .B(_05698_),
    .C(_05593_),
    .Y(_05704_));
 AND3x1_ASAP7_75t_R _23389_ (.A(net305),
    .B(_05564_),
    .C(_05698_),
    .Y(_05705_));
 AO21x1_ASAP7_75t_R _23390_ (.A1(_13894_),
    .A2(_05700_),
    .B(_05705_),
    .Y(_05706_));
 AND2x2_ASAP7_75t_R _23391_ (.A(_13523_),
    .B(net305),
    .Y(_05707_));
 AND2x2_ASAP7_75t_R _23392_ (.A(_05564_),
    .B(_05698_),
    .Y(_05708_));
 AO221x1_ASAP7_75t_R _23393_ (.A1(_05707_),
    .A2(_05708_),
    .B1(_05700_),
    .B2(_05608_),
    .C(_14180_),
    .Y(_05709_));
 OA21x2_ASAP7_75t_R _23394_ (.A1(_14179_),
    .A2(_05706_),
    .B(_05709_),
    .Y(_05710_));
 AND2x2_ASAP7_75t_R _23395_ (.A(_14179_),
    .B(_14238_),
    .Y(_05711_));
 AND2x2_ASAP7_75t_R _23396_ (.A(_05612_),
    .B(_05711_),
    .Y(_05712_));
 OA211x2_ASAP7_75t_R _23397_ (.A1(_13525_),
    .A2(_05608_),
    .B(_14239_),
    .C(_14180_),
    .Y(_05713_));
 OA211x2_ASAP7_75t_R _23398_ (.A1(_05712_),
    .A2(_05713_),
    .B(_05584_),
    .C(_05602_),
    .Y(_05714_));
 OA211x2_ASAP7_75t_R _23399_ (.A1(_05684_),
    .A2(_05698_),
    .B(_05647_),
    .C(_05645_),
    .Y(_05715_));
 OR5x1_ASAP7_75t_R _23400_ (.A(_05701_),
    .B(_05704_),
    .C(_05710_),
    .D(_05714_),
    .E(_05715_),
    .Y(_05716_));
 AND2x2_ASAP7_75t_R _23401_ (.A(_05667_),
    .B(_05682_),
    .Y(_05717_));
 AO21x1_ASAP7_75t_R _23402_ (.A1(_05669_),
    .A2(_05651_),
    .B(_05717_),
    .Y(_05718_));
 TAPCELL_ASAP7_75t_R TAP_1040 ();
 AND3x1_ASAP7_75t_R _23404_ (.A(net310),
    .B(_05634_),
    .C(_05645_),
    .Y(_05720_));
 OR3x1_ASAP7_75t_R _23405_ (.A(_05683_),
    .B(_05718_),
    .C(_05720_),
    .Y(_05721_));
 AND2x2_ASAP7_75t_R _23406_ (.A(_05666_),
    .B(_05721_),
    .Y(_05722_));
 OR4x2_ASAP7_75t_R _23407_ (.A(_05690_),
    .B(_05697_),
    .C(_05716_),
    .D(_05722_),
    .Y(_05723_));
 INVx3_ASAP7_75t_R _23408_ (.A(_01311_),
    .Y(_05724_));
 OR5x2_ASAP7_75t_R _23409_ (.A(_01317_),
    .B(_00172_),
    .C(_13470_),
    .D(_13463_),
    .E(_13803_),
    .Y(_05725_));
 TAPCELL_ASAP7_75t_R TAP_1039 ();
 OR3x4_ASAP7_75t_R _23411_ (.A(_14799_),
    .B(_14806_),
    .C(_05725_),
    .Y(_05727_));
 OR3x4_ASAP7_75t_R _23412_ (.A(_14808_),
    .B(_14799_),
    .C(_05725_),
    .Y(_05728_));
 OR3x1_ASAP7_75t_R _23413_ (.A(_14383_),
    .B(_14802_),
    .C(_14803_),
    .Y(_05729_));
 OR4x1_ASAP7_75t_R _23414_ (.A(_01997_),
    .B(_14808_),
    .C(_05729_),
    .D(_05725_),
    .Y(_05730_));
 TAPCELL_ASAP7_75t_R TAP_1038 ();
 NOR2x1_ASAP7_75t_R _23416_ (.A(_17810_),
    .B(_02140_),
    .Y(_05732_));
 AO21x1_ASAP7_75t_R _23417_ (.A1(_05728_),
    .A2(_05730_),
    .B(_05732_),
    .Y(_05733_));
 INVx1_ASAP7_75t_R _23418_ (.A(_02285_),
    .Y(_05734_));
 OAI21x1_ASAP7_75t_R _23419_ (.A1(_05734_),
    .A2(_02284_),
    .B(_02283_),
    .Y(_05735_));
 OA21x2_ASAP7_75t_R _23420_ (.A1(_01313_),
    .A2(_02284_),
    .B(_05735_),
    .Y(_05736_));
 AND2x2_ASAP7_75t_R _23421_ (.A(_14797_),
    .B(_05570_),
    .Y(_05737_));
 AND4x1_ASAP7_75t_R _23422_ (.A(_02288_),
    .B(_14653_),
    .C(_18380_),
    .D(_05737_),
    .Y(_05738_));
 NOR2x2_ASAP7_75t_R _23423_ (.A(_05736_),
    .B(_05738_),
    .Y(_05739_));
 OR3x1_ASAP7_75t_R _23424_ (.A(_01317_),
    .B(_13804_),
    .C(_05739_),
    .Y(_05740_));
 OA211x2_ASAP7_75t_R _23425_ (.A1(_05724_),
    .A2(_05727_),
    .B(_05733_),
    .C(_05740_),
    .Y(_05741_));
 OA211x2_ASAP7_75t_R _23426_ (.A1(_01317_),
    .A2(_14842_),
    .B(_05723_),
    .C(_05741_),
    .Y(_05742_));
 NOR2x1_ASAP7_75t_R _23427_ (.A(_05557_),
    .B(_05742_),
    .Y(\id_stage_i.controller_i.illegal_insn_d ));
 TAPCELL_ASAP7_75t_R TAP_1037 ();
 INVx3_ASAP7_75t_R _23429_ (.A(_01721_),
    .Y(_05744_));
 AND4x2_ASAP7_75t_R _23430_ (.A(_13802_),
    .B(_05546_),
    .C(_14813_),
    .D(_14814_),
    .Y(_05745_));
 NOR2x2_ASAP7_75t_R _23431_ (.A(_05744_),
    .B(_05745_),
    .Y(_05746_));
 AO21x1_ASAP7_75t_R _23432_ (.A1(_14842_),
    .A2(_05746_),
    .B(_01317_),
    .Y(_05747_));
 AND3x2_ASAP7_75t_R _23433_ (.A(_05723_),
    .B(_05741_),
    .C(_05747_),
    .Y(_05748_));
 NOR2x1_ASAP7_75t_R _23434_ (.A(_05557_),
    .B(_05748_),
    .Y(\id_stage_i.controller_i.exc_req_d ));
 TAPCELL_ASAP7_75t_R TAP_1036 ();
 INVx1_ASAP7_75t_R _23436_ (.A(_01731_),
    .Y(_05750_));
 TAPCELL_ASAP7_75t_R TAP_1035 ();
 AND2x6_ASAP7_75t_R _23438_ (.A(_14797_),
    .B(_14842_),
    .Y(_05752_));
 AND3x2_ASAP7_75t_R _23439_ (.A(_01713_),
    .B(_14828_),
    .C(_05752_),
    .Y(_05753_));
 AND2x2_ASAP7_75t_R _23440_ (.A(_01608_),
    .B(_05753_),
    .Y(_05754_));
 INVx1_ASAP7_75t_R _23441_ (.A(_05754_),
    .Y(_05755_));
 TAPCELL_ASAP7_75t_R TAP_1034 ();
 NAND2x1_ASAP7_75t_R _23443_ (.A(_00277_),
    .B(net3030),
    .Y(_05757_));
 AO21x2_ASAP7_75t_R _23444_ (.A1(_01609_),
    .A2(_05755_),
    .B(_05757_),
    .Y(_05758_));
 OA211x2_ASAP7_75t_R _23445_ (.A1(_13446_),
    .A2(_05754_),
    .B(_00277_),
    .C(net3030),
    .Y(_05759_));
 AND3x4_ASAP7_75t_R _23446_ (.A(_13574_),
    .B(_14828_),
    .C(_05759_),
    .Y(_05760_));
 AO21x1_ASAP7_75t_R _23447_ (.A1(_05750_),
    .A2(_05758_),
    .B(_05760_),
    .Y(_00007_));
 TAPCELL_ASAP7_75t_R TAP_1033 ();
 INVx2_ASAP7_75t_R _23449_ (.A(_01730_),
    .Y(_05762_));
 AND2x2_ASAP7_75t_R _23450_ (.A(_00282_),
    .B(_14828_),
    .Y(_05763_));
 AND3x4_ASAP7_75t_R _23451_ (.A(_00281_),
    .B(_05759_),
    .C(_05763_),
    .Y(_05764_));
 AO21x1_ASAP7_75t_R _23452_ (.A1(_05762_),
    .A2(_05758_),
    .B(_05764_),
    .Y(_00006_));
 INVx2_ASAP7_75t_R _23453_ (.A(_01357_),
    .Y(_05765_));
 AND3x4_ASAP7_75t_R _23454_ (.A(_13570_),
    .B(_13534_),
    .C(_13537_),
    .Y(_05766_));
 TAPCELL_ASAP7_75t_R TAP_1032 ();
 TAPCELL_ASAP7_75t_R TAP_1031 ();
 NAND2x2_ASAP7_75t_R _23457_ (.A(_05752_),
    .B(_05766_),
    .Y(_05769_));
 TAPCELL_ASAP7_75t_R TAP_1030 ();
 NAND2x2_ASAP7_75t_R _23459_ (.A(_01322_),
    .B(_17825_),
    .Y(_05771_));
 TAPCELL_ASAP7_75t_R TAP_1029 ();
 INVx3_ASAP7_75t_R _23461_ (.A(_01318_),
    .Y(_05773_));
 OR2x4_ASAP7_75t_R _23462_ (.A(_01319_),
    .B(_05773_),
    .Y(_05774_));
 OR3x1_ASAP7_75t_R _23463_ (.A(_05769_),
    .B(_05771_),
    .C(_05774_),
    .Y(_05775_));
 INVx2_ASAP7_75t_R _23464_ (.A(_01873_),
    .Y(_05776_));
 AND3x4_ASAP7_75t_R _23465_ (.A(_14797_),
    .B(_14842_),
    .C(_05766_),
    .Y(_05777_));
 TAPCELL_ASAP7_75t_R TAP_1028 ();
 AND2x6_ASAP7_75t_R _23467_ (.A(_05776_),
    .B(_05777_),
    .Y(_05779_));
 TAPCELL_ASAP7_75t_R TAP_1027 ();
 AO21x1_ASAP7_75t_R _23469_ (.A1(_05765_),
    .A2(_05775_),
    .B(_05779_),
    .Y(_00005_));
 INVx4_ASAP7_75t_R _23470_ (.A(_00284_),
    .Y(_05781_));
 INVx2_ASAP7_75t_R _23471_ (.A(_01872_),
    .Y(_05782_));
 INVx5_ASAP7_75t_R _23472_ (.A(_00676_),
    .Y(net178));
 TAPCELL_ASAP7_75t_R TAP_1026 ();
 TAPCELL_ASAP7_75t_R TAP_1025 ();
 TAPCELL_ASAP7_75t_R TAP_1024 ();
 OR4x1_ASAP7_75t_R _23476_ (.A(net289),
    .B(net180),
    .C(net262),
    .D(_18555_),
    .Y(_05786_));
 OR5x1_ASAP7_75t_R _23477_ (.A(net293),
    .B(net154),
    .C(net259),
    .D(net156),
    .E(_05786_),
    .Y(_05787_));
 OR4x1_ASAP7_75t_R _23478_ (.A(net2179),
    .B(net2171),
    .C(net2152),
    .D(net2138),
    .Y(_05788_));
 OR5x1_ASAP7_75t_R _23479_ (.A(net178),
    .B(net261),
    .C(net258),
    .D(_05787_),
    .E(_05788_),
    .Y(_05789_));
 INVx1_ASAP7_75t_R _23480_ (.A(_05789_),
    .Y(_05790_));
 XOR2x2_ASAP7_75t_R _23481_ (.A(_02264_),
    .B(_02223_),
    .Y(_05791_));
 XOR2x2_ASAP7_75t_R _23482_ (.A(_02262_),
    .B(_02222_),
    .Y(_05792_));
 XOR2x2_ASAP7_75t_R _23483_ (.A(_02224_),
    .B(_02266_),
    .Y(_05793_));
 AND5x1_ASAP7_75t_R _23484_ (.A(_05404_),
    .B(_05790_),
    .C(_05791_),
    .D(_05792_),
    .E(_05793_),
    .Y(_05794_));
 XNOR2x2_ASAP7_75t_R _23485_ (.A(_00818_),
    .B(_02275_),
    .Y(_05795_));
 XOR2x2_ASAP7_75t_R _23486_ (.A(_02272_),
    .B(_02226_),
    .Y(_05796_));
 XOR2x2_ASAP7_75t_R _23487_ (.A(_02270_),
    .B(_02225_),
    .Y(_05797_));
 XNOR2x2_ASAP7_75t_R _23488_ (.A(_00679_),
    .B(_02268_),
    .Y(_05798_));
 AND4x1_ASAP7_75t_R _23489_ (.A(_05795_),
    .B(_05796_),
    .C(_05797_),
    .D(_05798_),
    .Y(_05799_));
 AND5x1_ASAP7_75t_R _23490_ (.A(_15778_),
    .B(_04747_),
    .C(_04968_),
    .D(_05185_),
    .E(_05799_),
    .Y(_05800_));
 AND5x2_ASAP7_75t_R _23491_ (.A(_16263_),
    .B(_16509_),
    .C(_04517_),
    .D(_05794_),
    .E(_05800_),
    .Y(_05801_));
 NAND2x2_ASAP7_75t_R _23492_ (.A(_05542_),
    .B(_05801_),
    .Y(_05802_));
 AND3x1_ASAP7_75t_R _23493_ (.A(_05782_),
    .B(_05777_),
    .C(_05802_),
    .Y(_05803_));
 AO21x1_ASAP7_75t_R _23494_ (.A1(_05781_),
    .A2(_05769_),
    .B(_05803_),
    .Y(_00004_));
 TAPCELL_ASAP7_75t_R TAP_1023 ();
 OA211x2_ASAP7_75t_R _23496_ (.A1(_01872_),
    .A2(_05802_),
    .B(_05777_),
    .C(_00285_),
    .Y(_05805_));
 AOI21x1_ASAP7_75t_R _23497_ (.A1(_01728_),
    .A2(_05769_),
    .B(_05805_),
    .Y(_00003_));
 TAPCELL_ASAP7_75t_R TAP_1022 ();
 TAPCELL_ASAP7_75t_R TAP_1021 ();
 NAND2x2_ASAP7_75t_R _23500_ (.A(_05765_),
    .B(_05777_),
    .Y(_05808_));
 TAPCELL_ASAP7_75t_R TAP_1020 ();
 OR3x1_ASAP7_75t_R _23502_ (.A(_05771_),
    .B(_05774_),
    .C(_05808_),
    .Y(_05810_));
 OAI21x1_ASAP7_75t_R _23503_ (.A1(_01727_),
    .A2(_05777_),
    .B(_05810_),
    .Y(_00002_));
 INVx5_ASAP7_75t_R _23504_ (.A(_05792_),
    .Y(net171));
 INVx4_ASAP7_75t_R _23505_ (.A(_05791_),
    .Y(net175));
 INVx4_ASAP7_75t_R _23506_ (.A(_05793_),
    .Y(net177));
 INVx3_ASAP7_75t_R _23507_ (.A(_05798_),
    .Y(net179));
 CKINVDCx5p33_ASAP7_75t_R _23508_ (.A(_05797_),
    .Y(net151));
 INVx6_ASAP7_75t_R _23509_ (.A(_05796_),
    .Y(net153));
 INVx3_ASAP7_75t_R _23510_ (.A(_05795_),
    .Y(net157));
 AND3x2_ASAP7_75t_R _23511_ (.A(_13456_),
    .B(_14828_),
    .C(_14842_),
    .Y(net218));
 TAPCELL_ASAP7_75t_R TAP_1019 ();
 INVx4_ASAP7_75t_R _23513_ (.A(_17818_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ));
 INVx1_ASAP7_75t_R _23514_ (.A(_02291_),
    .Y(_17821_));
 INVx2_ASAP7_75t_R _23515_ (.A(\ex_block_i.alu_adder_result_ex_o[0] ),
    .Y(_16721_));
 INVx4_ASAP7_75t_R _23516_ (.A(net296),
    .Y(_16717_));
 TAPCELL_ASAP7_75t_R TAP_1018 ();
 AND2x6_ASAP7_75t_R _23518_ (.A(_01314_),
    .B(_01875_),
    .Y(_05813_));
 TAPCELL_ASAP7_75t_R TAP_1017 ();
 NOR3x2_ASAP7_75t_R _23520_ (.B(_05546_),
    .C(_05547_),
    .Y(_05815_),
    .A(_05545_));
 OR2x2_ASAP7_75t_R _23521_ (.A(_01874_),
    .B(_05815_),
    .Y(_05816_));
 AND2x6_ASAP7_75t_R _23522_ (.A(_05813_),
    .B(_05816_),
    .Y(_05817_));
 TAPCELL_ASAP7_75t_R TAP_1016 ();
 OAI22x1_ASAP7_75t_R _23524_ (.A1(_00324_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00816_),
    .Y(_17826_));
 NAND2x2_ASAP7_75t_R _23525_ (.A(_01314_),
    .B(_01875_),
    .Y(_05819_));
 AND3x1_ASAP7_75t_R _23526_ (.A(_15933_),
    .B(_15971_),
    .C(_05819_),
    .Y(_05820_));
 AO21x2_ASAP7_75t_R _23527_ (.A1(_13886_),
    .A2(_05813_),
    .B(_05820_),
    .Y(_05821_));
 TAPCELL_ASAP7_75t_R TAP_1015 ();
 AND2x4_ASAP7_75t_R _23529_ (.A(_15994_),
    .B(_16017_),
    .Y(_05823_));
 NAND2x2_ASAP7_75t_R _23530_ (.A(_01314_),
    .B(_01874_),
    .Y(_05824_));
 TAPCELL_ASAP7_75t_R TAP_1014 ();
 AND3x1_ASAP7_75t_R _23532_ (.A(_01314_),
    .B(_01874_),
    .C(_13981_),
    .Y(_05826_));
 AO21x2_ASAP7_75t_R _23533_ (.A1(_05823_),
    .A2(_05824_),
    .B(_05826_),
    .Y(_05827_));
 TAPCELL_ASAP7_75t_R TAP_1013 ();
 AND2x2_ASAP7_75t_R _23535_ (.A(_05821_),
    .B(_05827_),
    .Y(_17827_));
 OAI22x1_ASAP7_75t_R _23536_ (.A1(_00291_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00849_),
    .Y(_17833_));
 TAPCELL_ASAP7_75t_R TAP_1012 ();
 TAPCELL_ASAP7_75t_R TAP_1011 ();
 OAI22x1_ASAP7_75t_R _23539_ (.A1(_00663_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00881_),
    .Y(_17840_));
 TAPCELL_ASAP7_75t_R TAP_1010 ();
 AND2x2_ASAP7_75t_R _23541_ (.A(_14169_),
    .B(_05813_),
    .Y(_05832_));
 AO21x2_ASAP7_75t_R _23542_ (.A1(_16213_),
    .A2(_05819_),
    .B(_05832_),
    .Y(_05833_));
 TAPCELL_ASAP7_75t_R TAP_1009 ();
 TAPCELL_ASAP7_75t_R TAP_1008 ();
 NAND2x1_ASAP7_75t_R _23545_ (.A(_05827_),
    .B(_05833_),
    .Y(_16764_));
 OAI22x1_ASAP7_75t_R _23546_ (.A1(_00665_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00914_),
    .Y(_17844_));
 AND2x2_ASAP7_75t_R _23547_ (.A(_14233_),
    .B(_05813_),
    .Y(_05836_));
 AO21x2_ASAP7_75t_R _23548_ (.A1(_16324_),
    .A2(_05819_),
    .B(_05836_),
    .Y(_05837_));
 TAPCELL_ASAP7_75t_R TAP_1007 ();
 AND2x2_ASAP7_75t_R _23550_ (.A(_05827_),
    .B(net2370),
    .Y(_17845_));
 AO21x1_ASAP7_75t_R _23551_ (.A1(_01314_),
    .A2(_01874_),
    .B(_16138_),
    .Y(_05839_));
 OA21x2_ASAP7_75t_R _23552_ (.A1(_13767_),
    .A2(_05824_),
    .B(_05839_),
    .Y(_05840_));
 TAPCELL_ASAP7_75t_R TAP_1006 ();
 NAND2x1_ASAP7_75t_R _23554_ (.A(_05833_),
    .B(_05840_),
    .Y(_16767_));
 TAPCELL_ASAP7_75t_R TAP_1005 ();
 OAI22x1_ASAP7_75t_R _23556_ (.A1(_00668_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00946_),
    .Y(_17859_));
 INVx1_ASAP7_75t_R _23557_ (.A(_16261_),
    .Y(_05843_));
 AND3x1_ASAP7_75t_R _23558_ (.A(_01314_),
    .B(_01874_),
    .C(_14921_),
    .Y(_05844_));
 AO21x2_ASAP7_75t_R _23559_ (.A1(_05843_),
    .A2(_05824_),
    .B(_05844_),
    .Y(_05845_));
 TAPCELL_ASAP7_75t_R TAP_1004 ();
 NAND2x1_ASAP7_75t_R _23561_ (.A(_05833_),
    .B(_05845_),
    .Y(_16774_));
 TAPCELL_ASAP7_75t_R TAP_1003 ();
 OAI22x1_ASAP7_75t_R _23563_ (.A1(_00670_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_00979_),
    .Y(_17869_));
 NOR2x1_ASAP7_75t_R _23564_ (.A(_16568_),
    .B(_05813_),
    .Y(_05848_));
 AO21x2_ASAP7_75t_R _23565_ (.A1(_14355_),
    .A2(_05813_),
    .B(_05848_),
    .Y(_05849_));
 TAPCELL_ASAP7_75t_R TAP_1002 ();
 AND2x2_ASAP7_75t_R _23567_ (.A(_05827_),
    .B(net2253),
    .Y(_16784_));
 AND2x2_ASAP7_75t_R _23568_ (.A(_14290_),
    .B(_05813_),
    .Y(_05851_));
 AO21x2_ASAP7_75t_R _23569_ (.A1(_16456_),
    .A2(_05819_),
    .B(_05851_),
    .Y(_05852_));
 TAPCELL_ASAP7_75t_R TAP_1001 ();
 AND2x2_ASAP7_75t_R _23571_ (.A(_05840_),
    .B(_05852_),
    .Y(_16785_));
 AND2x2_ASAP7_75t_R _23572_ (.A(net2370),
    .B(_05845_),
    .Y(_16786_));
 AO21x1_ASAP7_75t_R _23573_ (.A1(_01314_),
    .A2(_01874_),
    .B(_16378_),
    .Y(_05854_));
 OA21x2_ASAP7_75t_R _23574_ (.A1(_14980_),
    .A2(_05824_),
    .B(_05854_),
    .Y(_05855_));
 TAPCELL_ASAP7_75t_R TAP_1000 ();
 NAND2x1_ASAP7_75t_R _23576_ (.A(_05833_),
    .B(_05855_),
    .Y(_16788_));
 TAPCELL_ASAP7_75t_R TAP_999 ();
 OAI22x1_ASAP7_75t_R _23578_ (.A1(_00672_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01011_),
    .Y(_17875_));
 AND3x1_ASAP7_75t_R _23579_ (.A(_16647_),
    .B(_16678_),
    .C(_05819_),
    .Y(_05858_));
 AO21x2_ASAP7_75t_R _23580_ (.A1(_14420_),
    .A2(_05813_),
    .B(_05858_),
    .Y(_05859_));
 TAPCELL_ASAP7_75t_R TAP_998 ();
 AND2x2_ASAP7_75t_R _23582_ (.A(_05827_),
    .B(_05859_),
    .Y(_17872_));
 AND2x2_ASAP7_75t_R _23583_ (.A(_05840_),
    .B(net2253),
    .Y(_16805_));
 AND2x2_ASAP7_75t_R _23584_ (.A(_05845_),
    .B(_05852_),
    .Y(_16806_));
 AND2x2_ASAP7_75t_R _23585_ (.A(net2370),
    .B(_05855_),
    .Y(_16807_));
 OA21x2_ASAP7_75t_R _23586_ (.A1(_13626_),
    .A2(_16481_),
    .B(_16506_),
    .Y(_05861_));
 AND3x1_ASAP7_75t_R _23587_ (.A(_01314_),
    .B(_01874_),
    .C(_15050_),
    .Y(_05862_));
 AO21x2_ASAP7_75t_R _23588_ (.A1(_05861_),
    .A2(_05824_),
    .B(_05862_),
    .Y(_05863_));
 TAPCELL_ASAP7_75t_R TAP_997 ();
 NAND2x1_ASAP7_75t_R _23590_ (.A(_05833_),
    .B(_05863_),
    .Y(_16809_));
 TAPCELL_ASAP7_75t_R TAP_996 ();
 OAI22x1_ASAP7_75t_R _23592_ (.A1(_00674_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01045_),
    .Y(_17887_));
 AND2x2_ASAP7_75t_R _23593_ (.A(_14479_),
    .B(_05813_),
    .Y(_05866_));
 AO21x2_ASAP7_75t_R _23594_ (.A1(_04576_),
    .A2(_05819_),
    .B(_05866_),
    .Y(_05867_));
 TAPCELL_ASAP7_75t_R TAP_995 ();
 AND2x2_ASAP7_75t_R _23596_ (.A(_05827_),
    .B(_05867_),
    .Y(_17881_));
 AND2x2_ASAP7_75t_R _23597_ (.A(_05840_),
    .B(_05859_),
    .Y(_17882_));
 AND2x2_ASAP7_75t_R _23598_ (.A(_05845_),
    .B(_05849_),
    .Y(_16824_));
 AND2x2_ASAP7_75t_R _23599_ (.A(_05852_),
    .B(_05855_),
    .Y(_16825_));
 AND2x2_ASAP7_75t_R _23600_ (.A(_05837_),
    .B(_05863_),
    .Y(_16826_));
 AO21x1_ASAP7_75t_R _23601_ (.A1(_01314_),
    .A2(_01874_),
    .B(_16617_),
    .Y(_05869_));
 OA21x2_ASAP7_75t_R _23602_ (.A1(_15103_),
    .A2(_05824_),
    .B(_05869_),
    .Y(_05870_));
 TAPCELL_ASAP7_75t_R TAP_994 ();
 NAND2x1_ASAP7_75t_R _23604_ (.A(_05833_),
    .B(_05870_),
    .Y(_16828_));
 TAPCELL_ASAP7_75t_R TAP_993 ();
 OAI22x1_ASAP7_75t_R _23606_ (.A1(_00677_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01077_),
    .Y(_17894_));
 AND3x1_ASAP7_75t_R _23607_ (.A(_04664_),
    .B(_04696_),
    .C(_05819_),
    .Y(_05873_));
 AO21x2_ASAP7_75t_R _23608_ (.A1(_14539_),
    .A2(_05813_),
    .B(_05873_),
    .Y(_05874_));
 TAPCELL_ASAP7_75t_R TAP_992 ();
 TAPCELL_ASAP7_75t_R TAP_991 ();
 NAND2x1_ASAP7_75t_R _23611_ (.A(_05827_),
    .B(_05874_),
    .Y(_16842_));
 AND2x2_ASAP7_75t_R _23612_ (.A(net2253),
    .B(net2345),
    .Y(_16846_));
 AND2x2_ASAP7_75t_R _23613_ (.A(_05852_),
    .B(_05863_),
    .Y(_16847_));
 AND2x2_ASAP7_75t_R _23614_ (.A(_05837_),
    .B(_05870_),
    .Y(_16848_));
 AO22x2_ASAP7_75t_R _23615_ (.A1(_16692_),
    .A2(_16703_),
    .B1(_04504_),
    .B2(_04513_),
    .Y(_05877_));
 AO21x1_ASAP7_75t_R _23616_ (.A1(_01314_),
    .A2(_01874_),
    .B(_05877_),
    .Y(_05878_));
 OA21x2_ASAP7_75t_R _23617_ (.A1(_15167_),
    .A2(_05824_),
    .B(_05878_),
    .Y(_05879_));
 TAPCELL_ASAP7_75t_R TAP_990 ();
 NAND2x2_ASAP7_75t_R _23619_ (.A(_05833_),
    .B(_05879_),
    .Y(_16854_));
 TAPCELL_ASAP7_75t_R TAP_989 ();
 OAI22x1_ASAP7_75t_R _23621_ (.A1(_00680_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01110_),
    .Y(_17899_));
 NOR2x1_ASAP7_75t_R _23622_ (.A(_04808_),
    .B(_05813_),
    .Y(_05882_));
 AO21x2_ASAP7_75t_R _23623_ (.A1(_14597_),
    .A2(_05813_),
    .B(_05882_),
    .Y(_05883_));
 TAPCELL_ASAP7_75t_R TAP_988 ();
 AND2x2_ASAP7_75t_R _23625_ (.A(_05827_),
    .B(_05883_),
    .Y(_17900_));
 NAND2x1_ASAP7_75t_R _23626_ (.A(_05840_),
    .B(_05874_),
    .Y(_16872_));
 AND2x2_ASAP7_75t_R _23627_ (.A(net2253),
    .B(_05863_),
    .Y(_16877_));
 AND2x2_ASAP7_75t_R _23628_ (.A(_05852_),
    .B(_05870_),
    .Y(_16878_));
 AND2x2_ASAP7_75t_R _23629_ (.A(net2370),
    .B(net2353),
    .Y(_16879_));
 NAND2x2_ASAP7_75t_R _23630_ (.A(_15196_),
    .B(_15222_),
    .Y(_05885_));
 NOR2x1_ASAP7_75t_R _23631_ (.A(_05885_),
    .B(_05824_),
    .Y(_05886_));
 AO21x2_ASAP7_75t_R _23632_ (.A1(_04624_),
    .A2(_05824_),
    .B(_05886_),
    .Y(_05887_));
 TAPCELL_ASAP7_75t_R TAP_987 ();
 NAND2x2_ASAP7_75t_R _23634_ (.A(_05833_),
    .B(net2317),
    .Y(_16881_));
 TAPCELL_ASAP7_75t_R TAP_986 ();
 TAPCELL_ASAP7_75t_R TAP_985 ();
 TAPCELL_ASAP7_75t_R TAP_984 ();
 OAI22x1_ASAP7_75t_R _23638_ (.A1(_00682_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01142_),
    .Y(_17916_));
 NAND2x1_ASAP7_75t_R _23639_ (.A(net2337),
    .B(_05874_),
    .Y(_16896_));
 AND2x2_ASAP7_75t_R _23640_ (.A(_05849_),
    .B(_05870_),
    .Y(_16901_));
 AND2x2_ASAP7_75t_R _23641_ (.A(_05852_),
    .B(net2353),
    .Y(_16902_));
 AND2x2_ASAP7_75t_R _23642_ (.A(_05837_),
    .B(net2316),
    .Y(_16903_));
 OA21x2_ASAP7_75t_R _23643_ (.A1(net378),
    .A2(_04723_),
    .B(_04744_),
    .Y(_05892_));
 AND3x1_ASAP7_75t_R _23644_ (.A(_01314_),
    .B(_01874_),
    .C(_15279_),
    .Y(_05893_));
 AO21x2_ASAP7_75t_R _23645_ (.A1(_05892_),
    .A2(_05824_),
    .B(_05893_),
    .Y(_05894_));
 TAPCELL_ASAP7_75t_R TAP_983 ();
 TAPCELL_ASAP7_75t_R TAP_982 ();
 NAND2x1_ASAP7_75t_R _23648_ (.A(net2223),
    .B(_05894_),
    .Y(_16909_));
 TAPCELL_ASAP7_75t_R TAP_981 ();
 OAI22x1_ASAP7_75t_R _23650_ (.A1(_00684_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01176_),
    .Y(_17928_));
 AO211x2_ASAP7_75t_R _23651_ (.A1(_14666_),
    .A2(_14677_),
    .B(_14689_),
    .C(_14702_),
    .Y(_05898_));
 AND3x1_ASAP7_75t_R _23652_ (.A(_04995_),
    .B(_05027_),
    .C(_05819_),
    .Y(_05899_));
 AO21x2_ASAP7_75t_R _23653_ (.A1(_05898_),
    .A2(_05813_),
    .B(_05899_),
    .Y(_05900_));
 TAPCELL_ASAP7_75t_R TAP_980 ();
 TAPCELL_ASAP7_75t_R TAP_979 ();
 NAND2x1_ASAP7_75t_R _23656_ (.A(_05827_),
    .B(_05900_),
    .Y(_16926_));
 NAND2x1_ASAP7_75t_R _23657_ (.A(net2346),
    .B(_05874_),
    .Y(_16929_));
 AND2x2_ASAP7_75t_R _23658_ (.A(net2253),
    .B(net2353),
    .Y(_16934_));
 AND2x2_ASAP7_75t_R _23659_ (.A(_05852_),
    .B(net2316),
    .Y(_16935_));
 AND2x2_ASAP7_75t_R _23660_ (.A(net2370),
    .B(_05894_),
    .Y(_16936_));
 AO21x1_ASAP7_75t_R _23661_ (.A1(_01314_),
    .A2(_01874_),
    .B(_04854_),
    .Y(_05903_));
 OA21x2_ASAP7_75t_R _23662_ (.A1(_15331_),
    .A2(_05824_),
    .B(_05903_),
    .Y(_05904_));
 TAPCELL_ASAP7_75t_R TAP_978 ();
 TAPCELL_ASAP7_75t_R TAP_977 ();
 NAND2x1_ASAP7_75t_R _23665_ (.A(net2223),
    .B(_05904_),
    .Y(_16942_));
 OAI22x1_ASAP7_75t_R _23666_ (.A1(_00686_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01208_),
    .Y(_17942_));
 AND3x2_ASAP7_75t_R _23667_ (.A(_05104_),
    .B(_05135_),
    .C(_05819_),
    .Y(_05907_));
 AO21x2_ASAP7_75t_R _23668_ (.A1(_15487_),
    .A2(_05813_),
    .B(_05907_),
    .Y(_05908_));
 TAPCELL_ASAP7_75t_R TAP_976 ();
 TAPCELL_ASAP7_75t_R TAP_975 ();
 AND2x2_ASAP7_75t_R _23671_ (.A(_05827_),
    .B(_05908_),
    .Y(_17943_));
 NAND2x1_ASAP7_75t_R _23672_ (.A(_05840_),
    .B(_05900_),
    .Y(_16958_));
 NAND2x1_ASAP7_75t_R _23673_ (.A(net2285),
    .B(_05874_),
    .Y(_16961_));
 AND2x2_ASAP7_75t_R _23674_ (.A(_05849_),
    .B(net2316),
    .Y(_16966_));
 AND2x2_ASAP7_75t_R _23675_ (.A(_05852_),
    .B(_05894_),
    .Y(_16967_));
 AND2x2_ASAP7_75t_R _23676_ (.A(_05837_),
    .B(_05904_),
    .Y(_16968_));
 AND3x1_ASAP7_75t_R _23677_ (.A(_01314_),
    .B(_01874_),
    .C(_15396_),
    .Y(_05911_));
 AO21x2_ASAP7_75t_R _23678_ (.A1(_04965_),
    .A2(_05824_),
    .B(_05911_),
    .Y(_05912_));
 TAPCELL_ASAP7_75t_R TAP_974 ();
 TAPCELL_ASAP7_75t_R TAP_973 ();
 NAND2x1_ASAP7_75t_R _23681_ (.A(net2224),
    .B(_05912_),
    .Y(_16976_));
 TAPCELL_ASAP7_75t_R TAP_972 ();
 OAI22x1_ASAP7_75t_R _23683_ (.A1(_00718_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01242_),
    .Y(_17963_));
 NAND2x1_ASAP7_75t_R _23684_ (.A(net2338),
    .B(_05900_),
    .Y(_16995_));
 NAND2x1_ASAP7_75t_R _23685_ (.A(_05870_),
    .B(_05874_),
    .Y(_17003_));
 AND2x4_ASAP7_75t_R _23686_ (.A(_05849_),
    .B(_05894_),
    .Y(_17008_));
 AND2x4_ASAP7_75t_R _23687_ (.A(_05852_),
    .B(_05904_),
    .Y(_17009_));
 AND2x2_ASAP7_75t_R _23688_ (.A(_05837_),
    .B(_05912_),
    .Y(_17007_));
 AND3x1_ASAP7_75t_R _23689_ (.A(_01314_),
    .B(_01874_),
    .C(_14783_),
    .Y(_05916_));
 AO21x2_ASAP7_75t_R _23690_ (.A1(_05075_),
    .A2(_05824_),
    .B(_05916_),
    .Y(_05917_));
 TAPCELL_ASAP7_75t_R TAP_971 ();
 TAPCELL_ASAP7_75t_R TAP_970 ();
 NAND2x1_ASAP7_75t_R _23693_ (.A(net2223),
    .B(_05917_),
    .Y(_17017_));
 TAPCELL_ASAP7_75t_R TAP_969 ();
 OAI22x1_ASAP7_75t_R _23695_ (.A1(_00750_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01274_),
    .Y(_17979_));
 OR2x2_ASAP7_75t_R _23696_ (.A(_15723_),
    .B(_05819_),
    .Y(_05921_));
 OAI21x1_ASAP7_75t_R _23697_ (.A1(_05355_),
    .A2(_05813_),
    .B(_05921_),
    .Y(_05922_));
 TAPCELL_ASAP7_75t_R TAP_968 ();
 NAND2x1_ASAP7_75t_R _23699_ (.A(_05827_),
    .B(_05922_),
    .Y(_17030_));
 NAND2x1_ASAP7_75t_R _23700_ (.A(net2345),
    .B(_05900_),
    .Y(_17036_));
 NAND2x1_ASAP7_75t_R _23701_ (.A(_05874_),
    .B(net2354),
    .Y(_17046_));
 AND2x2_ASAP7_75t_R _23702_ (.A(net2206),
    .B(_05904_),
    .Y(_17049_));
 AND2x2_ASAP7_75t_R _23703_ (.A(net2234),
    .B(net2270),
    .Y(_17051_));
 AND2x2_ASAP7_75t_R _23704_ (.A(net2295),
    .B(_05917_),
    .Y(_17050_));
 AO22x2_ASAP7_75t_R _23705_ (.A1(_05150_),
    .A2(_05161_),
    .B1(_05172_),
    .B2(_05181_),
    .Y(_05924_));
 AO21x1_ASAP7_75t_R _23706_ (.A1(_01314_),
    .A2(_01874_),
    .B(_05924_),
    .Y(_05925_));
 OA21x2_ASAP7_75t_R _23707_ (.A1(_14099_),
    .A2(_05824_),
    .B(_05925_),
    .Y(_05926_));
 TAPCELL_ASAP7_75t_R TAP_967 ();
 TAPCELL_ASAP7_75t_R TAP_966 ();
 NAND2x1_ASAP7_75t_R _23710_ (.A(net2223),
    .B(_05926_),
    .Y(_17063_));
 OAI22x1_ASAP7_75t_R _23711_ (.A1(_00783_),
    .A2(_05548_),
    .B1(_05817_),
    .B2(_01308_),
    .Y(_17995_));
 AO21x1_ASAP7_75t_R _23712_ (.A1(_15807_),
    .A2(_15838_),
    .B(_05819_),
    .Y(_05929_));
 OA21x2_ASAP7_75t_R _23713_ (.A1(_05454_),
    .A2(_05813_),
    .B(_05929_),
    .Y(_05930_));
 TAPCELL_ASAP7_75t_R TAP_965 ();
 AND2x2_ASAP7_75t_R _23715_ (.A(_05827_),
    .B(_05930_),
    .Y(_17996_));
 AND2x2_ASAP7_75t_R _23716_ (.A(_05840_),
    .B(_05922_),
    .Y(_17078_));
 NOR2x1_ASAP7_75t_R _23717_ (.A(_15590_),
    .B(_05819_),
    .Y(_05932_));
 AO21x2_ASAP7_75t_R _23718_ (.A1(_05244_),
    .A2(_05819_),
    .B(_05932_),
    .Y(_05933_));
 TAPCELL_ASAP7_75t_R TAP_964 ();
 TAPCELL_ASAP7_75t_R TAP_963 ();
 AND2x2_ASAP7_75t_R _23721_ (.A(net2339),
    .B(_05933_),
    .Y(_17079_));
 AND2x2_ASAP7_75t_R _23722_ (.A(net2348),
    .B(_05908_),
    .Y(_17080_));
 NAND2x1_ASAP7_75t_R _23723_ (.A(net2286),
    .B(_05900_),
    .Y(_17084_));
 NAND2x1_ASAP7_75t_R _23724_ (.A(_05874_),
    .B(net2318),
    .Y(_17093_));
 AND2x2_ASAP7_75t_R _23725_ (.A(net2206),
    .B(net2271),
    .Y(_17096_));
 AND2x2_ASAP7_75t_R _23726_ (.A(net2234),
    .B(_05917_),
    .Y(_17097_));
 AND2x2_ASAP7_75t_R _23727_ (.A(net2295),
    .B(_05926_),
    .Y(_17098_));
 NOR2x2_ASAP7_75t_R _23728_ (.A(_05270_),
    .B(_05291_),
    .Y(_05936_));
 AND3x1_ASAP7_75t_R _23729_ (.A(_01314_),
    .B(_01874_),
    .C(_15643_),
    .Y(_05937_));
 AO21x2_ASAP7_75t_R _23730_ (.A1(_05936_),
    .A2(_05824_),
    .B(_05937_),
    .Y(_05938_));
 TAPCELL_ASAP7_75t_R TAP_962 ();
 TAPCELL_ASAP7_75t_R TAP_961 ();
 NAND2x1_ASAP7_75t_R _23733_ (.A(net2226),
    .B(_05938_),
    .Y(_17108_));
 TAPCELL_ASAP7_75t_R TAP_960 ();
 AND3x1_ASAP7_75t_R _23735_ (.A(_13483_),
    .B(_00283_),
    .C(_13484_),
    .Y(_05942_));
 OA21x2_ASAP7_75t_R _23736_ (.A1(_13571_),
    .A2(_05942_),
    .B(_13817_),
    .Y(_05943_));
 AND2x6_ASAP7_75t_R _23737_ (.A(_05454_),
    .B(_05943_),
    .Y(_05944_));
 TAPCELL_ASAP7_75t_R TAP_959 ();
 NAND2x2_ASAP7_75t_R _23739_ (.A(_05819_),
    .B(_05944_),
    .Y(_05946_));
 TAPCELL_ASAP7_75t_R TAP_958 ();
 AND2x2_ASAP7_75t_R _23741_ (.A(_05840_),
    .B(_05930_),
    .Y(_17125_));
 AND2x2_ASAP7_75t_R _23742_ (.A(net2339),
    .B(_05922_),
    .Y(_17126_));
 AND2x2_ASAP7_75t_R _23743_ (.A(net2348),
    .B(_05933_),
    .Y(_17127_));
 NAND2x1_ASAP7_75t_R _23744_ (.A(net2286),
    .B(_05908_),
    .Y(_17132_));
 TAPCELL_ASAP7_75t_R TAP_957 ();
 NAND2x1_ASAP7_75t_R _23746_ (.A(net2190),
    .B(net2318),
    .Y(_17141_));
 AND2x2_ASAP7_75t_R _23747_ (.A(_05859_),
    .B(net2271),
    .Y(_17146_));
 AND2x2_ASAP7_75t_R _23748_ (.A(net2207),
    .B(_05917_),
    .Y(_17147_));
 AND2x2_ASAP7_75t_R _23749_ (.A(net2234),
    .B(_05926_),
    .Y(_17148_));
 NAND2x1_ASAP7_75t_R _23750_ (.A(net2295),
    .B(_05938_),
    .Y(_17158_));
 TAPCELL_ASAP7_75t_R TAP_956 ();
 NAND2x1_ASAP7_75t_R _23752_ (.A(_00281_),
    .B(_13546_),
    .Y(_05949_));
 AOI21x1_ASAP7_75t_R _23753_ (.A1(_13485_),
    .A2(_05949_),
    .B(_13538_),
    .Y(_05950_));
 AND3x4_ASAP7_75t_R _23754_ (.A(_05513_),
    .B(_05824_),
    .C(_05950_),
    .Y(_05951_));
 TAPCELL_ASAP7_75t_R TAP_955 ();
 TAPCELL_ASAP7_75t_R TAP_954 ();
 NAND2x2_ASAP7_75t_R _23757_ (.A(net2245),
    .B(_05951_),
    .Y(_17213_));
 INVx2_ASAP7_75t_R _23758_ (.A(_17213_),
    .Y(_17166_));
 OA22x2_ASAP7_75t_R _23759_ (.A1(_01314_),
    .A2(_00034_),
    .B1(_05548_),
    .B2(_00849_),
    .Y(_17176_));
 AND2x2_ASAP7_75t_R _23760_ (.A(net2348),
    .B(_05922_),
    .Y(_17181_));
 AND2x2_ASAP7_75t_R _23761_ (.A(net2286),
    .B(_05933_),
    .Y(_17182_));
 AND2x2_ASAP7_75t_R _23762_ (.A(net2349),
    .B(_05908_),
    .Y(_17183_));
 NAND2x1_ASAP7_75t_R _23763_ (.A(net2355),
    .B(_05900_),
    .Y(_17187_));
 NAND2x1_ASAP7_75t_R _23764_ (.A(_05874_),
    .B(net2324),
    .Y(_17198_));
 AND2x2_ASAP7_75t_R _23765_ (.A(net2207),
    .B(_05926_),
    .Y(_17203_));
 AND2x2_ASAP7_75t_R _23766_ (.A(net2234),
    .B(_05938_),
    .Y(_17204_));
 AO21x1_ASAP7_75t_R _23767_ (.A1(_01314_),
    .A2(_01874_),
    .B(_05400_),
    .Y(_05954_));
 OA21x2_ASAP7_75t_R _23768_ (.A1(_15773_),
    .A2(_05824_),
    .B(_05954_),
    .Y(_05955_));
 TAPCELL_ASAP7_75t_R TAP_953 ();
 AND2x2_ASAP7_75t_R _23770_ (.A(net2295),
    .B(_05955_),
    .Y(_17205_));
 AO22x2_ASAP7_75t_R _23771_ (.A1(_15853_),
    .A2(_15862_),
    .B1(_15873_),
    .B2(_15884_),
    .Y(_05957_));
 AO21x1_ASAP7_75t_R _23772_ (.A1(_01314_),
    .A2(_01874_),
    .B(_05513_),
    .Y(_05958_));
 OA21x2_ASAP7_75t_R _23773_ (.A1(_05957_),
    .A2(_05824_),
    .B(_05958_),
    .Y(_05959_));
 TAPCELL_ASAP7_75t_R TAP_952 ();
 TAPCELL_ASAP7_75t_R TAP_951 ();
 NAND2x1_ASAP7_75t_R _23776_ (.A(net2225),
    .B(_05959_),
    .Y(_17214_));
 OR3x4_ASAP7_75t_R _23777_ (.A(_13372_),
    .B(_13419_),
    .C(_13441_),
    .Y(_05962_));
 NOR2x1_ASAP7_75t_R _23778_ (.A(_16087_),
    .B(_05813_),
    .Y(_05963_));
 AO21x2_ASAP7_75t_R _23779_ (.A1(_05962_),
    .A2(_05813_),
    .B(_05963_),
    .Y(_05964_));
 TAPCELL_ASAP7_75t_R TAP_950 ();
 NAND2x1_ASAP7_75t_R _23781_ (.A(_05951_),
    .B(net2185),
    .Y(_17215_));
 INVx1_ASAP7_75t_R _23782_ (.A(_17215_),
    .Y(_17262_));
 AO21x2_ASAP7_75t_R _23783_ (.A1(_13485_),
    .A2(_05949_),
    .B(_13538_),
    .Y(_05966_));
 OR3x4_ASAP7_75t_R _23784_ (.A(_01314_),
    .B(_00034_),
    .C(_05966_),
    .Y(_05967_));
 TAPCELL_ASAP7_75t_R TAP_949 ();
 OA21x2_ASAP7_75t_R _23786_ (.A1(_00881_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17226_));
 AND2x2_ASAP7_75t_R _23787_ (.A(net2287),
    .B(_05922_),
    .Y(_17231_));
 AND2x2_ASAP7_75t_R _23788_ (.A(net2349),
    .B(_05933_),
    .Y(_17232_));
 AND2x2_ASAP7_75t_R _23789_ (.A(net2355),
    .B(_05908_),
    .Y(_17233_));
 NAND2x1_ASAP7_75t_R _23790_ (.A(net2318),
    .B(_05900_),
    .Y(_17237_));
 NAND2x1_ASAP7_75t_R _23791_ (.A(_05874_),
    .B(net2271),
    .Y(_17247_));
 NAND2x1_ASAP7_75t_R _23792_ (.A(net2208),
    .B(_05938_),
    .Y(_17252_));
 AND2x2_ASAP7_75t_R _23793_ (.A(net2223),
    .B(_05951_),
    .Y(_17263_));
 OA21x2_ASAP7_75t_R _23794_ (.A1(_00914_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17277_));
 AND2x2_ASAP7_75t_R _23795_ (.A(net2349),
    .B(_05922_),
    .Y(_17282_));
 AND2x2_ASAP7_75t_R _23796_ (.A(net2355),
    .B(_05933_),
    .Y(_17283_));
 AND2x2_ASAP7_75t_R _23797_ (.A(net2318),
    .B(_05908_),
    .Y(_17284_));
 NAND2x1_ASAP7_75t_R _23798_ (.A(net2365),
    .B(_05900_),
    .Y(_17288_));
 NAND2x1_ASAP7_75t_R _23799_ (.A(_05874_),
    .B(_05917_),
    .Y(_17298_));
 TAPCELL_ASAP7_75t_R TAP_948 ();
 NAND2x1_ASAP7_75t_R _23801_ (.A(net2207),
    .B(_05955_),
    .Y(_17303_));
 NAND2x2_ASAP7_75t_R _23802_ (.A(net2295),
    .B(_05951_),
    .Y(_17305_));
 INVx1_ASAP7_75t_R _23803_ (.A(_17305_),
    .Y(_17392_));
 OA21x2_ASAP7_75t_R _23804_ (.A1(_00946_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17321_));
 AND2x2_ASAP7_75t_R _23805_ (.A(net2355),
    .B(_05922_),
    .Y(_17326_));
 AND2x2_ASAP7_75t_R _23806_ (.A(net2318),
    .B(_05933_),
    .Y(_17327_));
 AND2x2_ASAP7_75t_R _23807_ (.A(net2365),
    .B(_05908_),
    .Y(_17328_));
 NAND2x1_ASAP7_75t_R _23808_ (.A(_05900_),
    .B(net2326),
    .Y(_17332_));
 NAND2x1_ASAP7_75t_R _23809_ (.A(_05874_),
    .B(_05926_),
    .Y(_17342_));
 NAND2x1_ASAP7_75t_R _23810_ (.A(net2207),
    .B(_05959_),
    .Y(_17347_));
 NAND2x1_ASAP7_75t_R _23811_ (.A(net2234),
    .B(_05951_),
    .Y(_17348_));
 INVx1_ASAP7_75t_R _23812_ (.A(_17348_),
    .Y(_17393_));
 OA21x2_ASAP7_75t_R _23813_ (.A1(_00979_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17365_));
 NAND2x1_ASAP7_75t_R _23814_ (.A(net2319),
    .B(_05922_),
    .Y(_17370_));
 NAND2x1_ASAP7_75t_R _23815_ (.A(_05900_),
    .B(net2272),
    .Y(_17377_));
 NAND2x1_ASAP7_75t_R _23816_ (.A(_05874_),
    .B(net2308),
    .Y(_17387_));
 AND2x2_ASAP7_75t_R _23817_ (.A(net2207),
    .B(_05951_),
    .Y(_17394_));
 TAPCELL_ASAP7_75t_R TAP_947 ();
 OA21x2_ASAP7_75t_R _23819_ (.A1(_01011_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17413_));
 NAND2x1_ASAP7_75t_R _23820_ (.A(net2368),
    .B(_05922_),
    .Y(_17418_));
 NAND2x1_ASAP7_75t_R _23821_ (.A(_05900_),
    .B(_05917_),
    .Y(_17425_));
 NAND2x1_ASAP7_75t_R _23822_ (.A(_05874_),
    .B(_05955_),
    .Y(_17434_));
 NAND2x2_ASAP7_75t_R _23823_ (.A(_05859_),
    .B(_05951_),
    .Y(_17436_));
 INVx1_ASAP7_75t_R _23824_ (.A(_17436_),
    .Y(_17513_));
 OA21x2_ASAP7_75t_R _23825_ (.A1(_01045_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17456_));
 NAND2x1_ASAP7_75t_R _23826_ (.A(net2328),
    .B(_05922_),
    .Y(_17461_));
 NAND2x1_ASAP7_75t_R _23827_ (.A(_05900_),
    .B(_05926_),
    .Y(_17468_));
 NAND2x1_ASAP7_75t_R _23828_ (.A(_05874_),
    .B(_05959_),
    .Y(_17477_));
 NAND2x1_ASAP7_75t_R _23829_ (.A(_05867_),
    .B(_05951_),
    .Y(_17478_));
 INVx1_ASAP7_75t_R _23830_ (.A(_17478_),
    .Y(_17514_));
 OA21x2_ASAP7_75t_R _23831_ (.A1(_01077_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17492_));
 NAND2x1_ASAP7_75t_R _23832_ (.A(net2274),
    .B(_05922_),
    .Y(_17497_));
 NAND2x1_ASAP7_75t_R _23833_ (.A(_05900_),
    .B(net2309),
    .Y(_17504_));
 AND2x2_ASAP7_75t_R _23834_ (.A(_05874_),
    .B(_05951_),
    .Y(_17515_));
 OA21x2_ASAP7_75t_R _23835_ (.A1(_01110_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17534_));
 NAND2x1_ASAP7_75t_R _23836_ (.A(_05917_),
    .B(_05922_),
    .Y(_17539_));
 NAND2x1_ASAP7_75t_R _23837_ (.A(_05900_),
    .B(_05955_),
    .Y(_17546_));
 NAND2x2_ASAP7_75t_R _23838_ (.A(net2190),
    .B(_05951_),
    .Y(_17548_));
 INVx1_ASAP7_75t_R _23839_ (.A(_17548_),
    .Y(_17612_));
 OA21x2_ASAP7_75t_R _23840_ (.A1(_01142_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17568_));
 NAND2x1_ASAP7_75t_R _23841_ (.A(_05922_),
    .B(_05926_),
    .Y(_17573_));
 NAND2x1_ASAP7_75t_R _23842_ (.A(_05900_),
    .B(_05959_),
    .Y(_17580_));
 NOR2x1_ASAP7_75t_R _23843_ (.A(_14651_),
    .B(_05819_),
    .Y(_05971_));
 AO21x2_ASAP7_75t_R _23844_ (.A1(_04916_),
    .A2(_05819_),
    .B(_05971_),
    .Y(_05972_));
 TAPCELL_ASAP7_75t_R TAP_946 ();
 NAND2x1_ASAP7_75t_R _23846_ (.A(_05951_),
    .B(_05972_),
    .Y(_17581_));
 INVx1_ASAP7_75t_R _23847_ (.A(_17581_),
    .Y(_17613_));
 OA21x2_ASAP7_75t_R _23848_ (.A1(_01176_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17600_));
 NAND2x1_ASAP7_75t_R _23849_ (.A(_05922_),
    .B(net2305),
    .Y(_17605_));
 AND2x2_ASAP7_75t_R _23850_ (.A(_05900_),
    .B(_05951_),
    .Y(_17614_));
 OA21x2_ASAP7_75t_R _23851_ (.A1(_01208_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17630_));
 NAND2x1_ASAP7_75t_R _23852_ (.A(_05922_),
    .B(_05955_),
    .Y(_17635_));
 NAND2x2_ASAP7_75t_R _23853_ (.A(_05908_),
    .B(_05951_),
    .Y(_17637_));
 INVx1_ASAP7_75t_R _23854_ (.A(_17637_),
    .Y(_17684_));
 OA21x2_ASAP7_75t_R _23855_ (.A1(_01242_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17658_));
 NAND2x1_ASAP7_75t_R _23856_ (.A(_05922_),
    .B(_05959_),
    .Y(_17663_));
 NAND2x1_ASAP7_75t_R _23857_ (.A(_05933_),
    .B(_05951_),
    .Y(_17664_));
 INVx1_ASAP7_75t_R _23858_ (.A(_17664_),
    .Y(_17685_));
 OA21x2_ASAP7_75t_R _23859_ (.A1(_01274_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17680_));
 AND2x2_ASAP7_75t_R _23860_ (.A(_05922_),
    .B(_05951_),
    .Y(_17686_));
 OA21x2_ASAP7_75t_R _23861_ (.A1(_01308_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17710_));
 OA21x2_ASAP7_75t_R _23862_ (.A1(_01677_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_17735_));
 INVx1_ASAP7_75t_R _23863_ (.A(_17868_),
    .Y(_16773_));
 OA21x2_ASAP7_75t_R _23864_ (.A1(_01375_),
    .A2(_16773_),
    .B(_01386_),
    .Y(_05974_));
 OA21x2_ASAP7_75t_R _23865_ (.A1(_01385_),
    .A2(_05974_),
    .B(_02313_),
    .Y(_05975_));
 AND3x1_ASAP7_75t_R _23866_ (.A(_01427_),
    .B(_02326_),
    .C(_02322_),
    .Y(_05976_));
 OA211x2_ASAP7_75t_R _23867_ (.A1(_01398_),
    .A2(_05975_),
    .B(_05976_),
    .C(_01411_),
    .Y(_05977_));
 AO21x1_ASAP7_75t_R _23868_ (.A1(net2334),
    .A2(_02322_),
    .B(_01420_),
    .Y(_05978_));
 AO21x1_ASAP7_75t_R _23869_ (.A1(_01427_),
    .A2(_05978_),
    .B(_01426_),
    .Y(_05979_));
 AO21x1_ASAP7_75t_R _23870_ (.A1(_02326_),
    .A2(_05979_),
    .B(_01432_),
    .Y(_05980_));
 OA21x2_ASAP7_75t_R _23871_ (.A1(_05977_),
    .A2(_05980_),
    .B(_01437_),
    .Y(_05981_));
 OA21x2_ASAP7_75t_R _23872_ (.A1(_01436_),
    .A2(_05981_),
    .B(_02330_),
    .Y(_05982_));
 OR3x1_ASAP7_75t_R _23873_ (.A(_00015_),
    .B(_00009_),
    .C(_00019_),
    .Y(_05983_));
 OR2x2_ASAP7_75t_R _23874_ (.A(_00015_),
    .B(_00016_),
    .Y(_05984_));
 AO21x1_ASAP7_75t_R _23875_ (.A1(_02336_),
    .A2(_05984_),
    .B(_00019_),
    .Y(_05985_));
 AND3x1_ASAP7_75t_R _23876_ (.A(_00025_),
    .B(_00032_),
    .C(_02342_),
    .Y(_05986_));
 OA211x2_ASAP7_75t_R _23877_ (.A1(_05982_),
    .A2(_05983_),
    .B(_05985_),
    .C(_05986_),
    .Y(_05987_));
 AND3x1_ASAP7_75t_R _23878_ (.A(_00024_),
    .B(_00032_),
    .C(_02342_),
    .Y(_05988_));
 AO21x1_ASAP7_75t_R _23879_ (.A1(_00032_),
    .A2(_00029_),
    .B(_05988_),
    .Y(_05989_));
 OR3x1_ASAP7_75t_R _23880_ (.A(_00031_),
    .B(net2163),
    .C(_00036_),
    .Y(_05990_));
 OR3x1_ASAP7_75t_R _23881_ (.A(net2163),
    .B(_00036_),
    .C(_02344_),
    .Y(_05991_));
 OA21x2_ASAP7_75t_R _23882_ (.A1(net2164),
    .A2(_00039_),
    .B(_05991_),
    .Y(_05992_));
 OA31x2_ASAP7_75t_R _23883_ (.A1(_05987_),
    .A2(_05989_),
    .A3(_05990_),
    .B1(_05992_),
    .Y(_05993_));
 AND3x1_ASAP7_75t_R _23884_ (.A(_00045_),
    .B(_02347_),
    .C(_02350_),
    .Y(_05994_));
 AND3x1_ASAP7_75t_R _23885_ (.A(_00045_),
    .B(_00041_),
    .C(_02350_),
    .Y(_05995_));
 AO21x1_ASAP7_75t_R _23886_ (.A1(_00044_),
    .A2(_02350_),
    .B(_05995_),
    .Y(_05996_));
 AO21x1_ASAP7_75t_R _23887_ (.A1(_05993_),
    .A2(_05994_),
    .B(_05996_),
    .Y(_05997_));
 OR3x1_ASAP7_75t_R _23888_ (.A(net2134),
    .B(_00049_),
    .C(_00054_),
    .Y(_05998_));
 OR2x2_ASAP7_75t_R _23889_ (.A(_00052_),
    .B(_00053_),
    .Y(_05999_));
 AO21x1_ASAP7_75t_R _23890_ (.A1(_02353_),
    .A2(_05999_),
    .B(_00054_),
    .Y(_06000_));
 OA21x2_ASAP7_75t_R _23891_ (.A1(_05997_),
    .A2(_05998_),
    .B(_06000_),
    .Y(_06001_));
 AND3x1_ASAP7_75t_R _23892_ (.A(_00056_),
    .B(_00059_),
    .C(_02354_),
    .Y(_06002_));
 AND3x1_ASAP7_75t_R _23893_ (.A(_00055_),
    .B(_00059_),
    .C(_02354_),
    .Y(_06003_));
 AO221x1_ASAP7_75t_R _23894_ (.A1(_00059_),
    .A2(_00057_),
    .B1(_06001_),
    .B2(_06002_),
    .C(_06003_),
    .Y(_06004_));
 OA21x2_ASAP7_75t_R _23895_ (.A1(_00058_),
    .A2(_06004_),
    .B(_02355_),
    .Y(_06005_));
 OA21x2_ASAP7_75t_R _23896_ (.A1(_00060_),
    .A2(_06005_),
    .B(_00062_),
    .Y(_06006_));
 OA21x2_ASAP7_75t_R _23897_ (.A1(_00061_),
    .A2(_06006_),
    .B(_02356_),
    .Y(_06007_));
 OA21x2_ASAP7_75t_R _23898_ (.A1(_00063_),
    .A2(_06007_),
    .B(_00065_),
    .Y(_06008_));
 OA21x2_ASAP7_75t_R _23899_ (.A1(_00064_),
    .A2(_06008_),
    .B(_00067_),
    .Y(_17750_));
 INVx13_ASAP7_75t_R _23900_ (.A(net2126),
    .Y(_17486_));
 CKINVDCx12_ASAP7_75t_R _23901_ (.A(net2160),
    .Y(_17526_));
 INVx1_ASAP7_75t_R _23902_ (.A(_02357_),
    .Y(_18324_));
 INVx1_ASAP7_75t_R _23903_ (.A(_02064_),
    .Y(\cs_registers_i.mhpmcounter[2][34] ));
 INVx1_ASAP7_75t_R _23904_ (.A(_02170_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[34] ));
 INVx1_ASAP7_75t_R _23905_ (.A(_01486_),
    .Y(\cs_registers_i.mhpmcounter[2][2] ));
 INVx1_ASAP7_75t_R _23906_ (.A(_01517_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[2] ));
 INVx1_ASAP7_75t_R _23907_ (.A(_02062_),
    .Y(\cs_registers_i.mhpmcounter[2][36] ));
 INVx1_ASAP7_75t_R _23908_ (.A(_02168_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[36] ));
 INVx1_ASAP7_75t_R _23909_ (.A(_01484_),
    .Y(\cs_registers_i.mhpmcounter[2][4] ));
 INVx1_ASAP7_75t_R _23910_ (.A(_01515_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[4] ));
 INVx1_ASAP7_75t_R _23911_ (.A(_02060_),
    .Y(\cs_registers_i.mhpmcounter[2][38] ));
 INVx1_ASAP7_75t_R _23912_ (.A(_02166_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[38] ));
 INVx1_ASAP7_75t_R _23913_ (.A(_01482_),
    .Y(\cs_registers_i.mhpmcounter[2][6] ));
 INVx1_ASAP7_75t_R _23914_ (.A(_01513_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[6] ));
 INVx1_ASAP7_75t_R _23915_ (.A(_02058_),
    .Y(\cs_registers_i.mhpmcounter[2][40] ));
 INVx1_ASAP7_75t_R _23916_ (.A(_02164_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[40] ));
 INVx1_ASAP7_75t_R _23917_ (.A(_01480_),
    .Y(\cs_registers_i.mhpmcounter[2][8] ));
 INVx1_ASAP7_75t_R _23918_ (.A(_01511_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[8] ));
 INVx1_ASAP7_75t_R _23919_ (.A(_02056_),
    .Y(\cs_registers_i.mhpmcounter[2][42] ));
 INVx1_ASAP7_75t_R _23920_ (.A(_02162_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[42] ));
 INVx1_ASAP7_75t_R _23921_ (.A(_01478_),
    .Y(\cs_registers_i.mhpmcounter[2][10] ));
 INVx1_ASAP7_75t_R _23922_ (.A(_01509_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[10] ));
 INVx1_ASAP7_75t_R _23923_ (.A(_02052_),
    .Y(\cs_registers_i.mhpmcounter[2][46] ));
 INVx1_ASAP7_75t_R _23924_ (.A(_02158_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[46] ));
 INVx1_ASAP7_75t_R _23925_ (.A(_01474_),
    .Y(\cs_registers_i.mhpmcounter[2][14] ));
 INVx1_ASAP7_75t_R _23926_ (.A(_01505_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[14] ));
 INVx1_ASAP7_75t_R _23927_ (.A(_02050_),
    .Y(\cs_registers_i.mhpmcounter[2][48] ));
 INVx1_ASAP7_75t_R _23928_ (.A(_02156_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[48] ));
 INVx1_ASAP7_75t_R _23929_ (.A(_01472_),
    .Y(\cs_registers_i.mhpmcounter[2][16] ));
 INVx1_ASAP7_75t_R _23930_ (.A(_01503_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[16] ));
 INVx1_ASAP7_75t_R _23931_ (.A(_02048_),
    .Y(\cs_registers_i.mhpmcounter[2][50] ));
 INVx1_ASAP7_75t_R _23932_ (.A(_02154_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[50] ));
 INVx1_ASAP7_75t_R _23933_ (.A(_01470_),
    .Y(\cs_registers_i.mhpmcounter[2][18] ));
 INVx1_ASAP7_75t_R _23934_ (.A(_01501_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[18] ));
 INVx1_ASAP7_75t_R _23935_ (.A(_02046_),
    .Y(\cs_registers_i.mhpmcounter[2][52] ));
 INVx1_ASAP7_75t_R _23936_ (.A(_02152_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[52] ));
 INVx1_ASAP7_75t_R _23937_ (.A(_01468_),
    .Y(\cs_registers_i.mhpmcounter[2][20] ));
 INVx1_ASAP7_75t_R _23938_ (.A(_01499_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[20] ));
 INVx1_ASAP7_75t_R _23939_ (.A(_02044_),
    .Y(\cs_registers_i.mhpmcounter[2][54] ));
 INVx1_ASAP7_75t_R _23940_ (.A(_02150_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[54] ));
 INVx1_ASAP7_75t_R _23941_ (.A(_01466_),
    .Y(\cs_registers_i.mhpmcounter[2][22] ));
 INVx1_ASAP7_75t_R _23942_ (.A(_01497_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[22] ));
 INVx1_ASAP7_75t_R _23943_ (.A(_02042_),
    .Y(\cs_registers_i.mhpmcounter[2][56] ));
 INVx1_ASAP7_75t_R _23944_ (.A(_02148_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[56] ));
 INVx1_ASAP7_75t_R _23945_ (.A(_01464_),
    .Y(\cs_registers_i.mhpmcounter[2][24] ));
 INVx1_ASAP7_75t_R _23946_ (.A(_01495_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[24] ));
 INVx1_ASAP7_75t_R _23947_ (.A(_02040_),
    .Y(\cs_registers_i.mhpmcounter[2][58] ));
 INVx1_ASAP7_75t_R _23948_ (.A(_02146_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[58] ));
 INVx1_ASAP7_75t_R _23949_ (.A(_01462_),
    .Y(\cs_registers_i.mhpmcounter[2][26] ));
 INVx1_ASAP7_75t_R _23950_ (.A(_01493_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[26] ));
 INVx1_ASAP7_75t_R _23951_ (.A(_02038_),
    .Y(\cs_registers_i.mhpmcounter[2][60] ));
 INVx1_ASAP7_75t_R _23952_ (.A(_02144_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[60] ));
 INVx1_ASAP7_75t_R _23953_ (.A(_01460_),
    .Y(\cs_registers_i.mhpmcounter[2][28] ));
 INVx1_ASAP7_75t_R _23954_ (.A(_01491_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[28] ));
 INVx1_ASAP7_75t_R _23955_ (.A(_02036_),
    .Y(\cs_registers_i.mhpmcounter[2][62] ));
 INVx1_ASAP7_75t_R _23956_ (.A(_02142_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[62] ));
 INVx1_ASAP7_75t_R _23957_ (.A(_01458_),
    .Y(\cs_registers_i.mhpmcounter[2][30] ));
 INVx1_ASAP7_75t_R _23958_ (.A(_01489_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[30] ));
 INVx1_ASAP7_75t_R _23959_ (.A(_02391_),
    .Y(_18478_));
 OR3x1_ASAP7_75t_R _23960_ (.A(_01485_),
    .B(_01486_),
    .C(_02391_),
    .Y(_06009_));
 INVx1_ASAP7_75t_R _23961_ (.A(_06009_),
    .Y(_18479_));
 OR5x1_ASAP7_75t_R _23962_ (.A(_01483_),
    .B(_01484_),
    .C(_01485_),
    .D(_01486_),
    .E(_02391_),
    .Y(_06010_));
 INVx1_ASAP7_75t_R _23963_ (.A(_06010_),
    .Y(_18480_));
 OR3x2_ASAP7_75t_R _23964_ (.A(_01481_),
    .B(_01482_),
    .C(_06010_),
    .Y(_06011_));
 INVx1_ASAP7_75t_R _23965_ (.A(_06011_),
    .Y(_18481_));
 OR2x2_ASAP7_75t_R _23966_ (.A(_01479_),
    .B(_01480_),
    .Y(_06012_));
 OR2x2_ASAP7_75t_R _23967_ (.A(_06011_),
    .B(_06012_),
    .Y(_06013_));
 INVx1_ASAP7_75t_R _23968_ (.A(_06013_),
    .Y(_18482_));
 OR2x2_ASAP7_75t_R _23969_ (.A(_01477_),
    .B(_01478_),
    .Y(_06014_));
 OR3x1_ASAP7_75t_R _23970_ (.A(_06011_),
    .B(_06012_),
    .C(_06014_),
    .Y(_06015_));
 INVx1_ASAP7_75t_R _23971_ (.A(_06015_),
    .Y(_18483_));
 OR2x2_ASAP7_75t_R _23972_ (.A(_01475_),
    .B(_01476_),
    .Y(_06016_));
 NOR2x1_ASAP7_75t_R _23973_ (.A(_06015_),
    .B(_06016_),
    .Y(_18484_));
 OR2x2_ASAP7_75t_R _23974_ (.A(_01473_),
    .B(_01474_),
    .Y(_06017_));
 OR5x2_ASAP7_75t_R _23975_ (.A(_06011_),
    .B(_06012_),
    .C(_06014_),
    .D(_06016_),
    .E(_06017_),
    .Y(_06018_));
 INVx1_ASAP7_75t_R _23976_ (.A(_06018_),
    .Y(_18485_));
 OR3x1_ASAP7_75t_R _23977_ (.A(_01471_),
    .B(_01472_),
    .C(_06018_),
    .Y(_06019_));
 INVx1_ASAP7_75t_R _23978_ (.A(_06019_),
    .Y(_18486_));
 OR5x2_ASAP7_75t_R _23979_ (.A(_01469_),
    .B(_01470_),
    .C(_01471_),
    .D(_01472_),
    .E(_06018_),
    .Y(_06020_));
 INVx1_ASAP7_75t_R _23980_ (.A(_06020_),
    .Y(_18487_));
 INVx1_ASAP7_75t_R _23981_ (.A(_01467_),
    .Y(_06021_));
 AND3x1_ASAP7_75t_R _23982_ (.A(_06021_),
    .B(\cs_registers_i.mhpmcounter[2][20] ),
    .C(_18487_),
    .Y(_18488_));
 OR5x2_ASAP7_75t_R _23983_ (.A(_01465_),
    .B(_01466_),
    .C(_01467_),
    .D(_01468_),
    .E(_06020_),
    .Y(_06022_));
 INVx1_ASAP7_75t_R _23984_ (.A(_06022_),
    .Y(_18489_));
 OR3x1_ASAP7_75t_R _23985_ (.A(_01463_),
    .B(_01464_),
    .C(_06022_),
    .Y(_06023_));
 INVx1_ASAP7_75t_R _23986_ (.A(_06023_),
    .Y(_18490_));
 OR5x1_ASAP7_75t_R _23987_ (.A(_01461_),
    .B(_01462_),
    .C(_01463_),
    .D(_01464_),
    .E(_06022_),
    .Y(_06024_));
 INVx1_ASAP7_75t_R _23988_ (.A(_06024_),
    .Y(_18491_));
 INVx1_ASAP7_75t_R _23989_ (.A(_01459_),
    .Y(_06025_));
 AND3x1_ASAP7_75t_R _23990_ (.A(_06025_),
    .B(\cs_registers_i.mhpmcounter[2][28] ),
    .C(_18491_),
    .Y(_18492_));
 OR5x1_ASAP7_75t_R _23991_ (.A(_01457_),
    .B(_01458_),
    .C(_01459_),
    .D(_01460_),
    .E(_06024_),
    .Y(_06026_));
 INVx1_ASAP7_75t_R _23992_ (.A(_06026_),
    .Y(_18493_));
 INVx1_ASAP7_75t_R _23993_ (.A(_02065_),
    .Y(_06027_));
 AND3x1_ASAP7_75t_R _23994_ (.A(_06027_),
    .B(\cs_registers_i.mhpmcounter[2][32] ),
    .C(_18493_),
    .Y(_18494_));
 OR5x2_ASAP7_75t_R _23995_ (.A(_02063_),
    .B(_02064_),
    .C(_02065_),
    .D(_02066_),
    .E(_06026_),
    .Y(_06028_));
 INVx1_ASAP7_75t_R _23996_ (.A(_06028_),
    .Y(_18495_));
 INVx1_ASAP7_75t_R _23997_ (.A(_02061_),
    .Y(_06029_));
 AND3x1_ASAP7_75t_R _23998_ (.A(_06029_),
    .B(\cs_registers_i.mhpmcounter[2][36] ),
    .C(_18495_),
    .Y(_18496_));
 OR5x2_ASAP7_75t_R _23999_ (.A(_02059_),
    .B(_02060_),
    .C(_02061_),
    .D(_02062_),
    .E(_06028_),
    .Y(_06030_));
 INVx1_ASAP7_75t_R _24000_ (.A(_06030_),
    .Y(_18497_));
 OR3x1_ASAP7_75t_R _24001_ (.A(_02057_),
    .B(_02058_),
    .C(_06030_),
    .Y(_06031_));
 INVx1_ASAP7_75t_R _24002_ (.A(_06031_),
    .Y(_18498_));
 OR5x1_ASAP7_75t_R _24003_ (.A(_02055_),
    .B(_02056_),
    .C(_02057_),
    .D(_02058_),
    .E(_06030_),
    .Y(_06032_));
 INVx1_ASAP7_75t_R _24004_ (.A(_06032_),
    .Y(_18499_));
 INVx1_ASAP7_75t_R _24005_ (.A(_02053_),
    .Y(_06033_));
 AND3x1_ASAP7_75t_R _24006_ (.A(_06033_),
    .B(\cs_registers_i.mhpmcounter[2][44] ),
    .C(_18499_),
    .Y(_18500_));
 OR5x1_ASAP7_75t_R _24007_ (.A(_02051_),
    .B(_02052_),
    .C(_02053_),
    .D(_02054_),
    .E(_06032_),
    .Y(_06034_));
 INVx1_ASAP7_75t_R _24008_ (.A(_06034_),
    .Y(_18501_));
 OR3x1_ASAP7_75t_R _24009_ (.A(_02049_),
    .B(_02050_),
    .C(_06034_),
    .Y(_06035_));
 INVx1_ASAP7_75t_R _24010_ (.A(_06035_),
    .Y(_18502_));
 OR3x2_ASAP7_75t_R _24011_ (.A(_02047_),
    .B(_02048_),
    .C(_06035_),
    .Y(_06036_));
 INVx1_ASAP7_75t_R _24012_ (.A(_06036_),
    .Y(_18503_));
 OR3x1_ASAP7_75t_R _24013_ (.A(_02045_),
    .B(_02046_),
    .C(_06036_),
    .Y(_06037_));
 INVx1_ASAP7_75t_R _24014_ (.A(_06037_),
    .Y(_18504_));
 OR5x2_ASAP7_75t_R _24015_ (.A(_02043_),
    .B(_02044_),
    .C(_02045_),
    .D(_02046_),
    .E(_06036_),
    .Y(_06038_));
 INVx1_ASAP7_75t_R _24016_ (.A(_06038_),
    .Y(_18505_));
 OR3x1_ASAP7_75t_R _24017_ (.A(_02041_),
    .B(_02042_),
    .C(_06038_),
    .Y(_06039_));
 INVx1_ASAP7_75t_R _24018_ (.A(_06039_),
    .Y(_18506_));
 OR5x2_ASAP7_75t_R _24019_ (.A(_02039_),
    .B(_02040_),
    .C(_02041_),
    .D(_02042_),
    .E(_06038_),
    .Y(_06040_));
 INVx1_ASAP7_75t_R _24020_ (.A(_06040_),
    .Y(_18507_));
 NOR3x1_ASAP7_75t_R _24021_ (.A(_02037_),
    .B(_02038_),
    .C(_06040_),
    .Y(_18508_));
 INVx1_ASAP7_75t_R _24022_ (.A(_02455_),
    .Y(_18509_));
 OR3x1_ASAP7_75t_R _24023_ (.A(_01516_),
    .B(_01517_),
    .C(_02455_),
    .Y(_06041_));
 INVx1_ASAP7_75t_R _24024_ (.A(_06041_),
    .Y(_18510_));
 OR5x2_ASAP7_75t_R _24025_ (.A(_01514_),
    .B(_01515_),
    .C(_01516_),
    .D(_01517_),
    .E(_02455_),
    .Y(_06042_));
 INVx1_ASAP7_75t_R _24026_ (.A(_06042_),
    .Y(_18511_));
 OR2x2_ASAP7_75t_R _24027_ (.A(_01512_),
    .B(_01513_),
    .Y(_06043_));
 OR2x2_ASAP7_75t_R _24028_ (.A(_06042_),
    .B(_06043_),
    .Y(_06044_));
 INVx1_ASAP7_75t_R _24029_ (.A(_06044_),
    .Y(_18512_));
 OR2x2_ASAP7_75t_R _24030_ (.A(_01510_),
    .B(_01511_),
    .Y(_06045_));
 OR3x1_ASAP7_75t_R _24031_ (.A(_06042_),
    .B(_06043_),
    .C(_06045_),
    .Y(_06046_));
 INVx1_ASAP7_75t_R _24032_ (.A(_06046_),
    .Y(_18513_));
 OR2x2_ASAP7_75t_R _24033_ (.A(_01508_),
    .B(_01509_),
    .Y(_06047_));
 OR2x2_ASAP7_75t_R _24034_ (.A(_06046_),
    .B(_06047_),
    .Y(_06048_));
 INVx1_ASAP7_75t_R _24035_ (.A(_06048_),
    .Y(_18514_));
 OR2x2_ASAP7_75t_R _24036_ (.A(_01506_),
    .B(_01507_),
    .Y(_06049_));
 OR5x2_ASAP7_75t_R _24037_ (.A(_06042_),
    .B(_06043_),
    .C(_06045_),
    .D(_06047_),
    .E(_06049_),
    .Y(_06050_));
 INVx1_ASAP7_75t_R _24038_ (.A(_06050_),
    .Y(_18515_));
 OR2x2_ASAP7_75t_R _24039_ (.A(_01504_),
    .B(_01505_),
    .Y(_06051_));
 OR2x2_ASAP7_75t_R _24040_ (.A(_06050_),
    .B(_06051_),
    .Y(_06052_));
 INVx1_ASAP7_75t_R _24041_ (.A(_06052_),
    .Y(_18516_));
 OR2x2_ASAP7_75t_R _24042_ (.A(_01502_),
    .B(_01503_),
    .Y(_06053_));
 OR3x1_ASAP7_75t_R _24043_ (.A(_06050_),
    .B(_06051_),
    .C(_06053_),
    .Y(_06054_));
 INVx1_ASAP7_75t_R _24044_ (.A(_06054_),
    .Y(_18517_));
 OR2x2_ASAP7_75t_R _24045_ (.A(_01500_),
    .B(_01501_),
    .Y(_06055_));
 OR2x2_ASAP7_75t_R _24046_ (.A(_06054_),
    .B(_06055_),
    .Y(_06056_));
 INVx1_ASAP7_75t_R _24047_ (.A(_06056_),
    .Y(_18518_));
 OR2x2_ASAP7_75t_R _24048_ (.A(_01498_),
    .B(_01499_),
    .Y(_06057_));
 OR5x2_ASAP7_75t_R _24049_ (.A(_06050_),
    .B(_06051_),
    .C(_06053_),
    .D(_06055_),
    .E(_06057_),
    .Y(_06058_));
 INVx1_ASAP7_75t_R _24050_ (.A(_06058_),
    .Y(_18519_));
 OR2x2_ASAP7_75t_R _24051_ (.A(_01496_),
    .B(_01497_),
    .Y(_06059_));
 OR2x2_ASAP7_75t_R _24052_ (.A(_06058_),
    .B(_06059_),
    .Y(_06060_));
 INVx1_ASAP7_75t_R _24053_ (.A(_06060_),
    .Y(_18520_));
 OR4x2_ASAP7_75t_R _24054_ (.A(_01494_),
    .B(_01495_),
    .C(_06058_),
    .D(_06059_),
    .Y(_06061_));
 INVx1_ASAP7_75t_R _24055_ (.A(_06061_),
    .Y(_18521_));
 OR2x2_ASAP7_75t_R _24056_ (.A(_01492_),
    .B(_01493_),
    .Y(_06062_));
 OR2x2_ASAP7_75t_R _24057_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 INVx1_ASAP7_75t_R _24058_ (.A(_06063_),
    .Y(_18522_));
 OR2x2_ASAP7_75t_R _24059_ (.A(_01490_),
    .B(_01491_),
    .Y(_06064_));
 NOR2x1_ASAP7_75t_R _24060_ (.A(_06063_),
    .B(_06064_),
    .Y(_18523_));
 OR5x2_ASAP7_75t_R _24061_ (.A(_01488_),
    .B(_01489_),
    .C(_06061_),
    .D(_06062_),
    .E(_06064_),
    .Y(_06065_));
 TAPCELL_ASAP7_75t_R TAP_945 ();
 INVx1_ASAP7_75t_R _24063_ (.A(_06065_),
    .Y(_18524_));
 OR3x1_ASAP7_75t_R _24064_ (.A(_02171_),
    .B(_02172_),
    .C(_06065_),
    .Y(_06067_));
 INVx1_ASAP7_75t_R _24065_ (.A(_06067_),
    .Y(_18525_));
 OR4x2_ASAP7_75t_R _24066_ (.A(_02169_),
    .B(_02170_),
    .C(_02171_),
    .D(_02172_),
    .Y(_06068_));
 NOR2x1_ASAP7_75t_R _24067_ (.A(_06065_),
    .B(_06068_),
    .Y(_18526_));
 OR3x2_ASAP7_75t_R _24068_ (.A(_02167_),
    .B(_02168_),
    .C(_06068_),
    .Y(_06069_));
 NOR2x1_ASAP7_75t_R _24069_ (.A(_06065_),
    .B(_06069_),
    .Y(_18527_));
 OR2x2_ASAP7_75t_R _24070_ (.A(_02165_),
    .B(_02166_),
    .Y(_06070_));
 NOR3x1_ASAP7_75t_R _24071_ (.A(_06065_),
    .B(_06069_),
    .C(_06070_),
    .Y(_18528_));
 INVx1_ASAP7_75t_R _24072_ (.A(_02163_),
    .Y(_06071_));
 AND3x1_ASAP7_75t_R _24073_ (.A(_06071_),
    .B(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .C(_18528_),
    .Y(_18529_));
 INVx1_ASAP7_75t_R _24074_ (.A(_02161_),
    .Y(_06072_));
 AND3x1_ASAP7_75t_R _24075_ (.A(_06072_),
    .B(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .C(_18529_),
    .Y(_18530_));
 NOR2x1_ASAP7_75t_R _24076_ (.A(_02159_),
    .B(_02160_),
    .Y(_06073_));
 NAND2x1_ASAP7_75t_R _24077_ (.A(_18530_),
    .B(_06073_),
    .Y(_06074_));
 INVx1_ASAP7_75t_R _24078_ (.A(_06074_),
    .Y(_18531_));
 INVx1_ASAP7_75t_R _24079_ (.A(_02157_),
    .Y(_06075_));
 AND3x1_ASAP7_75t_R _24080_ (.A(_06075_),
    .B(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .C(_18531_),
    .Y(_18532_));
 OR5x2_ASAP7_75t_R _24081_ (.A(_02155_),
    .B(_02156_),
    .C(_02157_),
    .D(_02158_),
    .E(_06074_),
    .Y(_06076_));
 INVx1_ASAP7_75t_R _24082_ (.A(_06076_),
    .Y(_18533_));
 OR3x1_ASAP7_75t_R _24083_ (.A(_02153_),
    .B(_02154_),
    .C(_06076_),
    .Y(_06077_));
 INVx1_ASAP7_75t_R _24084_ (.A(_06077_),
    .Y(_18534_));
 OR3x4_ASAP7_75t_R _24085_ (.A(_02151_),
    .B(_02152_),
    .C(_06077_),
    .Y(_06078_));
 INVx1_ASAP7_75t_R _24086_ (.A(_06078_),
    .Y(_18535_));
 NOR3x2_ASAP7_75t_R _24087_ (.B(_02150_),
    .C(_06078_),
    .Y(_18536_),
    .A(_02149_));
 INVx1_ASAP7_75t_R _24088_ (.A(_02147_),
    .Y(_06079_));
 AND3x1_ASAP7_75t_R _24089_ (.A(_06079_),
    .B(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .C(_18536_),
    .Y(_18537_));
 INVx1_ASAP7_75t_R _24090_ (.A(_02145_),
    .Y(_06080_));
 AND3x1_ASAP7_75t_R _24091_ (.A(_06080_),
    .B(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .C(_18537_),
    .Y(_18538_));
 INVx1_ASAP7_75t_R _24092_ (.A(_02143_),
    .Y(_06081_));
 AND3x1_ASAP7_75t_R _24093_ (.A(_06081_),
    .B(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .C(_18538_),
    .Y(_18539_));
 INVx1_ASAP7_75t_R _24094_ (.A(_01606_),
    .Y(\cs_registers_i.pc_if_i[3] ));
 INVx1_ASAP7_75t_R _24095_ (.A(_01604_),
    .Y(\cs_registers_i.pc_if_i[5] ));
 INVx2_ASAP7_75t_R _24096_ (.A(_01602_),
    .Y(\cs_registers_i.pc_if_i[7] ));
 INVx1_ASAP7_75t_R _24097_ (.A(_01600_),
    .Y(\cs_registers_i.pc_if_i[9] ));
 INVx1_ASAP7_75t_R _24098_ (.A(_01598_),
    .Y(\cs_registers_i.pc_if_i[11] ));
 INVx2_ASAP7_75t_R _24099_ (.A(_01596_),
    .Y(\cs_registers_i.pc_if_i[13] ));
 INVx2_ASAP7_75t_R _24100_ (.A(_01594_),
    .Y(\cs_registers_i.pc_if_i[15] ));
 INVx2_ASAP7_75t_R _24101_ (.A(_01592_),
    .Y(\cs_registers_i.pc_if_i[17] ));
 INVx2_ASAP7_75t_R _24102_ (.A(_01590_),
    .Y(\cs_registers_i.pc_if_i[19] ));
 INVx2_ASAP7_75t_R _24103_ (.A(_01588_),
    .Y(\cs_registers_i.pc_if_i[21] ));
 INVx2_ASAP7_75t_R _24104_ (.A(_01586_),
    .Y(\cs_registers_i.pc_if_i[23] ));
 INVx2_ASAP7_75t_R _24105_ (.A(_01584_),
    .Y(\cs_registers_i.pc_if_i[25] ));
 INVx2_ASAP7_75t_R _24106_ (.A(_01582_),
    .Y(\cs_registers_i.pc_if_i[27] ));
 INVx2_ASAP7_75t_R _24107_ (.A(_01580_),
    .Y(\cs_registers_i.pc_if_i[29] ));
 INVx1_ASAP7_75t_R _24108_ (.A(_02519_),
    .Y(_18540_));
 OR3x1_ASAP7_75t_R _24109_ (.A(_00170_),
    .B(_00174_),
    .C(_02519_),
    .Y(_06082_));
 INVx1_ASAP7_75t_R _24110_ (.A(_06082_),
    .Y(_18541_));
 OR5x1_ASAP7_75t_R _24111_ (.A(_00170_),
    .B(_00174_),
    .C(_00177_),
    .D(_00180_),
    .E(_02519_),
    .Y(_06083_));
 INVx1_ASAP7_75t_R _24112_ (.A(_06083_),
    .Y(_18542_));
 OR3x1_ASAP7_75t_R _24113_ (.A(_00182_),
    .B(_00186_),
    .C(_06083_),
    .Y(_06084_));
 INVx1_ASAP7_75t_R _24114_ (.A(_06084_),
    .Y(_18543_));
 OR3x1_ASAP7_75t_R _24115_ (.A(_00189_),
    .B(_00193_),
    .C(_06084_),
    .Y(_06085_));
 INVx1_ASAP7_75t_R _24116_ (.A(_06085_),
    .Y(_18544_));
 OR5x1_ASAP7_75t_R _24117_ (.A(_00189_),
    .B(_00193_),
    .C(_00196_),
    .D(_00199_),
    .E(_06084_),
    .Y(_06086_));
 INVx1_ASAP7_75t_R _24118_ (.A(_06086_),
    .Y(_18545_));
 OR3x1_ASAP7_75t_R _24119_ (.A(_00201_),
    .B(_00204_),
    .C(_06086_),
    .Y(_06087_));
 INVx1_ASAP7_75t_R _24120_ (.A(_06087_),
    .Y(_18546_));
 OR3x1_ASAP7_75t_R _24121_ (.A(_00206_),
    .B(_00208_),
    .C(_06087_),
    .Y(_06088_));
 INVx1_ASAP7_75t_R _24122_ (.A(_06088_),
    .Y(_18547_));
 OR3x1_ASAP7_75t_R _24123_ (.A(_00209_),
    .B(_00211_),
    .C(_06088_),
    .Y(_06089_));
 INVx1_ASAP7_75t_R _24124_ (.A(_06089_),
    .Y(_18548_));
 OR3x1_ASAP7_75t_R _24125_ (.A(_00212_),
    .B(_00214_),
    .C(_06089_),
    .Y(_06090_));
 INVx1_ASAP7_75t_R _24126_ (.A(_06090_),
    .Y(_18549_));
 OR3x1_ASAP7_75t_R _24127_ (.A(_00215_),
    .B(_00217_),
    .C(_06090_),
    .Y(_06091_));
 INVx1_ASAP7_75t_R _24128_ (.A(_06091_),
    .Y(_18550_));
 OR3x1_ASAP7_75t_R _24129_ (.A(_00218_),
    .B(_00220_),
    .C(_06091_),
    .Y(_06092_));
 INVx1_ASAP7_75t_R _24130_ (.A(_06092_),
    .Y(_18551_));
 OR3x1_ASAP7_75t_R _24131_ (.A(_00221_),
    .B(_00223_),
    .C(_06092_),
    .Y(_06093_));
 INVx1_ASAP7_75t_R _24132_ (.A(_06093_),
    .Y(_18552_));
 OR3x1_ASAP7_75t_R _24133_ (.A(_00224_),
    .B(_00226_),
    .C(_06093_),
    .Y(_06094_));
 INVx1_ASAP7_75t_R _24134_ (.A(_06094_),
    .Y(_18553_));
 TAPCELL_ASAP7_75t_R TAP_944 ();
 TAPCELL_ASAP7_75t_R TAP_943 ();
 TAPCELL_ASAP7_75t_R TAP_942 ();
 TAPCELL_ASAP7_75t_R TAP_941 ();
 TAPCELL_ASAP7_75t_R TAP_940 ();
 TAPCELL_ASAP7_75t_R TAP_939 ();
 TAPCELL_ASAP7_75t_R TAP_938 ();
 TAPCELL_ASAP7_75t_R TAP_937 ();
 OA222x2_ASAP7_75t_R _24143_ (.A1(_00231_),
    .A2(_15972_),
    .B1(_04698_),
    .B2(_00232_),
    .C1(net294),
    .C2(_14540_),
    .Y(_06103_));
 NAND2x1_ASAP7_75t_R _24144_ (.A(net292),
    .B(_06103_),
    .Y(_06104_));
 OA21x2_ASAP7_75t_R _24145_ (.A1(net292),
    .A2(_13886_),
    .B(_06104_),
    .Y(net186));
 TAPCELL_ASAP7_75t_R TAP_936 ();
 CKINVDCx10_ASAP7_75t_R _24147_ (.A(net294),
    .Y(_06106_));
 NAND2x1_ASAP7_75t_R _24148_ (.A(_06106_),
    .B(_14597_),
    .Y(_06107_));
 OA211x2_ASAP7_75t_R _24149_ (.A1(_00231_),
    .A2(_16087_),
    .B(_06107_),
    .C(net292),
    .Y(_06108_));
 OAI21x1_ASAP7_75t_R _24150_ (.A1(_00232_),
    .A2(_04808_),
    .B(_06108_),
    .Y(_06109_));
 OA21x2_ASAP7_75t_R _24151_ (.A1(net292),
    .A2(_05962_),
    .B(_06109_),
    .Y(net197));
 INVx8_ASAP7_75t_R _24152_ (.A(_00231_),
    .Y(_06110_));
 TAPCELL_ASAP7_75t_R TAP_935 ();
 CKINVDCx8_ASAP7_75t_R _24154_ (.A(_00232_),
    .Y(_06112_));
 TAPCELL_ASAP7_75t_R TAP_934 ();
 CKINVDCx16_ASAP7_75t_R _24156_ (.A(_18555_),
    .Y(_06114_));
 AO21x1_ASAP7_75t_R _24157_ (.A1(_06106_),
    .A2(_14652_),
    .B(_06114_),
    .Y(_06115_));
 AO221x1_ASAP7_75t_R _24158_ (.A1(_06110_),
    .A2(_16213_),
    .B1(_04916_),
    .B2(_06112_),
    .C(_06115_),
    .Y(_06116_));
 OA21x2_ASAP7_75t_R _24159_ (.A1(net291),
    .A2(_14169_),
    .B(_06116_),
    .Y(net208));
 AOI22x1_ASAP7_75t_R _24160_ (.A1(_06106_),
    .A2(_05898_),
    .B1(_16324_),
    .B2(_06110_),
    .Y(_06117_));
 OA211x2_ASAP7_75t_R _24161_ (.A1(_00232_),
    .A2(_05028_),
    .B(_06117_),
    .C(net291),
    .Y(_06118_));
 INVx1_ASAP7_75t_R _24162_ (.A(_06118_),
    .Y(_06119_));
 OA21x2_ASAP7_75t_R _24163_ (.A1(net291),
    .A2(net2231),
    .B(_06119_),
    .Y(net211));
 OA222x2_ASAP7_75t_R _24164_ (.A1(_00231_),
    .A2(_16457_),
    .B1(_05136_),
    .B2(_00232_),
    .C1(net294),
    .C2(_15488_),
    .Y(_06120_));
 NAND2x1_ASAP7_75t_R _24165_ (.A(net292),
    .B(_06120_),
    .Y(_06121_));
 OA21x2_ASAP7_75t_R _24166_ (.A1(net292),
    .A2(net2218),
    .B(_06121_),
    .Y(net212));
 OA222x2_ASAP7_75t_R _24167_ (.A1(_00231_),
    .A2(net2182),
    .B1(_05245_),
    .B2(_00232_),
    .C1(net294),
    .C2(_15590_),
    .Y(_06122_));
 NAND2x1_ASAP7_75t_R _24168_ (.A(net291),
    .B(_06122_),
    .Y(_06123_));
 OA21x2_ASAP7_75t_R _24169_ (.A1(net291),
    .A2(_14355_),
    .B(_06123_),
    .Y(net213));
 OA222x2_ASAP7_75t_R _24170_ (.A1(_00231_),
    .A2(_16679_),
    .B1(_05355_),
    .B2(_00232_),
    .C1(net294),
    .C2(_15723_),
    .Y(_06124_));
 NAND2x1_ASAP7_75t_R _24171_ (.A(net292),
    .B(_06124_),
    .Y(_06125_));
 OA21x2_ASAP7_75t_R _24172_ (.A1(net292),
    .A2(_14420_),
    .B(_06125_),
    .Y(net214));
 TAPCELL_ASAP7_75t_R TAP_933 ();
 INVx1_ASAP7_75t_R _24174_ (.A(_05454_),
    .Y(_06127_));
 OA222x2_ASAP7_75t_R _24175_ (.A1(_00231_),
    .A2(_04577_),
    .B1(_06127_),
    .B2(_00232_),
    .C1(net294),
    .C2(_15839_),
    .Y(_06128_));
 NAND2x1_ASAP7_75t_R _24176_ (.A(net292),
    .B(_06128_),
    .Y(_06129_));
 OA21x2_ASAP7_75t_R _24177_ (.A1(net292),
    .A2(_14479_),
    .B(_06129_),
    .Y(net215));
 OAI21x1_ASAP7_75t_R _24178_ (.A1(net294),
    .A2(_15972_),
    .B(net291),
    .Y(_06130_));
 AO221x1_ASAP7_75t_R _24179_ (.A1(_06112_),
    .A2(_13886_),
    .B1(_04697_),
    .B2(_06110_),
    .C(_06130_),
    .Y(_06131_));
 OA21x2_ASAP7_75t_R _24180_ (.A1(net291),
    .A2(_14539_),
    .B(_06131_),
    .Y(net216));
 OA22x2_ASAP7_75t_R _24181_ (.A1(net294),
    .A2(_16087_),
    .B1(_04808_),
    .B2(_00231_),
    .Y(_06132_));
 OA211x2_ASAP7_75t_R _24182_ (.A1(_00232_),
    .A2(_13442_),
    .B(_06132_),
    .C(net292),
    .Y(_06133_));
 INVx1_ASAP7_75t_R _24183_ (.A(_06133_),
    .Y(_06134_));
 OA21x2_ASAP7_75t_R _24184_ (.A1(net291),
    .A2(_14597_),
    .B(_06134_),
    .Y(net217));
 TAPCELL_ASAP7_75t_R TAP_932 ();
 TAPCELL_ASAP7_75t_R TAP_931 ();
 AO21x1_ASAP7_75t_R _24187_ (.A1(_06112_),
    .A2(_14169_),
    .B(_06114_),
    .Y(_06137_));
 AO221x1_ASAP7_75t_R _24188_ (.A1(_06106_),
    .A2(_16213_),
    .B1(_04916_),
    .B2(_06110_),
    .C(_06137_),
    .Y(_06138_));
 OA21x2_ASAP7_75t_R _24189_ (.A1(net291),
    .A2(_14652_),
    .B(_06138_),
    .Y(net187));
 TAPCELL_ASAP7_75t_R TAP_930 ();
 TAPCELL_ASAP7_75t_R TAP_929 ();
 AOI22x1_ASAP7_75t_R _24192_ (.A1(_06112_),
    .A2(net2231),
    .B1(_16324_),
    .B2(_06106_),
    .Y(_06141_));
 OA211x2_ASAP7_75t_R _24193_ (.A1(_00231_),
    .A2(_05028_),
    .B(_06141_),
    .C(net291),
    .Y(_06142_));
 AOI21x1_ASAP7_75t_R _24194_ (.A1(_06114_),
    .A2(_14703_),
    .B(_06142_),
    .Y(net188));
 AO221x1_ASAP7_75t_R _24195_ (.A1(_06112_),
    .A2(net2218),
    .B1(_16456_),
    .B2(_06106_),
    .C(_06114_),
    .Y(_06143_));
 AND3x1_ASAP7_75t_R _24196_ (.A(_06110_),
    .B(_05104_),
    .C(_05135_),
    .Y(_06144_));
 OA22x2_ASAP7_75t_R _24197_ (.A1(net291),
    .A2(_15487_),
    .B1(_06143_),
    .B2(_06144_),
    .Y(net189));
 INVx1_ASAP7_75t_R _24198_ (.A(_14355_),
    .Y(_06145_));
 OA222x2_ASAP7_75t_R _24199_ (.A1(_00232_),
    .A2(_06145_),
    .B1(net2183),
    .B2(net294),
    .C1(_05245_),
    .C2(_00231_),
    .Y(_06146_));
 OR2x2_ASAP7_75t_R _24200_ (.A(net291),
    .B(_15590_),
    .Y(_06147_));
 OAI21x1_ASAP7_75t_R _24201_ (.A1(_06114_),
    .A2(_06146_),
    .B(_06147_),
    .Y(net190));
 INVx1_ASAP7_75t_R _24202_ (.A(_16679_),
    .Y(_06148_));
 AO32x1_ASAP7_75t_R _24203_ (.A1(_06110_),
    .A2(_05323_),
    .A3(_05354_),
    .B1(_06106_),
    .B2(_06148_),
    .Y(_06149_));
 AO21x1_ASAP7_75t_R _24204_ (.A1(_06112_),
    .A2(_14420_),
    .B(_06149_),
    .Y(_06150_));
 NOR2x1_ASAP7_75t_R _24205_ (.A(net292),
    .B(_15723_),
    .Y(_06151_));
 AO21x1_ASAP7_75t_R _24206_ (.A1(net292),
    .A2(_06150_),
    .B(_06151_),
    .Y(net191));
 AO221x1_ASAP7_75t_R _24207_ (.A1(_06112_),
    .A2(_14479_),
    .B1(_05454_),
    .B2(_06110_),
    .C(_06114_),
    .Y(_06152_));
 AOI21x1_ASAP7_75t_R _24208_ (.A1(_06106_),
    .A2(_04576_),
    .B(_06152_),
    .Y(_06153_));
 AOI21x1_ASAP7_75t_R _24209_ (.A1(_06114_),
    .A2(_15839_),
    .B(_06153_),
    .Y(net192));
 AO222x2_ASAP7_75t_R _24210_ (.A1(_06110_),
    .A2(_13886_),
    .B1(_14539_),
    .B2(_06112_),
    .C1(_04697_),
    .C2(_06106_),
    .Y(_06154_));
 AND3x1_ASAP7_75t_R _24211_ (.A(_06114_),
    .B(_15933_),
    .C(_15971_),
    .Y(_06155_));
 AO21x1_ASAP7_75t_R _24212_ (.A1(net291),
    .A2(_06154_),
    .B(_06155_),
    .Y(net193));
 AOI22x1_ASAP7_75t_R _24213_ (.A1(_06110_),
    .A2(_05962_),
    .B1(_14597_),
    .B2(_06112_),
    .Y(_06156_));
 OA211x2_ASAP7_75t_R _24214_ (.A1(net294),
    .A2(_04808_),
    .B(_06156_),
    .C(net292),
    .Y(_06157_));
 AOI21x1_ASAP7_75t_R _24215_ (.A1(_06114_),
    .A2(_16087_),
    .B(_06157_),
    .Y(net194));
 AO21x1_ASAP7_75t_R _24216_ (.A1(_06112_),
    .A2(_14652_),
    .B(_06114_),
    .Y(_06158_));
 AO221x1_ASAP7_75t_R _24217_ (.A1(_06110_),
    .A2(_14169_),
    .B1(_04916_),
    .B2(_06106_),
    .C(_06158_),
    .Y(_06159_));
 OA21x2_ASAP7_75t_R _24218_ (.A1(net291),
    .A2(_16213_),
    .B(_06159_),
    .Y(net195));
 AOI22x1_ASAP7_75t_R _24219_ (.A1(_06110_),
    .A2(net2231),
    .B1(_05898_),
    .B2(_06112_),
    .Y(_06160_));
 OA211x2_ASAP7_75t_R _24220_ (.A1(net294),
    .A2(_05028_),
    .B(_06160_),
    .C(net291),
    .Y(_06161_));
 AOI21x1_ASAP7_75t_R _24221_ (.A1(_06114_),
    .A2(_16329_),
    .B(_06161_),
    .Y(net196));
 INVx1_ASAP7_75t_R _24222_ (.A(net2220),
    .Y(_06162_));
 OA222x2_ASAP7_75t_R _24223_ (.A1(_00231_),
    .A2(_06162_),
    .B1(_15488_),
    .B2(_00232_),
    .C1(_05136_),
    .C2(net294),
    .Y(_06163_));
 NAND2x1_ASAP7_75t_R _24224_ (.A(net291),
    .B(_06163_),
    .Y(_06164_));
 OA21x2_ASAP7_75t_R _24225_ (.A1(net291),
    .A2(_16456_),
    .B(_06164_),
    .Y(net198));
 OA222x2_ASAP7_75t_R _24226_ (.A1(_00231_),
    .A2(_06145_),
    .B1(_15590_),
    .B2(_00232_),
    .C1(_05245_),
    .C2(net294),
    .Y(_06165_));
 OR2x2_ASAP7_75t_R _24227_ (.A(net291),
    .B(net2184),
    .Y(_06166_));
 OAI21x1_ASAP7_75t_R _24228_ (.A1(_06114_),
    .A2(_06165_),
    .B(_06166_),
    .Y(net199));
 OAI22x1_ASAP7_75t_R _24229_ (.A1(_00232_),
    .A2(_15723_),
    .B1(_05355_),
    .B2(net294),
    .Y(_06167_));
 AO21x1_ASAP7_75t_R _24230_ (.A1(_06110_),
    .A2(_14420_),
    .B(_06167_),
    .Y(_06168_));
 AND3x1_ASAP7_75t_R _24231_ (.A(_06114_),
    .B(_16647_),
    .C(_16678_),
    .Y(_06169_));
 AO21x1_ASAP7_75t_R _24232_ (.A1(net292),
    .A2(_06168_),
    .B(_06169_),
    .Y(net200));
 AOI22x1_ASAP7_75t_R _24233_ (.A1(_06110_),
    .A2(_14479_),
    .B1(_05454_),
    .B2(_06106_),
    .Y(_06170_));
 OA211x2_ASAP7_75t_R _24234_ (.A1(_00232_),
    .A2(_15839_),
    .B(_06170_),
    .C(net292),
    .Y(_06171_));
 AOI21x1_ASAP7_75t_R _24235_ (.A1(_06114_),
    .A2(_04577_),
    .B(_06171_),
    .Y(net201));
 OAI21x1_ASAP7_75t_R _24236_ (.A1(_00232_),
    .A2(_15972_),
    .B(net291),
    .Y(_06172_));
 AO221x1_ASAP7_75t_R _24237_ (.A1(_06106_),
    .A2(_13886_),
    .B1(_14539_),
    .B2(_06110_),
    .C(_06172_),
    .Y(_06173_));
 OA21x2_ASAP7_75t_R _24238_ (.A1(net291),
    .A2(_04697_),
    .B(_06173_),
    .Y(net202));
 AOI22x1_ASAP7_75t_R _24239_ (.A1(_06106_),
    .A2(_05962_),
    .B1(_14597_),
    .B2(_06110_),
    .Y(_06174_));
 OA211x2_ASAP7_75t_R _24240_ (.A1(_00232_),
    .A2(_16087_),
    .B(_06174_),
    .C(net292),
    .Y(_06175_));
 AOI21x1_ASAP7_75t_R _24241_ (.A1(_06114_),
    .A2(_04808_),
    .B(_06175_),
    .Y(net203));
 AO21x1_ASAP7_75t_R _24242_ (.A1(_06110_),
    .A2(_14652_),
    .B(_06114_),
    .Y(_06176_));
 AO221x1_ASAP7_75t_R _24243_ (.A1(_06106_),
    .A2(_14169_),
    .B1(_16213_),
    .B2(_06112_),
    .C(_06176_),
    .Y(_06177_));
 OA21x2_ASAP7_75t_R _24244_ (.A1(net291),
    .A2(_04916_),
    .B(_06177_),
    .Y(net204));
 AO222x2_ASAP7_75t_R _24245_ (.A1(_06110_),
    .A2(_05898_),
    .B1(_16324_),
    .B2(_06112_),
    .C1(_06106_),
    .C2(net2231),
    .Y(_06178_));
 AND3x1_ASAP7_75t_R _24246_ (.A(_06114_),
    .B(_04995_),
    .C(_05027_),
    .Y(_06179_));
 AO21x1_ASAP7_75t_R _24247_ (.A1(net291),
    .A2(_06178_),
    .B(_06179_),
    .Y(net205));
 AO222x2_ASAP7_75t_R _24248_ (.A1(_06110_),
    .A2(_15487_),
    .B1(_16456_),
    .B2(_06112_),
    .C1(_06106_),
    .C2(net2219),
    .Y(_06180_));
 AND3x1_ASAP7_75t_R _24249_ (.A(_06114_),
    .B(_05104_),
    .C(_05135_),
    .Y(_06181_));
 AO21x1_ASAP7_75t_R _24250_ (.A1(net291),
    .A2(_06180_),
    .B(_06181_),
    .Y(net206));
 OA222x2_ASAP7_75t_R _24251_ (.A1(_00231_),
    .A2(_15590_),
    .B1(net2182),
    .B2(_00232_),
    .C1(net294),
    .C2(_06145_),
    .Y(_06182_));
 NOR2x1_ASAP7_75t_R _24252_ (.A(_06114_),
    .B(_06182_),
    .Y(_06183_));
 AO21x1_ASAP7_75t_R _24253_ (.A1(_06114_),
    .A2(_05244_),
    .B(_06183_),
    .Y(net207));
 OAI22x1_ASAP7_75t_R _24254_ (.A1(_00231_),
    .A2(_15723_),
    .B1(_16679_),
    .B2(_00232_),
    .Y(_06184_));
 AO21x1_ASAP7_75t_R _24255_ (.A1(_06106_),
    .A2(_14420_),
    .B(_06184_),
    .Y(_06185_));
 AND3x1_ASAP7_75t_R _24256_ (.A(_06114_),
    .B(_05323_),
    .C(_05354_),
    .Y(_06186_));
 AO21x1_ASAP7_75t_R _24257_ (.A1(net292),
    .A2(_06185_),
    .B(_06186_),
    .Y(net209));
 AOI221x1_ASAP7_75t_R _24258_ (.A1(_06106_),
    .A2(_14479_),
    .B1(_04576_),
    .B2(_06112_),
    .C(_06114_),
    .Y(_06187_));
 OAI21x1_ASAP7_75t_R _24259_ (.A1(_00231_),
    .A2(_15839_),
    .B(_06187_),
    .Y(_06188_));
 OA21x2_ASAP7_75t_R _24260_ (.A1(net292),
    .A2(_05454_),
    .B(_06188_),
    .Y(net210));
 NAND2x2_ASAP7_75t_R _24261_ (.A(_00282_),
    .B(_14828_),
    .Y(_06189_));
 AND2x2_ASAP7_75t_R _24262_ (.A(_13483_),
    .B(_02534_),
    .Y(_06190_));
 AO21x1_ASAP7_75t_R _24263_ (.A1(_00281_),
    .A2(_06114_),
    .B(_06190_),
    .Y(_06191_));
 NAND2x1_ASAP7_75t_R _24264_ (.A(_02535_),
    .B(_06189_),
    .Y(_06192_));
 OA21x2_ASAP7_75t_R _24265_ (.A1(_06189_),
    .A2(_06191_),
    .B(_06192_),
    .Y(net181));
 INVx1_ASAP7_75t_R _24266_ (.A(_02536_),
    .Y(_06193_));
 NAND2x1_ASAP7_75t_R _24267_ (.A(_13483_),
    .B(_00233_),
    .Y(_06194_));
 OA211x2_ASAP7_75t_R _24268_ (.A1(_13483_),
    .A2(_06112_),
    .B(_05763_),
    .C(_06194_),
    .Y(_06195_));
 AO21x2_ASAP7_75t_R _24269_ (.A1(_06193_),
    .A2(_06189_),
    .B(_06195_),
    .Y(net182));
 OR3x1_ASAP7_75t_R _24270_ (.A(_13508_),
    .B(_00281_),
    .C(_00235_),
    .Y(_06196_));
 OAI21x1_ASAP7_75t_R _24271_ (.A1(_13483_),
    .A2(_00231_),
    .B(_06196_),
    .Y(_06197_));
 NAND2x1_ASAP7_75t_R _24272_ (.A(_13508_),
    .B(_02537_),
    .Y(_06198_));
 OA211x2_ASAP7_75t_R _24273_ (.A1(_13508_),
    .A2(_00234_),
    .B(_06189_),
    .C(_06198_),
    .Y(_06199_));
 AO21x2_ASAP7_75t_R _24274_ (.A1(_05763_),
    .A2(_06197_),
    .B(_06199_),
    .Y(net183));
 NAND2x1_ASAP7_75t_R _24275_ (.A(_13483_),
    .B(_00236_),
    .Y(_06200_));
 OA211x2_ASAP7_75t_R _24276_ (.A1(_13483_),
    .A2(_06106_),
    .B(_05763_),
    .C(_06200_),
    .Y(_06201_));
 AO21x2_ASAP7_75t_R _24277_ (.A1(_18554_),
    .A2(_06189_),
    .B(_06201_),
    .Y(net184));
 OA21x2_ASAP7_75t_R _24278_ (.A1(_13444_),
    .A2(_05753_),
    .B(_00277_),
    .Y(net185));
 AO21x1_ASAP7_75t_R _24279_ (.A1(_13496_),
    .A2(_13587_),
    .B(_13518_),
    .Y(_06202_));
 NAND3x1_ASAP7_75t_R _24280_ (.A(_01713_),
    .B(_14797_),
    .C(_06202_),
    .Y(_06203_));
 OA31x2_ASAP7_75t_R _24281_ (.A1(_14821_),
    .A2(_14841_),
    .A3(_06203_),
    .B1(_01710_),
    .Y(_06204_));
 OR2x6_ASAP7_75t_R _24282_ (.A(_01317_),
    .B(_01721_),
    .Y(_06205_));
 NAND2x1_ASAP7_75t_R _24283_ (.A(_14796_),
    .B(_06205_),
    .Y(_06206_));
 AND3x4_ASAP7_75t_R _24284_ (.A(_01719_),
    .B(_01724_),
    .C(_01725_),
    .Y(_06207_));
 NAND2x1_ASAP7_75t_R _24285_ (.A(_17810_),
    .B(_02140_),
    .Y(_06208_));
 OR3x1_ASAP7_75t_R _24286_ (.A(_02030_),
    .B(_17810_),
    .C(_02140_),
    .Y(_06209_));
 OA211x2_ASAP7_75t_R _24287_ (.A1(_02032_),
    .A2(_06208_),
    .B(_06209_),
    .C(_01311_),
    .Y(_06210_));
 NOR2x2_ASAP7_75t_R _24288_ (.A(_01317_),
    .B(_01721_),
    .Y(_06211_));
 OR3x1_ASAP7_75t_R _24289_ (.A(_14803_),
    .B(_06210_),
    .C(_06211_),
    .Y(_06212_));
 TAPCELL_ASAP7_75t_R TAP_928 ();
 INVx2_ASAP7_75t_R _24291_ (.A(_01312_),
    .Y(_06214_));
 NAND2x1_ASAP7_75t_R _24292_ (.A(_01740_),
    .B(_01741_),
    .Y(_06215_));
 OR5x2_ASAP7_75t_R _24293_ (.A(_06214_),
    .B(_06215_),
    .C(_13851_),
    .D(_14808_),
    .E(_05725_),
    .Y(_06216_));
 OR3x4_ASAP7_75t_R _24294_ (.A(_06207_),
    .B(_06212_),
    .C(_06216_),
    .Y(_06217_));
 NAND2x1_ASAP7_75t_R _24295_ (.A(_05557_),
    .B(_06217_),
    .Y(_06218_));
 OR3x4_ASAP7_75t_R _24296_ (.A(_14799_),
    .B(_14806_),
    .C(_05725_),
    .Y(_06219_));
 TAPCELL_ASAP7_75t_R TAP_927 ();
 OR3x4_ASAP7_75t_R _24298_ (.A(_14808_),
    .B(_14799_),
    .C(_05725_),
    .Y(_06221_));
 TAPCELL_ASAP7_75t_R TAP_926 ();
 AND3x1_ASAP7_75t_R _24300_ (.A(_06219_),
    .B(_06221_),
    .C(_06207_),
    .Y(_06223_));
 TAPCELL_ASAP7_75t_R TAP_925 ();
 INVx2_ASAP7_75t_R _24302_ (.A(_01714_),
    .Y(_06225_));
 TAPCELL_ASAP7_75t_R TAP_924 ();
 NAND2x2_ASAP7_75t_R _24304_ (.A(_01715_),
    .B(_01716_),
    .Y(_06227_));
 INVx1_ASAP7_75t_R _24305_ (.A(net3102),
    .Y(_06228_));
 AND2x2_ASAP7_75t_R _24306_ (.A(_06228_),
    .B(_02034_),
    .Y(_06229_));
 NOR2x2_ASAP7_75t_R _24307_ (.A(_01714_),
    .B(_06227_),
    .Y(_06230_));
 INVx1_ASAP7_75t_R _24308_ (.A(_06230_),
    .Y(_06231_));
 AO21x1_ASAP7_75t_R _24309_ (.A1(_01717_),
    .A2(_06229_),
    .B(_06231_),
    .Y(_06232_));
 OA21x2_ASAP7_75t_R _24310_ (.A1(_06225_),
    .A2(_06227_),
    .B(_06232_),
    .Y(_06233_));
 NOR2x2_ASAP7_75t_R _24311_ (.A(_01716_),
    .B(_01717_),
    .Y(_06234_));
 AND3x4_ASAP7_75t_R _24312_ (.A(_01714_),
    .B(_14793_),
    .C(_06234_),
    .Y(_06235_));
 INVx1_ASAP7_75t_R _24313_ (.A(_01453_),
    .Y(_06236_));
 OA211x2_ASAP7_75t_R _24314_ (.A1(net3131),
    .A2(_06236_),
    .B(_01718_),
    .C(_01311_),
    .Y(_06237_));
 AND2x2_ASAP7_75t_R _24315_ (.A(_06235_),
    .B(_06237_),
    .Y(_06238_));
 INVx1_ASAP7_75t_R _24316_ (.A(_01956_),
    .Y(_06239_));
 INVx1_ASAP7_75t_R _24317_ (.A(_01957_),
    .Y(_06240_));
 AO22x2_ASAP7_75t_R _24318_ (.A1(net3492),
    .A2(_06239_),
    .B1(_06240_),
    .B2(net141),
    .Y(_06241_));
 INVx1_ASAP7_75t_R _24319_ (.A(_01958_),
    .Y(_06242_));
 INVx1_ASAP7_75t_R _24320_ (.A(_01959_),
    .Y(_06243_));
 AO22x1_ASAP7_75t_R _24321_ (.A1(net140),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net3497),
    .Y(_06244_));
 INVx1_ASAP7_75t_R _24322_ (.A(_01960_),
    .Y(_06245_));
 INVx1_ASAP7_75t_R _24323_ (.A(_01961_),
    .Y(_06246_));
 AO22x1_ASAP7_75t_R _24324_ (.A1(net138),
    .A2(_06245_),
    .B1(_06246_),
    .B2(net137),
    .Y(_06247_));
 INVx1_ASAP7_75t_R _24325_ (.A(_01962_),
    .Y(_06248_));
 INVx1_ASAP7_75t_R _24326_ (.A(_01963_),
    .Y(_06249_));
 AO22x1_ASAP7_75t_R _24327_ (.A1(net136),
    .A2(_06248_),
    .B1(_06249_),
    .B2(net3299),
    .Y(_06250_));
 OR4x2_ASAP7_75t_R _24328_ (.A(net3493),
    .B(_06244_),
    .C(_06247_),
    .D(net3300),
    .Y(_06251_));
 INVx1_ASAP7_75t_R _24329_ (.A(net3505),
    .Y(_06252_));
 INVx2_ASAP7_75t_R _24330_ (.A(net3407),
    .Y(_06253_));
 OAI22x1_ASAP7_75t_R _24331_ (.A1(_06252_),
    .A2(_01952_),
    .B1(_01953_),
    .B2(net3408),
    .Y(_06254_));
 INVx1_ASAP7_75t_R _24332_ (.A(_01954_),
    .Y(_06255_));
 INVx1_ASAP7_75t_R _24333_ (.A(_01955_),
    .Y(_06256_));
 AO22x1_ASAP7_75t_R _24334_ (.A1(net3477),
    .A2(_06255_),
    .B1(_06256_),
    .B2(net143),
    .Y(_06257_));
 INVx1_ASAP7_75t_R _24335_ (.A(_01949_),
    .Y(_06258_));
 AND2x2_ASAP7_75t_R _24336_ (.A(net3354),
    .B(_06258_),
    .Y(_06259_));
 INVx1_ASAP7_75t_R _24337_ (.A(_01950_),
    .Y(_06260_));
 INVx1_ASAP7_75t_R _24338_ (.A(_01951_),
    .Y(_06261_));
 AO22x1_ASAP7_75t_R _24339_ (.A1(net3387),
    .A2(_06260_),
    .B1(_06261_),
    .B2(net3372),
    .Y(_06262_));
 OR4x2_ASAP7_75t_R _24340_ (.A(net3409),
    .B(_06257_),
    .C(net3355),
    .D(net3373),
    .Y(_06263_));
 INVx1_ASAP7_75t_R _24341_ (.A(net3513),
    .Y(_06264_));
 INVx2_ASAP7_75t_R _24342_ (.A(net3368),
    .Y(_06265_));
 OAI22x1_ASAP7_75t_R _24343_ (.A1(_06264_),
    .A2(_01946_),
    .B1(_01948_),
    .B2(net3369),
    .Y(_06266_));
 INVx1_ASAP7_75t_R _24344_ (.A(_01947_),
    .Y(_06267_));
 AO21x1_ASAP7_75t_R _24345_ (.A1(net3207),
    .A2(_06267_),
    .B(net2643),
    .Y(_06268_));
 OR2x2_ASAP7_75t_R _24346_ (.A(net3370),
    .B(net3208),
    .Y(_06269_));
 OR3x4_ASAP7_75t_R _24347_ (.A(net3301),
    .B(net3356),
    .C(net3209),
    .Y(_06270_));
 NAND2x2_ASAP7_75t_R _24348_ (.A(_06238_),
    .B(net3210),
    .Y(_06271_));
 OA211x2_ASAP7_75t_R _24349_ (.A1(_06218_),
    .A2(_06223_),
    .B(_06233_),
    .C(_06271_),
    .Y(_06272_));
 OA21x2_ASAP7_75t_R _24350_ (.A1(_06204_),
    .A2(_06206_),
    .B(_06272_),
    .Y(_06273_));
 TAPCELL_ASAP7_75t_R TAP_923 ();
 TAPCELL_ASAP7_75t_R TAP_922 ();
 TAPCELL_ASAP7_75t_R TAP_921 ();
 TAPCELL_ASAP7_75t_R TAP_920 ();
 NAND2x1_ASAP7_75t_R _24355_ (.A(net3487),
    .B(_06258_),
    .Y(_06278_));
 NAND2x1_ASAP7_75t_R _24356_ (.A(net3372),
    .B(_06261_),
    .Y(_06279_));
 INVx1_ASAP7_75t_R _24357_ (.A(_01952_),
    .Y(_06280_));
 NAND2x1_ASAP7_75t_R _24358_ (.A(net143),
    .B(_06256_),
    .Y(_06281_));
 NAND2x1_ASAP7_75t_R _24359_ (.A(net141),
    .B(_06240_),
    .Y(_06282_));
 INVx1_ASAP7_75t_R _24360_ (.A(net3497),
    .Y(_06283_));
 NAND2x1_ASAP7_75t_R _24361_ (.A(net137),
    .B(_06246_),
    .Y(_06284_));
 AO32x1_ASAP7_75t_R _24362_ (.A1(net136),
    .A2(_06248_),
    .A3(_06284_),
    .B1(net138),
    .B2(_06245_),
    .Y(_06285_));
 OA21x2_ASAP7_75t_R _24363_ (.A1(_06283_),
    .A2(_01959_),
    .B(_06285_),
    .Y(_06286_));
 AO21x1_ASAP7_75t_R _24364_ (.A1(net140),
    .A2(_06242_),
    .B(_06286_),
    .Y(_06287_));
 AO22x1_ASAP7_75t_R _24365_ (.A1(net142),
    .A2(_06239_),
    .B1(_06282_),
    .B2(_06287_),
    .Y(_06288_));
 AO22x1_ASAP7_75t_R _24366_ (.A1(net144),
    .A2(_06255_),
    .B1(_06281_),
    .B2(_06288_),
    .Y(_06289_));
 OA21x2_ASAP7_75t_R _24367_ (.A1(_06253_),
    .A2(_01953_),
    .B(_06289_),
    .Y(_06290_));
 AO21x1_ASAP7_75t_R _24368_ (.A1(net132),
    .A2(_06280_),
    .B(_06290_),
    .Y(_06291_));
 AO22x1_ASAP7_75t_R _24369_ (.A1(net3387),
    .A2(_06260_),
    .B1(_06279_),
    .B2(_06291_),
    .Y(_06292_));
 NOR2x1_ASAP7_75t_R _24370_ (.A(net3301),
    .B(net3356),
    .Y(_06293_));
 AOI221x1_ASAP7_75t_R _24371_ (.A1(net3131),
    .A2(_01718_),
    .B1(_06278_),
    .B2(net3388),
    .C(_06293_),
    .Y(_06294_));
 OR2x2_ASAP7_75t_R _24372_ (.A(_06271_),
    .B(net3489),
    .Y(_06295_));
 OAI21x1_ASAP7_75t_R _24373_ (.A1(_06204_),
    .A2(_06206_),
    .B(_06272_),
    .Y(_06296_));
 TAPCELL_ASAP7_75t_R TAP_919 ();
 TAPCELL_ASAP7_75t_R TAP_918 ();
 TAPCELL_ASAP7_75t_R TAP_917 ();
 NAND2x2_ASAP7_75t_R _24377_ (.A(_05557_),
    .B(_06207_),
    .Y(_06300_));
 OR2x6_ASAP7_75t_R _24378_ (.A(_06221_),
    .B(_06300_),
    .Y(_06301_));
 TAPCELL_ASAP7_75t_R TAP_916 ();
 TAPCELL_ASAP7_75t_R TAP_915 ();
 NAND2x2_ASAP7_75t_R _24381_ (.A(_14791_),
    .B(_14794_),
    .Y(_06304_));
 TAPCELL_ASAP7_75t_R TAP_914 ();
 TAPCELL_ASAP7_75t_R TAP_913 ();
 TAPCELL_ASAP7_75t_R TAP_912 ();
 OR2x6_ASAP7_75t_R _24385_ (.A(_06219_),
    .B(_06300_),
    .Y(_06308_));
 TAPCELL_ASAP7_75t_R TAP_911 ();
 OA22x2_ASAP7_75t_R _24387_ (.A1(_06304_),
    .A2(_05792_),
    .B1(_06308_),
    .B2(_01575_),
    .Y(_06310_));
 OA21x2_ASAP7_75t_R _24388_ (.A1(_01943_),
    .A2(_06301_),
    .B(_06310_),
    .Y(_06311_));
 AND3x4_ASAP7_75t_R _24389_ (.A(net3390),
    .B(_06296_),
    .C(_06311_),
    .Y(_06312_));
 AOI21x1_ASAP7_75t_R _24390_ (.A1(_01549_),
    .A2(net300),
    .B(net3391),
    .Y(_18605_));
 TAPCELL_ASAP7_75t_R TAP_910 ();
 TAPCELL_ASAP7_75t_R TAP_909 ();
 TAPCELL_ASAP7_75t_R TAP_908 ();
 NOR2x1_ASAP7_75t_R _24394_ (.A(net429),
    .B(_02201_),
    .Y(_06316_));
 AO21x1_ASAP7_75t_R _24395_ (.A1(net429),
    .A2(_18605_),
    .B(_06316_),
    .Y(net239));
 INVx2_ASAP7_75t_R _24396_ (.A(net174),
    .Y(_06317_));
 NAND3x2_ASAP7_75t_R _24397_ (.B(_01724_),
    .C(_01725_),
    .Y(_06318_),
    .A(_01719_));
 NAND2x2_ASAP7_75t_R _24398_ (.A(_05557_),
    .B(_06318_),
    .Y(_06319_));
 OA222x2_ASAP7_75t_R _24399_ (.A1(_06317_),
    .A2(_06304_),
    .B1(_06308_),
    .B2(_00081_),
    .C1(_06319_),
    .C2(_01311_),
    .Y(_06320_));
 AOI22x1_ASAP7_75t_R _24400_ (.A1(net3533),
    .A2(_06242_),
    .B1(_06243_),
    .B2(net3497),
    .Y(_06321_));
 AOI21x1_ASAP7_75t_R _24401_ (.A1(_06321_),
    .A2(_06247_),
    .B(net3493),
    .Y(_06322_));
 OA222x2_ASAP7_75t_R _24402_ (.A1(net3506),
    .A2(_01952_),
    .B1(net3478),
    .B2(_06322_),
    .C1(_01953_),
    .C2(net3408),
    .Y(_06323_));
 AO21x1_ASAP7_75t_R _24403_ (.A1(net3131),
    .A2(_01718_),
    .B(net3355),
    .Y(_06324_));
 NOR2x1_ASAP7_75t_R _24404_ (.A(_06293_),
    .B(_06324_),
    .Y(_06325_));
 OA21x2_ASAP7_75t_R _24405_ (.A1(net3373),
    .A2(net3507),
    .B(_06325_),
    .Y(_06326_));
 NOR2x1_ASAP7_75t_R _24406_ (.A(net3211),
    .B(net3508),
    .Y(_06327_));
 INVx1_ASAP7_75t_R _24407_ (.A(net3509),
    .Y(_06328_));
 OR3x1_ASAP7_75t_R _24408_ (.A(_01942_),
    .B(_06221_),
    .C(_06300_),
    .Y(_06329_));
 AND4x2_ASAP7_75t_R _24409_ (.A(_06296_),
    .B(_06320_),
    .C(net3510),
    .D(_06329_),
    .Y(_06330_));
 AOI21x1_ASAP7_75t_R _24410_ (.A1(_01548_),
    .A2(net300),
    .B(_06330_),
    .Y(_18575_));
 TAPCELL_ASAP7_75t_R TAP_907 ();
 NOR2x1_ASAP7_75t_R _24412_ (.A(net429),
    .B(_02200_),
    .Y(_06332_));
 AO21x1_ASAP7_75t_R _24413_ (.A1(net429),
    .A2(_18575_),
    .B(_06332_),
    .Y(net242));
 TAPCELL_ASAP7_75t_R TAP_906 ();
 OR2x2_ASAP7_75t_R _24415_ (.A(net3409),
    .B(net3478),
    .Y(_06334_));
 NOR2x1_ASAP7_75t_R _24416_ (.A(net3493),
    .B(net3498),
    .Y(_06335_));
 OA21x2_ASAP7_75t_R _24417_ (.A1(net3495),
    .A2(net3370),
    .B(net3499),
    .Y(_06336_));
 NOR2x1_ASAP7_75t_R _24418_ (.A(net3373),
    .B(_06324_),
    .Y(_06337_));
 OA21x2_ASAP7_75t_R _24419_ (.A1(net3479),
    .A2(net3500),
    .B(net3374),
    .Y(_06338_));
 AND2x4_ASAP7_75t_R _24420_ (.A(_05557_),
    .B(_06207_),
    .Y(_06339_));
 OAI22x1_ASAP7_75t_R _24421_ (.A1(_00084_),
    .A2(_05727_),
    .B1(_05728_),
    .B2(_01941_),
    .Y(_06340_));
 AOI22x1_ASAP7_75t_R _24422_ (.A1(_14796_),
    .A2(net175),
    .B1(_06339_),
    .B2(_06340_),
    .Y(_06341_));
 OA21x2_ASAP7_75t_R _24423_ (.A1(net3211),
    .A2(net3502),
    .B(_06341_),
    .Y(_06342_));
 AND2x2_ASAP7_75t_R _24424_ (.A(net299),
    .B(_06342_),
    .Y(_06343_));
 AOI21x1_ASAP7_75t_R _24425_ (.A1(_01547_),
    .A2(net300),
    .B(_06343_),
    .Y(_18577_));
 NOR2x1_ASAP7_75t_R _24426_ (.A(net429),
    .B(_02199_),
    .Y(_06344_));
 AO21x1_ASAP7_75t_R _24427_ (.A1(net429),
    .A2(_18577_),
    .B(_06344_),
    .Y(net243));
 INVx3_ASAP7_75t_R _24428_ (.A(net289),
    .Y(_06345_));
 OA22x2_ASAP7_75t_R _24429_ (.A1(_00087_),
    .A2(_05727_),
    .B1(_05728_),
    .B2(_01940_),
    .Y(_06346_));
 INVx1_ASAP7_75t_R _24430_ (.A(net3479),
    .Y(_06347_));
 OR3x1_ASAP7_75t_R _24431_ (.A(net3369),
    .B(_01948_),
    .C(net3301),
    .Y(_06348_));
 AND3x2_ASAP7_75t_R _24432_ (.A(net3480),
    .B(net3374),
    .C(_06348_),
    .Y(_06349_));
 OR2x2_ASAP7_75t_R _24433_ (.A(_06271_),
    .B(net3481),
    .Y(_06350_));
 OA21x2_ASAP7_75t_R _24434_ (.A1(_06300_),
    .A2(_06346_),
    .B(net3482),
    .Y(_06351_));
 OA211x2_ASAP7_75t_R _24435_ (.A1(_06345_),
    .A2(_06304_),
    .B(_06296_),
    .C(net3483),
    .Y(_06352_));
 AO21x2_ASAP7_75t_R _24436_ (.A1(_01546_),
    .A2(net300),
    .B(_06352_),
    .Y(_06353_));
 INVx4_ASAP7_75t_R _24437_ (.A(net429),
    .Y(_06354_));
 TAPCELL_ASAP7_75t_R TAP_905 ();
 AND2x2_ASAP7_75t_R _24439_ (.A(_06354_),
    .B(_02198_),
    .Y(_06356_));
 AOI21x1_ASAP7_75t_R _24440_ (.A1(net429),
    .A2(_06353_),
    .B(_06356_),
    .Y(net244));
 OA22x2_ASAP7_75t_R _24441_ (.A1(_00090_),
    .A2(_06219_),
    .B1(_06221_),
    .B2(_01939_),
    .Y(_06357_));
 OR3x2_ASAP7_75t_R _24442_ (.A(net3131),
    .B(net3301),
    .C(net3411),
    .Y(_06358_));
 NAND2x1_ASAP7_75t_R _24443_ (.A(_06238_),
    .B(net3412),
    .Y(_06359_));
 OA21x2_ASAP7_75t_R _24444_ (.A1(_06304_),
    .A2(_05793_),
    .B(net3413),
    .Y(_06360_));
 OA21x2_ASAP7_75t_R _24445_ (.A1(_06300_),
    .A2(_06357_),
    .B(_06360_),
    .Y(_06361_));
 AND2x2_ASAP7_75t_R _24446_ (.A(net299),
    .B(_06361_),
    .Y(_06362_));
 AOI21x1_ASAP7_75t_R _24447_ (.A1(_01545_),
    .A2(net300),
    .B(_06362_),
    .Y(_18579_));
 TAPCELL_ASAP7_75t_R TAP_904 ();
 NOR2x1_ASAP7_75t_R _24449_ (.A(net429),
    .B(_02197_),
    .Y(_06364_));
 AO21x1_ASAP7_75t_R _24450_ (.A1(net429),
    .A2(_18579_),
    .B(_06364_),
    .Y(net245));
 TAPCELL_ASAP7_75t_R TAP_903 ();
 NOR2x2_ASAP7_75t_R _24452_ (.A(_06219_),
    .B(_06300_),
    .Y(_06366_));
 INVx1_ASAP7_75t_R _24453_ (.A(_01574_),
    .Y(_06367_));
 AOI22x1_ASAP7_75t_R _24454_ (.A1(net178),
    .A2(_14796_),
    .B1(_06366_),
    .B2(_06367_),
    .Y(_06368_));
 AND2x2_ASAP7_75t_R _24455_ (.A(_01714_),
    .B(_14793_),
    .Y(_06369_));
 AO21x1_ASAP7_75t_R _24456_ (.A1(_05556_),
    .A2(_06318_),
    .B(_14791_),
    .Y(_06370_));
 INVx1_ASAP7_75t_R _24457_ (.A(_14806_),
    .Y(_06371_));
 INVx1_ASAP7_75t_R _24458_ (.A(_05725_),
    .Y(_06372_));
 INVx1_ASAP7_75t_R _24459_ (.A(_14799_),
    .Y(_06373_));
 OA211x2_ASAP7_75t_R _24460_ (.A1(_14813_),
    .A2(_06371_),
    .B(_06372_),
    .C(_06373_),
    .Y(_06374_));
 AO221x2_ASAP7_75t_R _24461_ (.A1(_06369_),
    .A2(_06370_),
    .B1(_06374_),
    .B2(_06339_),
    .C(_06230_),
    .Y(_06375_));
 OA211x2_ASAP7_75t_R _24462_ (.A1(_01938_),
    .A2(_06301_),
    .B(_06368_),
    .C(_06375_),
    .Y(_06376_));
 AND2x2_ASAP7_75t_R _24463_ (.A(net299),
    .B(_06376_),
    .Y(_06377_));
 AO21x1_ASAP7_75t_R _24464_ (.A1(_01544_),
    .A2(net301),
    .B(_06377_),
    .Y(_06378_));
 AND2x2_ASAP7_75t_R _24465_ (.A(_06354_),
    .B(_02196_),
    .Y(_06379_));
 AOI21x1_ASAP7_75t_R _24466_ (.A1(net429),
    .A2(_06378_),
    .B(_06379_),
    .Y(net246));
 AOI221x1_ASAP7_75t_R _24467_ (.A1(_06369_),
    .A2(_06370_),
    .B1(_06374_),
    .B2(_06339_),
    .C(_06230_),
    .Y(_06380_));
 INVx1_ASAP7_75t_R _24468_ (.A(_01937_),
    .Y(_06381_));
 INVx1_ASAP7_75t_R _24469_ (.A(_01573_),
    .Y(_06382_));
 AO32x1_ASAP7_75t_R _24470_ (.A1(_06381_),
    .A2(_13531_),
    .A3(_14807_),
    .B1(_06371_),
    .B2(_06382_),
    .Y(_06383_));
 AND3x1_ASAP7_75t_R _24471_ (.A(_06373_),
    .B(_06339_),
    .C(_06383_),
    .Y(_06384_));
 AND2x4_ASAP7_75t_R _24472_ (.A(_05557_),
    .B(_06318_),
    .Y(_06385_));
 AOI21x1_ASAP7_75t_R _24473_ (.A1(_01311_),
    .A2(_06385_),
    .B(_06235_),
    .Y(_06386_));
 OAI22x1_ASAP7_75t_R _24474_ (.A1(_06304_),
    .A2(_05798_),
    .B1(_06386_),
    .B2(_00095_),
    .Y(_06387_));
 AO221x2_ASAP7_75t_R _24475_ (.A1(net3089),
    .A2(_06380_),
    .B1(_06384_),
    .B2(_06372_),
    .C(_06387_),
    .Y(_06388_));
 NOR2x2_ASAP7_75t_R _24476_ (.A(net300),
    .B(_06388_),
    .Y(_06389_));
 AOI21x1_ASAP7_75t_R _24477_ (.A1(_01543_),
    .A2(net301),
    .B(net3090),
    .Y(_18581_));
 NOR2x1_ASAP7_75t_R _24478_ (.A(net429),
    .B(_02195_),
    .Y(_06390_));
 AO21x1_ASAP7_75t_R _24479_ (.A1(net429),
    .A2(_18581_),
    .B(_06390_),
    .Y(net247));
 INVx3_ASAP7_75t_R _24480_ (.A(net2202),
    .Y(_06391_));
 OA22x2_ASAP7_75t_R _24481_ (.A1(_01572_),
    .A2(_06219_),
    .B1(_06221_),
    .B2(_01936_),
    .Y(_06392_));
 OA222x2_ASAP7_75t_R _24482_ (.A1(_06391_),
    .A2(_06304_),
    .B1(_06300_),
    .B2(_06392_),
    .C1(_06386_),
    .C2(_00098_),
    .Y(_06393_));
 NOR2x1_ASAP7_75t_R _24483_ (.A(net3126),
    .B(_06375_),
    .Y(_06394_));
 AO21x2_ASAP7_75t_R _24484_ (.A1(_06375_),
    .A2(_06393_),
    .B(net3127),
    .Y(_06395_));
 OR2x2_ASAP7_75t_R _24485_ (.A(net300),
    .B(_06395_),
    .Y(_06396_));
 OA21x2_ASAP7_75t_R _24486_ (.A1(_01542_),
    .A2(net299),
    .B(_06396_),
    .Y(_06397_));
 AND2x2_ASAP7_75t_R _24487_ (.A(_06354_),
    .B(_02194_),
    .Y(_06398_));
 AOI21x1_ASAP7_75t_R _24488_ (.A1(net429),
    .A2(_06397_),
    .B(_06398_),
    .Y(net248));
 TAPCELL_ASAP7_75t_R TAP_902 ();
 OAI22x1_ASAP7_75t_R _24490_ (.A1(_01571_),
    .A2(_06219_),
    .B1(_06221_),
    .B2(_01935_),
    .Y(_06400_));
 OAI22x1_ASAP7_75t_R _24491_ (.A1(_06304_),
    .A2(_05797_),
    .B1(_06386_),
    .B2(_00101_),
    .Y(_06401_));
 AO21x1_ASAP7_75t_R _24492_ (.A1(_06339_),
    .A2(_06400_),
    .B(_06401_),
    .Y(_06402_));
 AOI211x1_ASAP7_75t_R _24493_ (.A1(net3026),
    .A2(_06380_),
    .B(_06402_),
    .C(_06273_),
    .Y(_06403_));
 AOI21x1_ASAP7_75t_R _24494_ (.A1(_01541_),
    .A2(net301),
    .B(_06403_),
    .Y(_18583_));
 NOR2x1_ASAP7_75t_R _24495_ (.A(net429),
    .B(_02193_),
    .Y(_06404_));
 AO21x1_ASAP7_75t_R _24496_ (.A1(net429),
    .A2(_18583_),
    .B(_06404_),
    .Y(net219));
 TAPCELL_ASAP7_75t_R TAP_901 ();
 NOR2x1_ASAP7_75t_R _24498_ (.A(net2922),
    .B(_06375_),
    .Y(_06406_));
 AND3x1_ASAP7_75t_R _24499_ (.A(net262),
    .B(_14791_),
    .C(_06369_),
    .Y(_06407_));
 AO21x1_ASAP7_75t_R _24500_ (.A1(_06225_),
    .A2(_01715_),
    .B(_06407_),
    .Y(_06408_));
 AO21x2_ASAP7_75t_R _24501_ (.A1(_05557_),
    .A2(_06318_),
    .B(_06235_),
    .Y(_06409_));
 INVx1_ASAP7_75t_R _24502_ (.A(_00657_),
    .Y(_06410_));
 AO21x1_ASAP7_75t_R _24503_ (.A1(_05724_),
    .A2(_06385_),
    .B(_06410_),
    .Y(_06411_));
 AOI22x1_ASAP7_75t_R _24504_ (.A1(_01716_),
    .A2(_06408_),
    .B1(_06409_),
    .B2(_06411_),
    .Y(_06412_));
 OAI22x1_ASAP7_75t_R _24505_ (.A1(_01570_),
    .A2(_06219_),
    .B1(_06221_),
    .B2(_01934_),
    .Y(_06413_));
 NAND2x1_ASAP7_75t_R _24506_ (.A(_06339_),
    .B(_06413_),
    .Y(_06414_));
 AND3x1_ASAP7_75t_R _24507_ (.A(_06375_),
    .B(_06412_),
    .C(_06414_),
    .Y(_06415_));
 OR3x4_ASAP7_75t_R _24508_ (.A(_06273_),
    .B(net2923),
    .C(_06415_),
    .Y(_06416_));
 OA21x2_ASAP7_75t_R _24509_ (.A1(_01540_),
    .A2(net299),
    .B(_06416_),
    .Y(_06417_));
 AND2x2_ASAP7_75t_R _24510_ (.A(_06354_),
    .B(_02192_),
    .Y(_06418_));
 AOI21x1_ASAP7_75t_R _24511_ (.A1(_00237_),
    .A2(_06417_),
    .B(_06418_),
    .Y(net220));
 NAND2x1_ASAP7_75t_R _24512_ (.A(net3161),
    .B(_06380_),
    .Y(_06419_));
 OR2x6_ASAP7_75t_R _24513_ (.A(_05727_),
    .B(_06300_),
    .Y(_06420_));
 TAPCELL_ASAP7_75t_R TAP_900 ();
 OA22x2_ASAP7_75t_R _24515_ (.A1(_06304_),
    .A2(_05796_),
    .B1(_06386_),
    .B2(_00656_),
    .Y(_06422_));
 OA21x2_ASAP7_75t_R _24516_ (.A1(_01569_),
    .A2(_06420_),
    .B(_06422_),
    .Y(_06423_));
 OA211x2_ASAP7_75t_R _24517_ (.A1(_01933_),
    .A2(_06301_),
    .B(net3162),
    .C(_06423_),
    .Y(_06424_));
 AND2x2_ASAP7_75t_R _24518_ (.A(net299),
    .B(_06424_),
    .Y(_06425_));
 AOI21x1_ASAP7_75t_R _24519_ (.A1(_01539_),
    .A2(net301),
    .B(_06425_),
    .Y(_18584_));
 NOR2x1_ASAP7_75t_R _24520_ (.A(net429),
    .B(_02191_),
    .Y(_06426_));
 AO21x1_ASAP7_75t_R _24521_ (.A1(net429),
    .A2(_18584_),
    .B(_06426_),
    .Y(net221));
 INVx1_ASAP7_75t_R _24522_ (.A(_02190_),
    .Y(_06427_));
 INVx3_ASAP7_75t_R _24523_ (.A(net154),
    .Y(_06428_));
 OA22x2_ASAP7_75t_R _24524_ (.A1(_01568_),
    .A2(_06219_),
    .B1(_06221_),
    .B2(_01932_),
    .Y(_06429_));
 OA222x2_ASAP7_75t_R _24525_ (.A1(_06428_),
    .A2(_06304_),
    .B1(_06300_),
    .B2(_06429_),
    .C1(_06386_),
    .C2(_00108_),
    .Y(_06430_));
 NOR2x1_ASAP7_75t_R _24526_ (.A(net3224),
    .B(_06375_),
    .Y(_06431_));
 AO21x2_ASAP7_75t_R _24527_ (.A1(_06375_),
    .A2(_06430_),
    .B(net3225),
    .Y(_06432_));
 NOR2x1_ASAP7_75t_R _24528_ (.A(net300),
    .B(_06432_),
    .Y(_06433_));
 NOR2x1_ASAP7_75t_R _24529_ (.A(_01538_),
    .B(net299),
    .Y(_06434_));
 OR3x1_ASAP7_75t_R _24530_ (.A(_06354_),
    .B(_06433_),
    .C(_06434_),
    .Y(_06435_));
 OA21x2_ASAP7_75t_R _24531_ (.A1(net429),
    .A2(_06427_),
    .B(_06435_),
    .Y(net222));
 NAND2x1_ASAP7_75t_R _24532_ (.A(net3166),
    .B(_06380_),
    .Y(_06436_));
 OA22x2_ASAP7_75t_R _24533_ (.A1(_06304_),
    .A2(_15778_),
    .B1(_06386_),
    .B2(_00111_),
    .Y(_06437_));
 OA21x2_ASAP7_75t_R _24534_ (.A1(_01567_),
    .A2(_06420_),
    .B(_06437_),
    .Y(_06438_));
 OA211x2_ASAP7_75t_R _24535_ (.A1(_01931_),
    .A2(_06301_),
    .B(net3167),
    .C(_06438_),
    .Y(_06439_));
 AND2x2_ASAP7_75t_R _24536_ (.A(net299),
    .B(_06439_),
    .Y(_06440_));
 AOI21x1_ASAP7_75t_R _24537_ (.A1(_01537_),
    .A2(net301),
    .B(net3168),
    .Y(_18586_));
 NOR2x1_ASAP7_75t_R _24538_ (.A(net429),
    .B(_02189_),
    .Y(_06441_));
 AO21x1_ASAP7_75t_R _24539_ (.A1(net429),
    .A2(_18586_),
    .B(_06441_),
    .Y(net223));
 NAND2x1_ASAP7_75t_R _24540_ (.A(net3194),
    .B(_06380_),
    .Y(_06442_));
 OA22x2_ASAP7_75t_R _24541_ (.A1(_00785_),
    .A2(_06304_),
    .B1(_06386_),
    .B2(_00114_),
    .Y(_06443_));
 OA21x2_ASAP7_75t_R _24542_ (.A1(_01566_),
    .A2(_06420_),
    .B(_06443_),
    .Y(_06444_));
 OA211x2_ASAP7_75t_R _24543_ (.A1(_01930_),
    .A2(_06301_),
    .B(net3195),
    .C(_06444_),
    .Y(_06445_));
 AND2x2_ASAP7_75t_R _24544_ (.A(net299),
    .B(_06445_),
    .Y(_06446_));
 AO21x1_ASAP7_75t_R _24545_ (.A1(_01536_),
    .A2(net301),
    .B(_06446_),
    .Y(_06447_));
 AND2x2_ASAP7_75t_R _24546_ (.A(_06354_),
    .B(_02188_),
    .Y(_06448_));
 AOI21x1_ASAP7_75t_R _24547_ (.A1(_00237_),
    .A2(_06447_),
    .B(_06448_),
    .Y(net224));
 INVx1_ASAP7_75t_R _24548_ (.A(net3043),
    .Y(_06449_));
 NOR2x2_ASAP7_75t_R _24549_ (.A(_06230_),
    .B(_06409_),
    .Y(_06450_));
 OA21x2_ASAP7_75t_R _24550_ (.A1(_01311_),
    .A2(_06319_),
    .B(_06231_),
    .Y(_06451_));
 AND2x2_ASAP7_75t_R _24551_ (.A(_00117_),
    .B(_06451_),
    .Y(_06452_));
 OA222x2_ASAP7_75t_R _24552_ (.A1(_06304_),
    .A2(_05795_),
    .B1(_06450_),
    .B2(_06452_),
    .C1(_06301_),
    .C2(_01929_),
    .Y(_06453_));
 OA21x2_ASAP7_75t_R _24553_ (.A1(_01565_),
    .A2(_06308_),
    .B(_06453_),
    .Y(_06454_));
 OA211x2_ASAP7_75t_R _24554_ (.A1(net3044),
    .A2(_06375_),
    .B(_06454_),
    .C(_06296_),
    .Y(_06455_));
 AOI21x1_ASAP7_75t_R _24555_ (.A1(_01535_),
    .A2(net301),
    .B(_06455_),
    .Y(_18588_));
 NOR2x1_ASAP7_75t_R _24556_ (.A(net429),
    .B(_02187_),
    .Y(_06456_));
 AO21x1_ASAP7_75t_R _24557_ (.A1(net429),
    .A2(_18588_),
    .B(_06456_),
    .Y(net225));
 NAND2x1_ASAP7_75t_R _24558_ (.A(net3199),
    .B(_06380_),
    .Y(_06457_));
 NAND2x1_ASAP7_75t_R _24559_ (.A(net259),
    .B(_14796_),
    .Y(_06458_));
 OA21x2_ASAP7_75t_R _24560_ (.A1(_00120_),
    .A2(_06386_),
    .B(_06458_),
    .Y(_06459_));
 OA21x2_ASAP7_75t_R _24561_ (.A1(_01564_),
    .A2(_06420_),
    .B(_06459_),
    .Y(_06460_));
 OA211x2_ASAP7_75t_R _24562_ (.A1(_01928_),
    .A2(_06301_),
    .B(net3200),
    .C(_06460_),
    .Y(_06461_));
 AND2x2_ASAP7_75t_R _24563_ (.A(net299),
    .B(_06461_),
    .Y(_06462_));
 AO21x2_ASAP7_75t_R _24564_ (.A1(_01534_),
    .A2(net301),
    .B(_06462_),
    .Y(_06463_));
 AND2x2_ASAP7_75t_R _24565_ (.A(_06354_),
    .B(_02186_),
    .Y(_06464_));
 AOI21x1_ASAP7_75t_R _24566_ (.A1(net429),
    .A2(_06463_),
    .B(_06464_),
    .Y(net226));
 INVx1_ASAP7_75t_R _24567_ (.A(_01563_),
    .Y(_06465_));
 TAPCELL_ASAP7_75t_R TAP_899 ();
 OAI22x1_ASAP7_75t_R _24569_ (.A1(_06304_),
    .A2(_16263_),
    .B1(_06386_),
    .B2(_00123_),
    .Y(_06467_));
 AOI221x1_ASAP7_75t_R _24570_ (.A1(_06465_),
    .A2(_06366_),
    .B1(_06380_),
    .B2(net3233),
    .C(_06467_),
    .Y(_06468_));
 OA211x2_ASAP7_75t_R _24571_ (.A1(_01927_),
    .A2(_06301_),
    .B(_06468_),
    .C(_06296_),
    .Y(_06469_));
 AOI21x1_ASAP7_75t_R _24572_ (.A1(_01533_),
    .A2(net301),
    .B(_06469_),
    .Y(_18590_));
 NOR2x1_ASAP7_75t_R _24573_ (.A(_00237_),
    .B(_02185_),
    .Y(_06470_));
 AO21x1_ASAP7_75t_R _24574_ (.A1(_00237_),
    .A2(_18590_),
    .B(_06470_),
    .Y(net227));
 NAND2x1_ASAP7_75t_R _24575_ (.A(net3172),
    .B(_06380_),
    .Y(_06471_));
 INVx3_ASAP7_75t_R _24576_ (.A(net160),
    .Y(_06472_));
 OA22x2_ASAP7_75t_R _24577_ (.A1(_06472_),
    .A2(_06304_),
    .B1(_06386_),
    .B2(_00126_),
    .Y(_06473_));
 OA211x2_ASAP7_75t_R _24578_ (.A1(_01562_),
    .A2(_06420_),
    .B(net3173),
    .C(_06473_),
    .Y(_06474_));
 OA211x2_ASAP7_75t_R _24579_ (.A1(_01926_),
    .A2(_06301_),
    .B(_06474_),
    .C(_06296_),
    .Y(_06475_));
 AOI21x1_ASAP7_75t_R _24580_ (.A1(_01532_),
    .A2(net301),
    .B(_06475_),
    .Y(_06476_));
 NOR2x1_ASAP7_75t_R _24581_ (.A(_00237_),
    .B(_02184_),
    .Y(_06477_));
 AO21x1_ASAP7_75t_R _24582_ (.A1(_00237_),
    .A2(_06476_),
    .B(_06477_),
    .Y(net228));
 INVx1_ASAP7_75t_R _24583_ (.A(net3204),
    .Y(_06478_));
 AND2x2_ASAP7_75t_R _24584_ (.A(_00129_),
    .B(_06451_),
    .Y(_06479_));
 OA222x2_ASAP7_75t_R _24585_ (.A1(_06304_),
    .A2(_16509_),
    .B1(_06450_),
    .B2(_06479_),
    .C1(_06301_),
    .C2(_01925_),
    .Y(_06480_));
 OA21x2_ASAP7_75t_R _24586_ (.A1(_01561_),
    .A2(_06308_),
    .B(_06480_),
    .Y(_06481_));
 OA211x2_ASAP7_75t_R _24587_ (.A1(net3205),
    .A2(_06375_),
    .B(_06481_),
    .C(_06296_),
    .Y(_06482_));
 AOI21x1_ASAP7_75t_R _24588_ (.A1(_01531_),
    .A2(net301),
    .B(_06482_),
    .Y(_18592_));
 TAPCELL_ASAP7_75t_R TAP_898 ();
 NOR2x1_ASAP7_75t_R _24590_ (.A(_00237_),
    .B(_02183_),
    .Y(_06484_));
 AO21x1_ASAP7_75t_R _24591_ (.A1(_00237_),
    .A2(_18592_),
    .B(_06484_),
    .Y(net229));
 INVx1_ASAP7_75t_R _24592_ (.A(_01560_),
    .Y(_06485_));
 NOR2x1_ASAP7_75t_R _24593_ (.A(_00132_),
    .B(_06386_),
    .Y(_06486_));
 AO21x1_ASAP7_75t_R _24594_ (.A1(net258),
    .A2(_14796_),
    .B(_06486_),
    .Y(_06487_));
 AOI221x1_ASAP7_75t_R _24595_ (.A1(_06485_),
    .A2(_06366_),
    .B1(_06380_),
    .B2(net3014),
    .C(_06487_),
    .Y(_06488_));
 OA211x2_ASAP7_75t_R _24596_ (.A1(_01924_),
    .A2(_06301_),
    .B(_06488_),
    .C(_06296_),
    .Y(_06489_));
 AOI21x1_ASAP7_75t_R _24597_ (.A1(_01530_),
    .A2(net301),
    .B(_06489_),
    .Y(_06490_));
 NOR2x1_ASAP7_75t_R _24598_ (.A(_00237_),
    .B(_02182_),
    .Y(_06491_));
 AO21x1_ASAP7_75t_R _24599_ (.A1(_00237_),
    .A2(_06490_),
    .B(_06491_),
    .Y(net230));
 INVx1_ASAP7_75t_R _24600_ (.A(_01559_),
    .Y(_06492_));
 OAI22x1_ASAP7_75t_R _24601_ (.A1(_06304_),
    .A2(_04517_),
    .B1(_06386_),
    .B2(_00135_),
    .Y(_06493_));
 AOI221x1_ASAP7_75t_R _24602_ (.A1(_06492_),
    .A2(_06366_),
    .B1(_06380_),
    .B2(net3220),
    .C(_06493_),
    .Y(_06494_));
 OA211x2_ASAP7_75t_R _24603_ (.A1(_01923_),
    .A2(_06301_),
    .B(_06494_),
    .C(_06296_),
    .Y(_06495_));
 AOI21x1_ASAP7_75t_R _24604_ (.A1(_01529_),
    .A2(net301),
    .B(_06495_),
    .Y(_18594_));
 NOR2x1_ASAP7_75t_R _24605_ (.A(net429),
    .B(_02181_),
    .Y(_06496_));
 AO21x1_ASAP7_75t_R _24606_ (.A1(net429),
    .A2(_18594_),
    .B(_06496_),
    .Y(net231));
 NAND2x1_ASAP7_75t_R _24607_ (.A(net3215),
    .B(_06380_),
    .Y(_06497_));
 INVx4_ASAP7_75t_R _24608_ (.A(net2177),
    .Y(_06498_));
 OA22x2_ASAP7_75t_R _24609_ (.A1(_06498_),
    .A2(_06304_),
    .B1(_06386_),
    .B2(_00138_),
    .Y(_06499_));
 OA21x2_ASAP7_75t_R _24610_ (.A1(_01558_),
    .A2(_06420_),
    .B(_06499_),
    .Y(_06500_));
 OA211x2_ASAP7_75t_R _24611_ (.A1(_01922_),
    .A2(_06301_),
    .B(net3216),
    .C(_06500_),
    .Y(_06501_));
 AND2x2_ASAP7_75t_R _24612_ (.A(net299),
    .B(_06501_),
    .Y(_06502_));
 AOI21x1_ASAP7_75t_R _24613_ (.A1(_01528_),
    .A2(net301),
    .B(_06502_),
    .Y(_06503_));
 NOR2x1_ASAP7_75t_R _24614_ (.A(_00237_),
    .B(_02180_),
    .Y(_06504_));
 AO21x1_ASAP7_75t_R _24615_ (.A1(_00237_),
    .A2(_06503_),
    .B(_06504_),
    .Y(net232));
 NAND2x1_ASAP7_75t_R _24616_ (.A(net3177),
    .B(_06380_),
    .Y(_06505_));
 OA22x2_ASAP7_75t_R _24617_ (.A1(_06304_),
    .A2(_04747_),
    .B1(_06386_),
    .B2(_00141_),
    .Y(_06506_));
 OA211x2_ASAP7_75t_R _24618_ (.A1(_01557_),
    .A2(_06420_),
    .B(net3178),
    .C(_06506_),
    .Y(_06507_));
 OA211x2_ASAP7_75t_R _24619_ (.A1(_01921_),
    .A2(_06301_),
    .B(_06507_),
    .C(_06296_),
    .Y(_06508_));
 AOI21x1_ASAP7_75t_R _24620_ (.A1(_01527_),
    .A2(net301),
    .B(_06508_),
    .Y(_18596_));
 NOR2x1_ASAP7_75t_R _24621_ (.A(_00237_),
    .B(_02179_),
    .Y(_06509_));
 AO21x1_ASAP7_75t_R _24622_ (.A1(_00237_),
    .A2(_18596_),
    .B(_06509_),
    .Y(net233));
 INVx1_ASAP7_75t_R _24623_ (.A(net3156),
    .Y(_06510_));
 INVx3_ASAP7_75t_R _24624_ (.A(net2175),
    .Y(_06511_));
 AO21x1_ASAP7_75t_R _24625_ (.A1(_00144_),
    .A2(_06451_),
    .B(_06450_),
    .Y(_06512_));
 OA21x2_ASAP7_75t_R _24626_ (.A1(_06511_),
    .A2(_06304_),
    .B(_06512_),
    .Y(_06513_));
 OA22x2_ASAP7_75t_R _24627_ (.A1(_01920_),
    .A2(_06301_),
    .B1(_06308_),
    .B2(_01556_),
    .Y(_06514_));
 OA211x2_ASAP7_75t_R _24628_ (.A1(net3157),
    .A2(_06375_),
    .B(_06513_),
    .C(_06514_),
    .Y(_06515_));
 AND2x2_ASAP7_75t_R _24629_ (.A(_01526_),
    .B(net301),
    .Y(_06516_));
 AOI21x1_ASAP7_75t_R _24630_ (.A1(net299),
    .A2(_06515_),
    .B(_06516_),
    .Y(_06517_));
 NOR2x1_ASAP7_75t_R _24631_ (.A(_00237_),
    .B(_02178_),
    .Y(_06518_));
 AO21x1_ASAP7_75t_R _24632_ (.A1(_00237_),
    .A2(_06517_),
    .B(_06518_),
    .Y(net234));
 TAPCELL_ASAP7_75t_R TAP_897 ();
 INVx1_ASAP7_75t_R _24634_ (.A(_01555_),
    .Y(_06520_));
 OAI22x1_ASAP7_75t_R _24635_ (.A1(_06304_),
    .A2(_04968_),
    .B1(_06386_),
    .B2(_00147_),
    .Y(_06521_));
 AOI221x1_ASAP7_75t_R _24636_ (.A1(_06520_),
    .A2(_06366_),
    .B1(_06380_),
    .B2(net3237),
    .C(_06521_),
    .Y(_06522_));
 OA211x2_ASAP7_75t_R _24637_ (.A1(_01919_),
    .A2(_06301_),
    .B(_06522_),
    .C(_06296_),
    .Y(_06523_));
 AOI21x1_ASAP7_75t_R _24638_ (.A1(_01525_),
    .A2(net301),
    .B(_06523_),
    .Y(_18598_));
 NOR2x1_ASAP7_75t_R _24639_ (.A(_00237_),
    .B(_02177_),
    .Y(_06524_));
 AO21x1_ASAP7_75t_R _24640_ (.A1(_00237_),
    .A2(_18598_),
    .B(_06524_),
    .Y(net235));
 INVx1_ASAP7_75t_R _24641_ (.A(net3146),
    .Y(_06525_));
 INVx4_ASAP7_75t_R _24642_ (.A(net2155),
    .Y(_06526_));
 AO21x1_ASAP7_75t_R _24643_ (.A1(_00150_),
    .A2(_06451_),
    .B(_06450_),
    .Y(_06527_));
 OA21x2_ASAP7_75t_R _24644_ (.A1(_06526_),
    .A2(_06304_),
    .B(_06527_),
    .Y(_06528_));
 OA22x2_ASAP7_75t_R _24645_ (.A1(_01918_),
    .A2(_06301_),
    .B1(_06308_),
    .B2(_01554_),
    .Y(_06529_));
 OA211x2_ASAP7_75t_R _24646_ (.A1(net3147),
    .A2(_06375_),
    .B(_06528_),
    .C(_06529_),
    .Y(_06530_));
 AND2x2_ASAP7_75t_R _24647_ (.A(_01524_),
    .B(net301),
    .Y(_06531_));
 AOI21x1_ASAP7_75t_R _24648_ (.A1(net299),
    .A2(_06530_),
    .B(_06531_),
    .Y(_06532_));
 NOR2x1_ASAP7_75t_R _24649_ (.A(net429),
    .B(_02176_),
    .Y(_06533_));
 AO21x1_ASAP7_75t_R _24650_ (.A1(net429),
    .A2(_06532_),
    .B(_06533_),
    .Y(net236));
 INVx1_ASAP7_75t_R _24651_ (.A(net3151),
    .Y(_06534_));
 AND2x2_ASAP7_75t_R _24652_ (.A(_00153_),
    .B(_06451_),
    .Y(_06535_));
 OA222x2_ASAP7_75t_R _24653_ (.A1(_06304_),
    .A2(_05185_),
    .B1(_06450_),
    .B2(_06535_),
    .C1(_06301_),
    .C2(_01917_),
    .Y(_06536_));
 OA21x2_ASAP7_75t_R _24654_ (.A1(_01553_),
    .A2(_06308_),
    .B(_06536_),
    .Y(_06537_));
 OA211x2_ASAP7_75t_R _24655_ (.A1(net3152),
    .A2(_06375_),
    .B(_06537_),
    .C(_06296_),
    .Y(_06538_));
 AOI21x1_ASAP7_75t_R _24656_ (.A1(_01523_),
    .A2(net301),
    .B(_06538_),
    .Y(_18600_));
 NOR2x1_ASAP7_75t_R _24657_ (.A(_00237_),
    .B(_02175_),
    .Y(_06539_));
 AO21x1_ASAP7_75t_R _24658_ (.A1(_00237_),
    .A2(_18600_),
    .B(_06539_),
    .Y(net237));
 NAND2x1_ASAP7_75t_R _24659_ (.A(net3189),
    .B(_06380_),
    .Y(_06540_));
 INVx2_ASAP7_75t_R _24660_ (.A(net2141),
    .Y(_06541_));
 OA22x2_ASAP7_75t_R _24661_ (.A1(_06541_),
    .A2(_06304_),
    .B1(_06386_),
    .B2(_00156_),
    .Y(_06542_));
 OA211x2_ASAP7_75t_R _24662_ (.A1(_01552_),
    .A2(_06420_),
    .B(net3190),
    .C(_06542_),
    .Y(_06543_));
 OA211x2_ASAP7_75t_R _24663_ (.A1(_01916_),
    .A2(_06301_),
    .B(_06543_),
    .C(_06296_),
    .Y(_06544_));
 AOI21x1_ASAP7_75t_R _24664_ (.A1(_01522_),
    .A2(net301),
    .B(_06544_),
    .Y(_06545_));
 NOR2x1_ASAP7_75t_R _24665_ (.A(_00237_),
    .B(_02174_),
    .Y(_06546_));
 AO21x1_ASAP7_75t_R _24666_ (.A1(_00237_),
    .A2(_06545_),
    .B(_06546_),
    .Y(net238));
 INVx1_ASAP7_75t_R _24667_ (.A(_01551_),
    .Y(_06547_));
 OAI22x1_ASAP7_75t_R _24668_ (.A1(_06304_),
    .A2(_05404_),
    .B1(_06386_),
    .B2(_00159_),
    .Y(_06548_));
 AOI221x1_ASAP7_75t_R _24669_ (.A1(_06547_),
    .A2(_06366_),
    .B1(_06380_),
    .B2(net3229),
    .C(_06548_),
    .Y(_06549_));
 OA211x2_ASAP7_75t_R _24670_ (.A1(_01915_),
    .A2(_06301_),
    .B(_06549_),
    .C(_06296_),
    .Y(_06550_));
 AOI21x1_ASAP7_75t_R _24671_ (.A1(_01521_),
    .A2(net301),
    .B(_06550_),
    .Y(_18602_));
 NOR2x1_ASAP7_75t_R _24672_ (.A(_00237_),
    .B(_02173_),
    .Y(_06551_));
 AO21x1_ASAP7_75t_R _24673_ (.A1(_00237_),
    .A2(_18602_),
    .B(_06551_),
    .Y(net240));
 INVx1_ASAP7_75t_R _24674_ (.A(net3063),
    .Y(_06552_));
 OR3x1_ASAP7_75t_R _24675_ (.A(_06304_),
    .B(_05540_),
    .C(_05541_),
    .Y(_06553_));
 OA22x2_ASAP7_75t_R _24676_ (.A1(_01914_),
    .A2(_06301_),
    .B1(_06308_),
    .B2(_01550_),
    .Y(_06554_));
 OA211x2_ASAP7_75t_R _24677_ (.A1(_00161_),
    .A2(_06386_),
    .B(_06554_),
    .C(_06375_),
    .Y(_06555_));
 AO221x2_ASAP7_75t_R _24678_ (.A1(net3064),
    .A2(_06380_),
    .B1(_06553_),
    .B2(_06555_),
    .C(_06273_),
    .Y(_06556_));
 OAI21x1_ASAP7_75t_R _24679_ (.A1(_01520_),
    .A2(net299),
    .B(net3065),
    .Y(_06557_));
 NAND2x1_ASAP7_75t_R _24680_ (.A(_06354_),
    .B(_01729_),
    .Y(_06558_));
 OA21x2_ASAP7_75t_R _24681_ (.A1(_06354_),
    .A2(_06557_),
    .B(_06558_),
    .Y(net241));
 TAPCELL_ASAP7_75t_R TAP_896 ();
 TAPCELL_ASAP7_75t_R TAP_895 ();
 AO21x1_ASAP7_75t_R _24684_ (.A1(_01815_),
    .A2(_01736_),
    .B(_00239_),
    .Y(_06561_));
 AND2x2_ASAP7_75t_R _24685_ (.A(_01714_),
    .B(_01717_),
    .Y(_06562_));
 NOR2x1_ASAP7_75t_R _24686_ (.A(_06227_),
    .B(_06562_),
    .Y(_06563_));
 OA21x2_ASAP7_75t_R _24687_ (.A1(_06369_),
    .A2(_06563_),
    .B(_00238_),
    .Y(_06564_));
 OAI21x1_ASAP7_75t_R _24688_ (.A1(net299),
    .A2(_06561_),
    .B(_06564_),
    .Y(_06565_));
 NAND2x2_ASAP7_75t_R _24689_ (.A(_00237_),
    .B(_06565_),
    .Y(net249));
 AOI21x1_ASAP7_75t_R _24690_ (.A1(_00238_),
    .A2(net2739),
    .B(_01736_),
    .Y(_06566_));
 AO21x1_ASAP7_75t_R _24691_ (.A1(net2758),
    .A2(net249),
    .B(_06566_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 INVx1_ASAP7_75t_R _24692_ (.A(net2758),
    .Y(_06567_));
 INVx1_ASAP7_75t_R _24693_ (.A(net249),
    .Y(_06568_));
 OR3x1_ASAP7_75t_R _24694_ (.A(net2759),
    .B(_01736_),
    .C(_06568_),
    .Y(_06569_));
 INVx2_ASAP7_75t_R _24695_ (.A(_01736_),
    .Y(_06570_));
 AND2x4_ASAP7_75t_R _24696_ (.A(net2739),
    .B(_06570_),
    .Y(_06571_));
 AOI21x1_ASAP7_75t_R _24697_ (.A1(_00238_),
    .A2(_06569_),
    .B(net2741),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 AO21x1_ASAP7_75t_R _24698_ (.A1(_01735_),
    .A2(net300),
    .B(net429),
    .Y(_06572_));
 INVx1_ASAP7_75t_R _24699_ (.A(_06572_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 TAPCELL_ASAP7_75t_R TAP_894 ();
 OR3x1_ASAP7_75t_R _24701_ (.A(net2759),
    .B(_01736_),
    .C(_06572_),
    .Y(_06574_));
 OA211x2_ASAP7_75t_R _24702_ (.A1(_00238_),
    .A2(net300),
    .B(_06574_),
    .C(_01848_),
    .Y(_06575_));
 OAI21x1_ASAP7_75t_R _24703_ (.A1(net2739),
    .A2(net299),
    .B(_06570_),
    .Y(_06576_));
 OA211x2_ASAP7_75t_R _24704_ (.A1(net2759),
    .A2(_06572_),
    .B(_06576_),
    .C(_01737_),
    .Y(_06577_));
 AO21x1_ASAP7_75t_R _24705_ (.A1(net2741),
    .A2(_06575_),
    .B(net2976),
    .Y(_06578_));
 INVx1_ASAP7_75t_R _24706_ (.A(net2977),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 NOR2x1_ASAP7_75t_R _24707_ (.A(net2741),
    .B(_06575_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 TAPCELL_ASAP7_75t_R TAP_893 ();
 CKINVDCx16_ASAP7_75t_R _24709_ (.A(net430),
    .Y(_06580_));
 TAPCELL_ASAP7_75t_R TAP_892 ();
 TAPCELL_ASAP7_75t_R TAP_891 ();
 TAPCELL_ASAP7_75t_R TAP_890 ();
 INVx1_ASAP7_75t_R _24713_ (.A(net2692),
    .Y(_06584_));
 TAPCELL_ASAP7_75t_R TAP_889 ();
 NAND2x1_ASAP7_75t_R _24715_ (.A(_00240_),
    .B(net2625),
    .Y(_06586_));
 OR3x1_ASAP7_75t_R _24716_ (.A(_00240_),
    .B(_01829_),
    .C(_01830_),
    .Y(_06587_));
 OA21x2_ASAP7_75t_R _24717_ (.A1(_06584_),
    .A2(_06586_),
    .B(_06587_),
    .Y(_06588_));
 CKINVDCx20_ASAP7_75t_R _24718_ (.A(net428),
    .Y(_06589_));
 TAPCELL_ASAP7_75t_R TAP_888 ();
 INVx2_ASAP7_75t_R _24720_ (.A(net2935),
    .Y(_06591_));
 AND2x2_ASAP7_75t_R _24721_ (.A(_00240_),
    .B(net2936),
    .Y(_06592_));
 AO21x1_ASAP7_75t_R _24722_ (.A1(_06589_),
    .A2(_01814_),
    .B(_06592_),
    .Y(_06593_));
 AND3x2_ASAP7_75t_R _24723_ (.A(_06580_),
    .B(_06588_),
    .C(_06593_),
    .Y(_17752_));
 OR3x1_ASAP7_75t_R _24724_ (.A(_00242_),
    .B(_01605_),
    .C(_01606_),
    .Y(_06594_));
 INVx1_ASAP7_75t_R _24725_ (.A(_06594_),
    .Y(_18561_));
 OR5x1_ASAP7_75t_R _24726_ (.A(_00242_),
    .B(_01603_),
    .C(_01604_),
    .D(_01605_),
    .E(_01606_),
    .Y(_06595_));
 INVx1_ASAP7_75t_R _24727_ (.A(_06595_),
    .Y(_18562_));
 OR3x1_ASAP7_75t_R _24728_ (.A(_01601_),
    .B(_01602_),
    .C(_06595_),
    .Y(_06596_));
 INVx1_ASAP7_75t_R _24729_ (.A(_06596_),
    .Y(_18563_));
 OR3x1_ASAP7_75t_R _24730_ (.A(_01599_),
    .B(_01600_),
    .C(_06596_),
    .Y(_06597_));
 INVx1_ASAP7_75t_R _24731_ (.A(_06597_),
    .Y(_18564_));
 OR3x1_ASAP7_75t_R _24732_ (.A(_01597_),
    .B(_01598_),
    .C(_06597_),
    .Y(_06598_));
 INVx1_ASAP7_75t_R _24733_ (.A(_06598_),
    .Y(_18565_));
 OR3x1_ASAP7_75t_R _24734_ (.A(_01595_),
    .B(_01596_),
    .C(_06598_),
    .Y(_06599_));
 INVx1_ASAP7_75t_R _24735_ (.A(_06599_),
    .Y(_18566_));
 OR3x1_ASAP7_75t_R _24736_ (.A(_01593_),
    .B(_01594_),
    .C(_06599_),
    .Y(_06600_));
 INVx1_ASAP7_75t_R _24737_ (.A(_06600_),
    .Y(_18567_));
 OR3x1_ASAP7_75t_R _24738_ (.A(_01591_),
    .B(_01592_),
    .C(_06600_),
    .Y(_06601_));
 INVx1_ASAP7_75t_R _24739_ (.A(_06601_),
    .Y(_18568_));
 OR3x1_ASAP7_75t_R _24740_ (.A(_01589_),
    .B(_01590_),
    .C(_06601_),
    .Y(_06602_));
 INVx1_ASAP7_75t_R _24741_ (.A(_06602_),
    .Y(_18569_));
 OR3x1_ASAP7_75t_R _24742_ (.A(_01587_),
    .B(_01588_),
    .C(_06602_),
    .Y(_06603_));
 INVx1_ASAP7_75t_R _24743_ (.A(_06603_),
    .Y(_18570_));
 OR3x1_ASAP7_75t_R _24744_ (.A(_01585_),
    .B(_01586_),
    .C(_06603_),
    .Y(_06604_));
 INVx1_ASAP7_75t_R _24745_ (.A(_06604_),
    .Y(_18571_));
 OR3x1_ASAP7_75t_R _24746_ (.A(_01583_),
    .B(_01584_),
    .C(_06604_),
    .Y(_06605_));
 INVx1_ASAP7_75t_R _24747_ (.A(_06605_),
    .Y(_18572_));
 OR3x1_ASAP7_75t_R _24748_ (.A(_01581_),
    .B(_01582_),
    .C(_06605_),
    .Y(_06606_));
 INVx1_ASAP7_75t_R _24749_ (.A(_06606_),
    .Y(_18573_));
 NOR3x2_ASAP7_75t_R _24750_ (.B(net3356),
    .C(net3209),
    .Y(_06607_),
    .A(net3301));
 AND2x2_ASAP7_75t_R _24751_ (.A(_06228_),
    .B(_01734_),
    .Y(_06608_));
 AO21x1_ASAP7_75t_R _24752_ (.A1(net3302),
    .A2(_06608_),
    .B(_01747_),
    .Y(net150));
 OR3x2_ASAP7_75t_R _24753_ (.A(_14808_),
    .B(_14804_),
    .C(_05725_),
    .Y(_06609_));
 INVx1_ASAP7_75t_R _24754_ (.A(_06374_),
    .Y(_06610_));
 INVx1_ASAP7_75t_R _24755_ (.A(_02287_),
    .Y(_06611_));
 AND2x2_ASAP7_75t_R _24756_ (.A(net2361),
    .B(net333),
    .Y(_06612_));
 AND5x1_ASAP7_75t_R _24757_ (.A(_02288_),
    .B(_06611_),
    .C(_06612_),
    .D(_05571_),
    .E(_06371_),
    .Y(_06613_));
 AND5x1_ASAP7_75t_R _24758_ (.A(net333),
    .B(_02287_),
    .C(_13390_),
    .D(_14813_),
    .E(_05571_),
    .Y(_06614_));
 OAI21x1_ASAP7_75t_R _24759_ (.A1(_06613_),
    .A2(_06614_),
    .B(_05737_),
    .Y(_06615_));
 AND4x2_ASAP7_75t_R _24760_ (.A(net3038),
    .B(_06609_),
    .C(_06610_),
    .D(_06615_),
    .Y(_06616_));
 AND3x1_ASAP7_75t_R _24761_ (.A(_05741_),
    .B(_05747_),
    .C(_06616_),
    .Y(_06617_));
 AO21x2_ASAP7_75t_R _24762_ (.A1(_05723_),
    .A2(_06617_),
    .B(_06304_),
    .Y(_06618_));
 TAPCELL_ASAP7_75t_R TAP_887 ();
 TAPCELL_ASAP7_75t_R TAP_886 ();
 AND4x2_ASAP7_75t_R _24765_ (.A(_01314_),
    .B(_01728_),
    .C(_13817_),
    .D(_05816_),
    .Y(_06621_));
 OA211x2_ASAP7_75t_R _24766_ (.A1(_01713_),
    .A2(_05553_),
    .B(_14828_),
    .C(_13459_),
    .Y(_06622_));
 AO21x1_ASAP7_75t_R _24767_ (.A1(_14797_),
    .A2(_06621_),
    .B(_06622_),
    .Y(_06623_));
 AO21x1_ASAP7_75t_R _24768_ (.A1(_14842_),
    .A2(_06623_),
    .B(_06202_),
    .Y(_06624_));
 AND5x1_ASAP7_75t_R _24769_ (.A(_15778_),
    .B(_16263_),
    .C(_04968_),
    .D(_05185_),
    .E(_05799_),
    .Y(_06625_));
 AND5x1_ASAP7_75t_R _24770_ (.A(_16509_),
    .B(_04517_),
    .C(_04747_),
    .D(_05794_),
    .E(_06625_),
    .Y(_06626_));
 OA21x2_ASAP7_75t_R _24771_ (.A1(_05540_),
    .A2(_05541_),
    .B(_06626_),
    .Y(_06627_));
 AND2x2_ASAP7_75t_R _24772_ (.A(_13588_),
    .B(_13614_),
    .Y(_06628_));
 AND3x2_ASAP7_75t_R _24773_ (.A(_13617_),
    .B(_13548_),
    .C(_13553_),
    .Y(_06629_));
 AND3x2_ASAP7_75t_R _24774_ (.A(_13613_),
    .B(_13594_),
    .C(_06629_),
    .Y(_06630_));
 OR3x1_ASAP7_75t_R _24775_ (.A(_13577_),
    .B(_13606_),
    .C(_06630_),
    .Y(_06631_));
 AO21x1_ASAP7_75t_R _24776_ (.A1(_13578_),
    .A2(_13582_),
    .B(_13583_),
    .Y(_06632_));
 AND2x2_ASAP7_75t_R _24777_ (.A(_13554_),
    .B(_13576_),
    .Y(_06633_));
 AOI211x1_ASAP7_75t_R _24778_ (.A1(_13599_),
    .A2(_13601_),
    .B(_13603_),
    .C(_13605_),
    .Y(_06634_));
 NAND3x2_ASAP7_75t_R _24779_ (.B(_13594_),
    .C(_06629_),
    .Y(_06635_),
    .A(_13613_));
 OR4x1_ASAP7_75t_R _24780_ (.A(_06632_),
    .B(_06633_),
    .C(_06634_),
    .D(_06635_),
    .Y(_06636_));
 AND3x1_ASAP7_75t_R _24781_ (.A(_06628_),
    .B(_06631_),
    .C(_06636_),
    .Y(_06637_));
 NOR2x2_ASAP7_75t_R _24782_ (.A(_13618_),
    .B(_06637_),
    .Y(_06638_));
 AOI21x1_ASAP7_75t_R _24783_ (.A1(_13483_),
    .A2(_06628_),
    .B(_06638_),
    .Y(_06639_));
 AND4x1_ASAP7_75t_R _24784_ (.A(_13476_),
    .B(_13587_),
    .C(_06627_),
    .D(_06639_),
    .Y(_06640_));
 INVx2_ASAP7_75t_R _24785_ (.A(_01310_),
    .Y(_06641_));
 AND2x2_ASAP7_75t_R _24786_ (.A(_06633_),
    .B(_06635_),
    .Y(_06642_));
 AOI22x1_ASAP7_75t_R _24787_ (.A1(_13605_),
    .A2(_06630_),
    .B1(_06642_),
    .B2(_13606_),
    .Y(_06643_));
 XNOR2x1_ASAP7_75t_R _24788_ (.B(_06643_),
    .Y(_06644_),
    .A(_17807_));
 NAND2x1_ASAP7_75t_R _24789_ (.A(_06641_),
    .B(_06644_),
    .Y(_06645_));
 AND3x1_ASAP7_75t_R _24790_ (.A(_13476_),
    .B(_13587_),
    .C(_06638_),
    .Y(_06646_));
 OA211x2_ASAP7_75t_R _24791_ (.A1(_06641_),
    .A2(net173),
    .B(_06645_),
    .C(_06646_),
    .Y(_06647_));
 OR3x1_ASAP7_75t_R _24792_ (.A(_06624_),
    .B(_06640_),
    .C(_06647_),
    .Y(_06648_));
 OAI21x1_ASAP7_75t_R _24793_ (.A1(_06641_),
    .A2(net173),
    .B(_06645_),
    .Y(_06649_));
 AO32x2_ASAP7_75t_R _24794_ (.A1(_13588_),
    .A2(_13562_),
    .A3(_06649_),
    .B1(_05802_),
    .B2(_13583_),
    .Y(_06650_));
 INVx1_ASAP7_75t_R _24795_ (.A(_14828_),
    .Y(_06651_));
 AO21x1_ASAP7_75t_R _24796_ (.A1(_01713_),
    .A2(_06651_),
    .B(_06621_),
    .Y(_06652_));
 AO21x1_ASAP7_75t_R _24797_ (.A1(_14797_),
    .A2(_06652_),
    .B(_06622_),
    .Y(_06653_));
 AND2x2_ASAP7_75t_R _24798_ (.A(_14842_),
    .B(_06653_),
    .Y(_06654_));
 OAI21x1_ASAP7_75t_R _24799_ (.A1(_06648_),
    .A2(_06650_),
    .B(_06654_),
    .Y(_06655_));
 NAND2x1_ASAP7_75t_R _24800_ (.A(_06618_),
    .B(_06655_),
    .Y(_06656_));
 OR3x1_ASAP7_75t_R _24801_ (.A(_06225_),
    .B(_14793_),
    .C(_01716_),
    .Y(_06657_));
 AND3x1_ASAP7_75t_R _24802_ (.A(_13459_),
    .B(_06232_),
    .C(_06657_),
    .Y(_06658_));
 INVx1_ASAP7_75t_R _24803_ (.A(_05801_),
    .Y(_06659_));
 OR3x1_ASAP7_75t_R _24804_ (.A(_13460_),
    .B(_13470_),
    .C(_13463_),
    .Y(_06660_));
 AO21x1_ASAP7_75t_R _24805_ (.A1(_13483_),
    .A2(_06628_),
    .B(_06660_),
    .Y(_06661_));
 OR3x1_ASAP7_75t_R _24806_ (.A(_06659_),
    .B(_06638_),
    .C(_06661_),
    .Y(_06662_));
 INVx1_ASAP7_75t_R _24807_ (.A(_06662_),
    .Y(_06663_));
 AND3x2_ASAP7_75t_R _24808_ (.A(_01714_),
    .B(_01715_),
    .C(_05556_),
    .Y(_06664_));
 OR3x1_ASAP7_75t_R _24809_ (.A(_05557_),
    .B(_06624_),
    .C(_06664_),
    .Y(_06665_));
 AO211x2_ASAP7_75t_R _24810_ (.A1(_05542_),
    .A2(_06663_),
    .B(_06647_),
    .C(_06665_),
    .Y(_06666_));
 OR3x1_ASAP7_75t_R _24811_ (.A(_05557_),
    .B(_06654_),
    .C(_06664_),
    .Y(_06667_));
 OAI21x1_ASAP7_75t_R _24812_ (.A1(_06650_),
    .A2(_06666_),
    .B(_06667_),
    .Y(_06668_));
 INVx1_ASAP7_75t_R _24813_ (.A(_02034_),
    .Y(_06669_));
 AO21x1_ASAP7_75t_R _24814_ (.A1(_13459_),
    .A2(_06669_),
    .B(net3102),
    .Y(_06670_));
 AND2x4_ASAP7_75t_R _24815_ (.A(_01311_),
    .B(net3103),
    .Y(_06671_));
 AO21x2_ASAP7_75t_R _24816_ (.A1(net3132),
    .A2(net3210),
    .B(net3104),
    .Y(_06672_));
 TAPCELL_ASAP7_75t_R TAP_885 ();
 TAPCELL_ASAP7_75t_R TAP_884 ();
 TAPCELL_ASAP7_75t_R TAP_883 ();
 AND2x2_ASAP7_75t_R _24820_ (.A(_06588_),
    .B(_06593_),
    .Y(_06676_));
 NOR2x1_ASAP7_75t_R _24821_ (.A(_00662_),
    .B(_06676_),
    .Y(_06677_));
 NAND2x2_ASAP7_75t_R _24822_ (.A(_01737_),
    .B(net2741),
    .Y(_06678_));
 OR3x1_ASAP7_75t_R _24823_ (.A(_00662_),
    .B(_00239_),
    .C(_06676_),
    .Y(_06679_));
 TAPCELL_ASAP7_75t_R TAP_882 ();
 TAPCELL_ASAP7_75t_R TAP_881 ();
 OA211x2_ASAP7_75t_R _24826_ (.A1(_06677_),
    .A2(_06678_),
    .B(_06679_),
    .C(_00240_),
    .Y(_06682_));
 AND3x1_ASAP7_75t_R _24827_ (.A(_00239_),
    .B(_06677_),
    .C(_06678_),
    .Y(_06683_));
 AOI211x1_ASAP7_75t_R _24828_ (.A1(_14794_),
    .A2(net3105),
    .B(_06682_),
    .C(_06683_),
    .Y(_06684_));
 AND2x6_ASAP7_75t_R _24829_ (.A(_06668_),
    .B(_06684_),
    .Y(_06685_));
 AND2x6_ASAP7_75t_R _24830_ (.A(_06618_),
    .B(_06685_),
    .Y(_06686_));
 TAPCELL_ASAP7_75t_R TAP_880 ();
 TAPCELL_ASAP7_75t_R TAP_879 ();
 AO32x1_ASAP7_75t_R _24833_ (.A1(_06218_),
    .A2(_06656_),
    .A3(_06658_),
    .B1(_06686_),
    .B2(_06273_),
    .Y(\if_stage_i.instr_valid_id_d ));
 AND2x2_ASAP7_75t_R _24834_ (.A(_06627_),
    .B(_06639_),
    .Y(_06689_));
 OA211x2_ASAP7_75t_R _24835_ (.A1(_06641_),
    .A2(net173),
    .B(_06638_),
    .C(_06645_),
    .Y(_06690_));
 NOR3x2_ASAP7_75t_R _24836_ (.B(_06690_),
    .C(_06650_),
    .Y(_06691_),
    .A(_06689_));
 NOR2x1_ASAP7_75t_R _24837_ (.A(_06660_),
    .B(_06691_),
    .Y(_06692_));
 AND4x1_ASAP7_75t_R _24838_ (.A(_01713_),
    .B(_06651_),
    .C(_05752_),
    .D(_06692_),
    .Y(\id_stage_i.branch_set_d ));
 INVx1_ASAP7_75t_R _24839_ (.A(_02566_),
    .Y(_18576_));
 AOI211x1_ASAP7_75t_R _24840_ (.A1(_01546_),
    .A2(net300),
    .B(_06352_),
    .C(_02566_),
    .Y(_06693_));
 AND2x2_ASAP7_75t_R _24841_ (.A(_18577_),
    .B(_06693_),
    .Y(_18578_));
 OR3x1_ASAP7_75t_R _24842_ (.A(_06342_),
    .B(_06361_),
    .C(_06376_),
    .Y(_06694_));
 NOR2x1_ASAP7_75t_R _24843_ (.A(net300),
    .B(_06694_),
    .Y(_06695_));
 OR3x1_ASAP7_75t_R _24844_ (.A(_01544_),
    .B(_01545_),
    .C(_01547_),
    .Y(_06696_));
 NOR2x1_ASAP7_75t_R _24845_ (.A(net299),
    .B(_06696_),
    .Y(_06697_));
 OA21x2_ASAP7_75t_R _24846_ (.A1(_06695_),
    .A2(_06697_),
    .B(_06693_),
    .Y(_18580_));
 NOR3x1_ASAP7_75t_R _24847_ (.A(_01542_),
    .B(_01543_),
    .C(net299),
    .Y(_06698_));
 INVx1_ASAP7_75t_R _24848_ (.A(_06395_),
    .Y(_06699_));
 AND3x1_ASAP7_75t_R _24849_ (.A(net299),
    .B(_06388_),
    .C(_06699_),
    .Y(_06700_));
 OA221x2_ASAP7_75t_R _24850_ (.A1(_06695_),
    .A2(_06697_),
    .B1(_06698_),
    .B2(_06700_),
    .C(_06693_),
    .Y(_18582_));
 NOR2x1_ASAP7_75t_R _24851_ (.A(_01540_),
    .B(_01541_),
    .Y(_06701_));
 NAND2x1_ASAP7_75t_R _24852_ (.A(_06412_),
    .B(_06414_),
    .Y(_06702_));
 AO32x2_ASAP7_75t_R _24853_ (.A1(net3026),
    .A2(net2922),
    .A3(_06380_),
    .B1(_06402_),
    .B2(_06702_),
    .Y(_06703_));
 AND2x2_ASAP7_75t_R _24854_ (.A(net299),
    .B(_06703_),
    .Y(_06704_));
 AO21x1_ASAP7_75t_R _24855_ (.A1(net301),
    .A2(_06701_),
    .B(_06704_),
    .Y(_06705_));
 AND2x2_ASAP7_75t_R _24856_ (.A(_18582_),
    .B(_06705_),
    .Y(_18585_));
 OR3x1_ASAP7_75t_R _24857_ (.A(_01538_),
    .B(_01539_),
    .C(net299),
    .Y(_06706_));
 OR3x1_ASAP7_75t_R _24858_ (.A(net301),
    .B(_06424_),
    .C(_06432_),
    .Y(_06707_));
 NAND2x1_ASAP7_75t_R _24859_ (.A(_06706_),
    .B(_06707_),
    .Y(_06708_));
 AND3x1_ASAP7_75t_R _24860_ (.A(_18582_),
    .B(_06705_),
    .C(_06708_),
    .Y(_18587_));
 OR3x1_ASAP7_75t_R _24861_ (.A(_01536_),
    .B(_01537_),
    .C(net299),
    .Y(_06709_));
 OR3x1_ASAP7_75t_R _24862_ (.A(net301),
    .B(_06439_),
    .C(_06445_),
    .Y(_06710_));
 NAND2x1_ASAP7_75t_R _24863_ (.A(_06709_),
    .B(_06710_),
    .Y(_06711_));
 AND2x2_ASAP7_75t_R _24864_ (.A(_18587_),
    .B(_06711_),
    .Y(_18589_));
 AOI211x1_ASAP7_75t_R _24865_ (.A1(_01535_),
    .A2(net301),
    .B(_06455_),
    .C(_06463_),
    .Y(_06712_));
 AND5x1_ASAP7_75t_R _24866_ (.A(_18582_),
    .B(_06705_),
    .C(_06708_),
    .D(_06711_),
    .E(_06712_),
    .Y(_18591_));
 AND3x1_ASAP7_75t_R _24867_ (.A(_18590_),
    .B(_06476_),
    .C(_18591_),
    .Y(_18593_));
 AND3x1_ASAP7_75t_R _24868_ (.A(_18592_),
    .B(_06490_),
    .C(_18593_),
    .Y(_18595_));
 AND3x1_ASAP7_75t_R _24869_ (.A(_18594_),
    .B(_06503_),
    .C(_18595_),
    .Y(_18597_));
 AND2x2_ASAP7_75t_R _24870_ (.A(_18596_),
    .B(_06517_),
    .Y(_06713_));
 AND2x2_ASAP7_75t_R _24871_ (.A(_18597_),
    .B(_06713_),
    .Y(_18599_));
 AND4x1_ASAP7_75t_R _24872_ (.A(_18598_),
    .B(_06532_),
    .C(_18597_),
    .D(_06713_),
    .Y(_18601_));
 AND3x1_ASAP7_75t_R _24873_ (.A(_18600_),
    .B(_06545_),
    .C(_18601_),
    .Y(_18603_));
 AND3x1_ASAP7_75t_R _24874_ (.A(_01311_),
    .B(net3302),
    .C(_06229_),
    .Y(_06714_));
 AND4x1_ASAP7_75t_R _24875_ (.A(_00238_),
    .B(_01736_),
    .C(_05552_),
    .D(_06664_),
    .Y(_06715_));
 OA21x2_ASAP7_75t_R _24876_ (.A1(_01717_),
    .A2(_06714_),
    .B(_06715_),
    .Y(_06716_));
 NAND2x1_ASAP7_75t_R _24877_ (.A(_06568_),
    .B(_06716_),
    .Y(core_busy_d));
 AND2x2_ASAP7_75t_R _24878_ (.A(clknet_leaf_26_clk_i),
    .B(\core_clock_gate_i.en_latch ),
    .Y(\core_clock_gate_i.clk_o ));
 INVx1_ASAP7_75t_R _24879_ (.A(net3963),
    .Y(_06717_));
 NAND2x1_ASAP7_75t_R _24880_ (.A(net3965),
    .B(net150),
    .Y(_00008_));
 AND2x2_ASAP7_75t_R _24881_ (.A(net2759),
    .B(net249),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 AND3x1_ASAP7_75t_R _24882_ (.A(_00240_),
    .B(net2696),
    .C(net2688),
    .Y(_06718_));
 TAPCELL_ASAP7_75t_R TAP_878 ();
 OA211x2_ASAP7_75t_R _24884_ (.A1(_01845_),
    .A2(_01846_),
    .B(_06589_),
    .C(_01814_),
    .Y(_06720_));
 NOR2x1_ASAP7_75t_R _24885_ (.A(_06592_),
    .B(_06720_),
    .Y(_06721_));
 OR3x4_ASAP7_75t_R _24886_ (.A(_06580_),
    .B(_06718_),
    .C(_06721_),
    .Y(_06722_));
 AND3x4_ASAP7_75t_R _24887_ (.A(_06668_),
    .B(net3106),
    .C(_06722_),
    .Y(_06723_));
 NAND2x2_ASAP7_75t_R _24888_ (.A(_06618_),
    .B(_06723_),
    .Y(_06724_));
 TAPCELL_ASAP7_75t_R TAP_877 ();
 TAPCELL_ASAP7_75t_R TAP_876 ();
 AND3x4_ASAP7_75t_R _24891_ (.A(net2739),
    .B(_06570_),
    .C(_01737_),
    .Y(_06727_));
 AND2x2_ASAP7_75t_R _24892_ (.A(_06589_),
    .B(_06727_),
    .Y(_06728_));
 CKINVDCx20_ASAP7_75t_R _24893_ (.A(_01815_),
    .Y(_06729_));
 AND3x4_ASAP7_75t_R _24894_ (.A(_06729_),
    .B(_06618_),
    .C(_06723_),
    .Y(_06730_));
 TAPCELL_ASAP7_75t_R TAP_875 ();
 TAPCELL_ASAP7_75t_R TAP_874 ();
 AO21x1_ASAP7_75t_R _24897_ (.A1(_06724_),
    .A2(_06728_),
    .B(_06730_),
    .Y(_06733_));
 CKINVDCx20_ASAP7_75t_R _24898_ (.A(_00239_),
    .Y(_06734_));
 TAPCELL_ASAP7_75t_R TAP_873 ();
 TAPCELL_ASAP7_75t_R TAP_872 ();
 OA21x2_ASAP7_75t_R _24901_ (.A1(_06727_),
    .A2(_06724_),
    .B(_06734_),
    .Y(_06737_));
 OA21x2_ASAP7_75t_R _24902_ (.A1(_06733_),
    .A2(_06737_),
    .B(net300),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 TAPCELL_ASAP7_75t_R TAP_871 ();
 TAPCELL_ASAP7_75t_R TAP_870 ();
 AND3x1_ASAP7_75t_R _24905_ (.A(_00239_),
    .B(_06618_),
    .C(_06723_),
    .Y(_06740_));
 AO21x1_ASAP7_75t_R _24906_ (.A1(_06678_),
    .A2(_06724_),
    .B(_06740_),
    .Y(_06741_));
 TAPCELL_ASAP7_75t_R TAP_869 ();
 TAPCELL_ASAP7_75t_R TAP_868 ();
 AOI221x1_ASAP7_75t_R _24909_ (.A1(_06678_),
    .A2(_06740_),
    .B1(_06741_),
    .B2(_00240_),
    .C(net299),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 AO21x1_ASAP7_75t_R _24910_ (.A1(_06734_),
    .A2(_06727_),
    .B(_06729_),
    .Y(_06744_));
 AND3x1_ASAP7_75t_R _24911_ (.A(net300),
    .B(_06724_),
    .C(_06744_),
    .Y(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 INVx1_ASAP7_75t_R _24912_ (.A(_00660_),
    .Y(\cs_registers_i.mhpmcounter[2][0] ));
 INVx1_ASAP7_75t_R _24913_ (.A(_00659_),
    .Y(\cs_registers_i.mcycle_counter_i.counter[0] ));
 INVx1_ASAP7_75t_R _24914_ (.A(_17754_),
    .Y(\cs_registers_i.pc_if_i[2] ));
 INVx1_ASAP7_75t_R _24915_ (.A(_17819_),
    .Y(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ));
 NAND2x1_ASAP7_75t_R _24916_ (.A(net2285),
    .B(_05883_),
    .Y(_16994_));
 TAPCELL_ASAP7_75t_R TAP_867 ();
 NAND2x1_ASAP7_75t_R _24918_ (.A(_05859_),
    .B(net2316),
    .Y(_17002_));
 TAPCELL_ASAP7_75t_R TAP_866 ();
 NAND2x1_ASAP7_75t_R _24920_ (.A(_05926_),
    .B(net2187),
    .Y(_17016_));
 TAPCELL_ASAP7_75t_R TAP_865 ();
 NAND2x1_ASAP7_75t_R _24922_ (.A(net2285),
    .B(_05972_),
    .Y(_17034_));
 NAND2x1_ASAP7_75t_R _24923_ (.A(_05859_),
    .B(net2364),
    .Y(_17044_));
 NAND2x1_ASAP7_75t_R _24924_ (.A(_05938_),
    .B(net2188),
    .Y(_17061_));
 NAND2x1_ASAP7_75t_R _24925_ (.A(net2349),
    .B(_05972_),
    .Y(_17082_));
 TAPCELL_ASAP7_75t_R TAP_864 ();
 NAND2x1_ASAP7_75t_R _24927_ (.A(_05867_),
    .B(net2365),
    .Y(_17091_));
 TAPCELL_ASAP7_75t_R TAP_863 ();
 NAND2x1_ASAP7_75t_R _24929_ (.A(net2246),
    .B(_05959_),
    .Y(_17107_));
 NAND2x2_ASAP7_75t_R _24930_ (.A(_05930_),
    .B(_05951_),
    .Y(_17712_));
 NAND2x1_ASAP7_75t_R _24931_ (.A(_05840_),
    .B(net2243),
    .Y(_16765_));
 NAND2x1_ASAP7_75t_R _24932_ (.A(_05845_),
    .B(net2243),
    .Y(_16768_));
 NAND2x1_ASAP7_75t_R _24933_ (.A(_05855_),
    .B(net2243),
    .Y(_16775_));
 NAND2x1_ASAP7_75t_R _24934_ (.A(_05863_),
    .B(_05964_),
    .Y(_16789_));
 NAND2x1_ASAP7_75t_R _24935_ (.A(_05870_),
    .B(net2243),
    .Y(_16810_));
 NAND2x1_ASAP7_75t_R _24936_ (.A(_05879_),
    .B(_05964_),
    .Y(_16829_));
 NAND2x1_ASAP7_75t_R _24937_ (.A(_05840_),
    .B(_05867_),
    .Y(_16843_));
 NAND2x2_ASAP7_75t_R _24938_ (.A(_05887_),
    .B(_05964_),
    .Y(_16855_));
 NAND2x1_ASAP7_75t_R _24939_ (.A(net2337),
    .B(_05867_),
    .Y(_16873_));
 NAND2x1_ASAP7_75t_R _24940_ (.A(_05894_),
    .B(_05964_),
    .Y(_16882_));
 NAND2x1_ASAP7_75t_R _24941_ (.A(net2345),
    .B(_05867_),
    .Y(_16897_));
 NAND2x2_ASAP7_75t_R _24942_ (.A(_05904_),
    .B(net2186),
    .Y(_16910_));
 NAND2x1_ASAP7_75t_R _24943_ (.A(_05840_),
    .B(_05972_),
    .Y(_16927_));
 NAND2x1_ASAP7_75t_R _24944_ (.A(net2285),
    .B(_05867_),
    .Y(_16930_));
 NAND2x1_ASAP7_75t_R _24945_ (.A(_05912_),
    .B(net2189),
    .Y(_16943_));
 NAND2x1_ASAP7_75t_R _24946_ (.A(net2338),
    .B(_05972_),
    .Y(_16959_));
 NAND2x1_ASAP7_75t_R _24947_ (.A(_05867_),
    .B(_05870_),
    .Y(_16962_));
 NAND2x1_ASAP7_75t_R _24948_ (.A(_05917_),
    .B(net2185),
    .Y(_16977_));
 NAND2x1_ASAP7_75t_R _24949_ (.A(net2338),
    .B(_05908_),
    .Y(_17031_));
 NAND2x1_ASAP7_75t_R _24950_ (.A(_05870_),
    .B(_05883_),
    .Y(_17035_));
 NAND2x1_ASAP7_75t_R _24951_ (.A(_05867_),
    .B(net2318),
    .Y(_17045_));
 NAND2x1_ASAP7_75t_R _24952_ (.A(net2245),
    .B(_05955_),
    .Y(_17062_));
 NAND2x1_ASAP7_75t_R _24953_ (.A(net2355),
    .B(net2190),
    .Y(_17083_));
 NAND2x1_ASAP7_75t_R _24954_ (.A(_05859_),
    .B(net2324),
    .Y(_17092_));
 OA22x2_ASAP7_75t_R _24955_ (.A1(_01314_),
    .A2(_01677_),
    .B1(_05548_),
    .B2(_00816_),
    .Y(_17122_));
 NAND2x1_ASAP7_75t_R _24956_ (.A(net2349),
    .B(_05900_),
    .Y(_17133_));
 NAND2x1_ASAP7_75t_R _24957_ (.A(_05874_),
    .B(net2365),
    .Y(_17142_));
 NAND2x1_ASAP7_75t_R _24958_ (.A(net2223),
    .B(_05955_),
    .Y(_17159_));
 OR2x2_ASAP7_75t_R _24959_ (.A(_05840_),
    .B(_05946_),
    .Y(_17177_));
 NAND2x1_ASAP7_75t_R _24960_ (.A(net2318),
    .B(_05972_),
    .Y(_17188_));
 NAND2x1_ASAP7_75t_R _24961_ (.A(_05867_),
    .B(net2271),
    .Y(_17199_));
 OR2x2_ASAP7_75t_R _24962_ (.A(net2340),
    .B(_05946_),
    .Y(_17227_));
 NAND2x1_ASAP7_75t_R _24963_ (.A(net2365),
    .B(_05972_),
    .Y(_17238_));
 NAND2x1_ASAP7_75t_R _24964_ (.A(_05867_),
    .B(_05917_),
    .Y(_17248_));
 NAND2x1_ASAP7_75t_R _24965_ (.A(net2235),
    .B(_05955_),
    .Y(_17253_));
 OR2x2_ASAP7_75t_R _24966_ (.A(net2348),
    .B(_05946_),
    .Y(_17278_));
 NAND2x1_ASAP7_75t_R _24967_ (.A(net2324),
    .B(_05972_),
    .Y(_17289_));
 NAND2x1_ASAP7_75t_R _24968_ (.A(_05867_),
    .B(_05926_),
    .Y(_17299_));
 NAND2x1_ASAP7_75t_R _24969_ (.A(net2234),
    .B(_05959_),
    .Y(_17304_));
 OR2x2_ASAP7_75t_R _24970_ (.A(net2287),
    .B(_05946_),
    .Y(_17322_));
 NAND2x1_ASAP7_75t_R _24971_ (.A(net2271),
    .B(_05972_),
    .Y(_17333_));
 NAND2x1_ASAP7_75t_R _24972_ (.A(_05867_),
    .B(_05938_),
    .Y(_17343_));
 OR2x2_ASAP7_75t_R _24973_ (.A(net2351),
    .B(_05946_),
    .Y(_17366_));
 NAND2x1_ASAP7_75t_R _24974_ (.A(net2368),
    .B(_05933_),
    .Y(_17371_));
 NAND2x1_ASAP7_75t_R _24975_ (.A(_05917_),
    .B(_05972_),
    .Y(_17378_));
 NAND2x1_ASAP7_75t_R _24976_ (.A(_05867_),
    .B(_05955_),
    .Y(_17388_));
 OR2x2_ASAP7_75t_R _24977_ (.A(net2356),
    .B(_05946_),
    .Y(_17414_));
 NAND2x1_ASAP7_75t_R _24978_ (.A(net2328),
    .B(_05933_),
    .Y(_17419_));
 NAND2x1_ASAP7_75t_R _24979_ (.A(_05926_),
    .B(_05972_),
    .Y(_17426_));
 NAND2x1_ASAP7_75t_R _24980_ (.A(_05867_),
    .B(_05959_),
    .Y(_17435_));
 OR2x2_ASAP7_75t_R _24981_ (.A(net2320),
    .B(_05946_),
    .Y(_17457_));
 NAND2x1_ASAP7_75t_R _24982_ (.A(net2273),
    .B(_05933_),
    .Y(_17462_));
 NAND2x1_ASAP7_75t_R _24983_ (.A(net2308),
    .B(_05972_),
    .Y(_17469_));
 OR2x2_ASAP7_75t_R _24984_ (.A(net2367),
    .B(_05946_),
    .Y(_17493_));
 NAND2x1_ASAP7_75t_R _24985_ (.A(_05917_),
    .B(_05933_),
    .Y(_17498_));
 NAND2x1_ASAP7_75t_R _24986_ (.A(_05955_),
    .B(_05972_),
    .Y(_17505_));
 OR2x2_ASAP7_75t_R _24987_ (.A(net2328),
    .B(_05946_),
    .Y(_17535_));
 NAND2x1_ASAP7_75t_R _24988_ (.A(_05926_),
    .B(_05933_),
    .Y(_17540_));
 NAND2x1_ASAP7_75t_R _24989_ (.A(_05959_),
    .B(_05972_),
    .Y(_17547_));
 OR2x2_ASAP7_75t_R _24990_ (.A(net2275),
    .B(_05946_),
    .Y(_17569_));
 NAND2x1_ASAP7_75t_R _24991_ (.A(_05933_),
    .B(net2305),
    .Y(_17574_));
 OR2x2_ASAP7_75t_R _24992_ (.A(_05917_),
    .B(_05946_),
    .Y(_17601_));
 NAND2x1_ASAP7_75t_R _24993_ (.A(_05933_),
    .B(_05955_),
    .Y(_17606_));
 OR2x2_ASAP7_75t_R _24994_ (.A(_05926_),
    .B(_05946_),
    .Y(_17631_));
 NAND2x1_ASAP7_75t_R _24995_ (.A(_05933_),
    .B(_05959_),
    .Y(_17636_));
 OR2x2_ASAP7_75t_R _24996_ (.A(net2305),
    .B(_05946_),
    .Y(_17659_));
 OR2x2_ASAP7_75t_R _24997_ (.A(_05946_),
    .B(_05955_),
    .Y(_17681_));
 OR2x2_ASAP7_75t_R _24998_ (.A(_05946_),
    .B(_05959_),
    .Y(_17711_));
 NAND2x1_ASAP7_75t_R _24999_ (.A(_05821_),
    .B(_05845_),
    .Y(_16766_));
 NAND2x1_ASAP7_75t_R _25000_ (.A(_05821_),
    .B(_05855_),
    .Y(_16769_));
 NAND2x1_ASAP7_75t_R _25001_ (.A(_05821_),
    .B(_05863_),
    .Y(_16776_));
 NAND2x1_ASAP7_75t_R _25002_ (.A(_05821_),
    .B(_05870_),
    .Y(_16790_));
 NAND2x1_ASAP7_75t_R _25003_ (.A(_05821_),
    .B(_05879_),
    .Y(_16811_));
 NAND2x1_ASAP7_75t_R _25004_ (.A(_05821_),
    .B(_05887_),
    .Y(_16830_));
 NAND2x1_ASAP7_75t_R _25005_ (.A(net2337),
    .B(_05859_),
    .Y(_16844_));
 NAND2x1_ASAP7_75t_R _25006_ (.A(_05821_),
    .B(_05894_),
    .Y(_16856_));
 NAND2x1_ASAP7_75t_R _25007_ (.A(net2345),
    .B(_05859_),
    .Y(_16874_));
 NAND2x1_ASAP7_75t_R _25008_ (.A(_05821_),
    .B(_05904_),
    .Y(_16883_));
 NAND2x1_ASAP7_75t_R _25009_ (.A(_05859_),
    .B(net2285),
    .Y(_16898_));
 NAND2x1_ASAP7_75t_R _25010_ (.A(net2245),
    .B(_05912_),
    .Y(_16911_));
 NAND2x1_ASAP7_75t_R _25011_ (.A(net2341),
    .B(_05883_),
    .Y(_16928_));
 NAND2x1_ASAP7_75t_R _25012_ (.A(_05859_),
    .B(_05870_),
    .Y(_16931_));
 NAND2x1_ASAP7_75t_R _25013_ (.A(net2245),
    .B(_05917_),
    .Y(_16944_));
 NAND2x1_ASAP7_75t_R _25014_ (.A(net2345),
    .B(_05883_),
    .Y(_16960_));
 NAND2x1_ASAP7_75t_R _25015_ (.A(_05859_),
    .B(net2353),
    .Y(_16963_));
 NAND2x1_ASAP7_75t_R _25016_ (.A(net2247),
    .B(_05926_),
    .Y(_16978_));
 NAND2x1_ASAP7_75t_R _25017_ (.A(net2347),
    .B(_05972_),
    .Y(_16996_));
 NAND2x1_ASAP7_75t_R _25018_ (.A(_05867_),
    .B(net2353),
    .Y(_17004_));
 NAND2x1_ASAP7_75t_R _25019_ (.A(net2245),
    .B(_05938_),
    .Y(_17018_));
 NAND2x1_ASAP7_75t_R _25020_ (.A(_05840_),
    .B(_05933_),
    .Y(_17032_));
 NAND2x1_ASAP7_75t_R _25021_ (.A(_05955_),
    .B(net2185),
    .Y(_17109_));
 OR2x2_ASAP7_75t_R _25022_ (.A(_05827_),
    .B(_05946_),
    .Y(_17123_));
 NAND2x1_ASAP7_75t_R _25023_ (.A(net2355),
    .B(_05972_),
    .Y(_17134_));
 NAND2x1_ASAP7_75t_R _25024_ (.A(_05867_),
    .B(net2324),
    .Y(_17143_));
 NAND2x1_ASAP7_75t_R _25025_ (.A(_05959_),
    .B(net2185),
    .Y(_17160_));
 OA211x2_ASAP7_75t_R _25026_ (.A1(_05982_),
    .A2(_05983_),
    .B(_05985_),
    .C(_00025_),
    .Y(_06750_));
 OA21x2_ASAP7_75t_R _25027_ (.A1(net2236),
    .A2(_06750_),
    .B(_02342_),
    .Y(_17175_));
 TAPCELL_ASAP7_75t_R TAP_862 ();
 NAND2x1_ASAP7_75t_R _25029_ (.A(net2340),
    .B(_05930_),
    .Y(_17178_));
 NAND2x1_ASAP7_75t_R _25030_ (.A(net2190),
    .B(net2365),
    .Y(_17189_));
 NAND2x1_ASAP7_75t_R _25031_ (.A(_05859_),
    .B(_05917_),
    .Y(_17200_));
 NAND2x1_ASAP7_75t_R _25032_ (.A(net2348),
    .B(_05930_),
    .Y(_17228_));
 NAND2x1_ASAP7_75t_R _25033_ (.A(net2191),
    .B(net2325),
    .Y(_17239_));
 NAND2x1_ASAP7_75t_R _25034_ (.A(_05859_),
    .B(_05926_),
    .Y(_17249_));
 NAND2x1_ASAP7_75t_R _25035_ (.A(net2296),
    .B(_05959_),
    .Y(_17254_));
 NAND2x1_ASAP7_75t_R _25036_ (.A(net2286),
    .B(_05930_),
    .Y(_17279_));
 NAND2x1_ASAP7_75t_R _25037_ (.A(net2190),
    .B(net2271),
    .Y(_17290_));
 NAND2x1_ASAP7_75t_R _25038_ (.A(_05859_),
    .B(_05938_),
    .Y(_17300_));
 NAND2x1_ASAP7_75t_R _25039_ (.A(net2350),
    .B(_05930_),
    .Y(_17323_));
 NAND2x1_ASAP7_75t_R _25040_ (.A(net2192),
    .B(_05917_),
    .Y(_17334_));
 NAND2x1_ASAP7_75t_R _25041_ (.A(_05859_),
    .B(_05955_),
    .Y(_17344_));
 NAND2x1_ASAP7_75t_R _25042_ (.A(net2356),
    .B(_05930_),
    .Y(_17367_));
 NAND2x1_ASAP7_75t_R _25043_ (.A(net2327),
    .B(_05908_),
    .Y(_17372_));
 NAND2x1_ASAP7_75t_R _25044_ (.A(net2190),
    .B(_05926_),
    .Y(_17379_));
 NAND2x1_ASAP7_75t_R _25045_ (.A(_05859_),
    .B(_05959_),
    .Y(_17389_));
 NAND2x1_ASAP7_75t_R _25046_ (.A(net2320),
    .B(_05930_),
    .Y(_17415_));
 NAND2x1_ASAP7_75t_R _25047_ (.A(_05908_),
    .B(net2272),
    .Y(_17420_));
 NAND2x1_ASAP7_75t_R _25048_ (.A(net2190),
    .B(net2308),
    .Y(_17427_));
 NAND2x1_ASAP7_75t_R _25049_ (.A(net2366),
    .B(_05930_),
    .Y(_17458_));
 NAND2x1_ASAP7_75t_R _25050_ (.A(_05908_),
    .B(_05917_),
    .Y(_17463_));
 NAND2x1_ASAP7_75t_R _25051_ (.A(net2190),
    .B(_05955_),
    .Y(_17470_));
 NAND2x1_ASAP7_75t_R _25052_ (.A(net2328),
    .B(_05930_),
    .Y(_17494_));
 NAND2x1_ASAP7_75t_R _25053_ (.A(_05908_),
    .B(_05926_),
    .Y(_17499_));
 NAND2x1_ASAP7_75t_R _25054_ (.A(net2190),
    .B(_05959_),
    .Y(_17506_));
 NAND2x1_ASAP7_75t_R _25055_ (.A(net2275),
    .B(_05930_),
    .Y(_17536_));
 NAND2x1_ASAP7_75t_R _25056_ (.A(_05908_),
    .B(net2307),
    .Y(_17541_));
 NAND2x1_ASAP7_75t_R _25057_ (.A(_05917_),
    .B(_05930_),
    .Y(_17570_));
 NAND2x1_ASAP7_75t_R _25058_ (.A(_05908_),
    .B(_05955_),
    .Y(_17575_));
 NAND2x1_ASAP7_75t_R _25059_ (.A(_05926_),
    .B(_05930_),
    .Y(_17602_));
 NAND2x1_ASAP7_75t_R _25060_ (.A(_05908_),
    .B(_05959_),
    .Y(_17607_));
 NAND2x1_ASAP7_75t_R _25061_ (.A(_05930_),
    .B(net2306),
    .Y(_17632_));
 NAND2x1_ASAP7_75t_R _25062_ (.A(_05930_),
    .B(_05955_),
    .Y(_17660_));
 NAND2x1_ASAP7_75t_R _25063_ (.A(_05930_),
    .B(_05959_),
    .Y(_17682_));
 NAND2x2_ASAP7_75t_R _25064_ (.A(_05454_),
    .B(_05943_),
    .Y(_06752_));
 OR3x4_ASAP7_75t_R _25065_ (.A(_05813_),
    .B(_06752_),
    .C(_05951_),
    .Y(_17736_));
 TAPCELL_ASAP7_75t_R TAP_861 ();
 TAPCELL_ASAP7_75t_R TAP_860 ();
 OR3x1_ASAP7_75t_R _25068_ (.A(_00663_),
    .B(net309),
    .C(_13815_),
    .Y(_06755_));
 OAI21x1_ASAP7_75t_R _25069_ (.A1(_13817_),
    .A2(_18336_),
    .B(_06755_),
    .Y(_17758_));
 TAPCELL_ASAP7_75t_R TAP_859 ();
 TAPCELL_ASAP7_75t_R TAP_858 ();
 XNOR2x1_ASAP7_75t_R _25072_ (.B(_14296_),
    .Y(_06758_),
    .A(_13620_));
 TAPCELL_ASAP7_75t_R TAP_857 ();
 INVx2_ASAP7_75t_R _25074_ (.A(_00668_),
    .Y(_06760_));
 INVx1_ASAP7_75t_R _25075_ (.A(_01448_),
    .Y(_06761_));
 OA222x2_ASAP7_75t_R _25076_ (.A1(_00285_),
    .A2(_06760_),
    .B1(_06761_),
    .B2(_13815_),
    .C1(_13986_),
    .C2(net2218),
    .Y(_06762_));
 OA211x2_ASAP7_75t_R _25077_ (.A1(_00284_),
    .A2(net2322),
    .B(_06762_),
    .C(_13817_),
    .Y(_06763_));
 AOI21x1_ASAP7_75t_R _25078_ (.A1(net309),
    .A2(_06758_),
    .B(_06763_),
    .Y(_17762_));
 XOR2x1_ASAP7_75t_R _25079_ (.A(_13620_),
    .Y(_06764_),
    .B(_18353_));
 INVx1_ASAP7_75t_R _25080_ (.A(_00672_),
    .Y(_06765_));
 INVx1_ASAP7_75t_R _25081_ (.A(_01446_),
    .Y(_06766_));
 OA222x2_ASAP7_75t_R _25082_ (.A1(_00285_),
    .A2(_06765_),
    .B1(_06766_),
    .B2(_13815_),
    .C1(_13986_),
    .C2(_14420_),
    .Y(_06767_));
 OA211x2_ASAP7_75t_R _25083_ (.A1(_00284_),
    .A2(_15167_),
    .B(_06767_),
    .C(_13817_),
    .Y(_06768_));
 AOI21x1_ASAP7_75t_R _25084_ (.A1(net309),
    .A2(_06764_),
    .B(_06768_),
    .Y(_17766_));
 AO221x1_ASAP7_75t_R _25085_ (.A1(_13775_),
    .A2(_00674_),
    .B1(_01445_),
    .B2(_13778_),
    .C(net309),
    .Y(_06769_));
 AO221x1_ASAP7_75t_R _25086_ (.A1(_13772_),
    .A2(_05629_),
    .B1(_05885_),
    .B2(_05781_),
    .C(_06769_),
    .Y(_06770_));
 OAI21x1_ASAP7_75t_R _25087_ (.A1(_13620_),
    .A2(_14481_),
    .B(net309),
    .Y(_06771_));
 AO22x2_ASAP7_75t_R _25088_ (.A1(_14002_),
    .A2(_14481_),
    .B1(_06770_),
    .B2(_06771_),
    .Y(_16728_));
 NOR2x1_ASAP7_75t_R _25089_ (.A(_00284_),
    .B(_15279_),
    .Y(_06772_));
 TAPCELL_ASAP7_75t_R TAP_856 ();
 AO221x1_ASAP7_75t_R _25091_ (.A1(_13775_),
    .A2(_00677_),
    .B1(_01444_),
    .B2(_13778_),
    .C(net309),
    .Y(_06774_));
 AO21x1_ASAP7_75t_R _25092_ (.A1(_13772_),
    .A2(_14540_),
    .B(_06774_),
    .Y(_06775_));
 NOR2x1_ASAP7_75t_R _25093_ (.A(_14002_),
    .B(_18363_),
    .Y(_06776_));
 AO21x1_ASAP7_75t_R _25094_ (.A1(_13620_),
    .A2(_18363_),
    .B(_06776_),
    .Y(_06777_));
 OA21x2_ASAP7_75t_R _25095_ (.A1(_06772_),
    .A2(_06775_),
    .B(_06777_),
    .Y(_17768_));
 OR3x1_ASAP7_75t_R _25096_ (.A(_00682_),
    .B(net309),
    .C(_13815_),
    .Y(_06778_));
 OAI21x1_ASAP7_75t_R _25097_ (.A1(_13817_),
    .A2(_18376_),
    .B(_06778_),
    .Y(_17772_));
 AO221x1_ASAP7_75t_R _25098_ (.A1(_13775_),
    .A2(_00686_),
    .B1(_02221_),
    .B2(_13778_),
    .C(net309),
    .Y(_06779_));
 TAPCELL_ASAP7_75t_R TAP_855 ();
 OAI22x1_ASAP7_75t_R _25100_ (.A1(_00284_),
    .A2(_14099_),
    .B1(_15487_),
    .B2(_13986_),
    .Y(_06781_));
 OAI21x1_ASAP7_75t_R _25101_ (.A1(_13620_),
    .A2(_18384_),
    .B(net309),
    .Y(_06782_));
 OA21x2_ASAP7_75t_R _25102_ (.A1(_06779_),
    .A2(_06781_),
    .B(_06782_),
    .Y(_06783_));
 AO21x1_ASAP7_75t_R _25103_ (.A1(_14002_),
    .A2(_18384_),
    .B(_06783_),
    .Y(_17776_));
 TAPCELL_ASAP7_75t_R TAP_854 ();
 OAI21x1_ASAP7_75t_R _25105_ (.A1(_13620_),
    .A2(_18395_),
    .B(net308),
    .Y(_06785_));
 AO221x1_ASAP7_75t_R _25106_ (.A1(_13775_),
    .A2(_00750_),
    .B1(_02219_),
    .B2(_13778_),
    .C(net308),
    .Y(_06786_));
 AOI21x1_ASAP7_75t_R _25107_ (.A1(_13772_),
    .A2(_15723_),
    .B(_06786_),
    .Y(_06787_));
 OAI21x1_ASAP7_75t_R _25108_ (.A1(_00284_),
    .A2(_15773_),
    .B(_06787_),
    .Y(_06788_));
 AO22x1_ASAP7_75t_R _25109_ (.A1(_14002_),
    .A2(_18395_),
    .B1(_06785_),
    .B2(_06788_),
    .Y(_17780_));
 NOR2x1_ASAP7_75t_R _25110_ (.A(_00284_),
    .B(_05957_),
    .Y(_06789_));
 AO221x1_ASAP7_75t_R _25111_ (.A1(_13775_),
    .A2(_00783_),
    .B1(_02218_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_06790_));
 OA22x2_ASAP7_75t_R _25112_ (.A1(_13986_),
    .A2(_15839_),
    .B1(_06789_),
    .B2(_06790_),
    .Y(_06791_));
 OAI22x1_ASAP7_75t_R _25113_ (.A1(_13620_),
    .A2(_15841_),
    .B1(_06791_),
    .B2(net308),
    .Y(_06792_));
 AOI21x1_ASAP7_75t_R _25114_ (.A1(_14002_),
    .A2(_15841_),
    .B(_06792_),
    .Y(_16740_));
 OR3x1_ASAP7_75t_R _25115_ (.A(_00816_),
    .B(net308),
    .C(_13815_),
    .Y(_06793_));
 OAI21x1_ASAP7_75t_R _25116_ (.A1(_13817_),
    .A2(_18404_),
    .B(_06793_),
    .Y(_17782_));
 XNOR2x1_ASAP7_75t_R _25117_ (.B(_18415_),
    .Y(_06794_),
    .A(_13620_));
 AO222x2_ASAP7_75t_R _25118_ (.A1(_13775_),
    .A2(_00881_),
    .B1(_02215_),
    .B2(_13778_),
    .C1(_16261_),
    .C2(_05781_),
    .Y(_06795_));
 NOR2x1_ASAP7_75t_R _25119_ (.A(_13986_),
    .B(_16213_),
    .Y(_06796_));
 OR3x1_ASAP7_75t_R _25120_ (.A(net309),
    .B(_06795_),
    .C(_06796_),
    .Y(_06797_));
 OA21x2_ASAP7_75t_R _25121_ (.A1(_13817_),
    .A2(_06794_),
    .B(_06797_),
    .Y(_17786_));
 TAPCELL_ASAP7_75t_R TAP_853 ();
 OR3x1_ASAP7_75t_R _25123_ (.A(_00946_),
    .B(net309),
    .C(_13815_),
    .Y(_06799_));
 OAI21x1_ASAP7_75t_R _25124_ (.A1(_13817_),
    .A2(_18424_),
    .B(_06799_),
    .Y(_17790_));
 OR3x1_ASAP7_75t_R _25125_ (.A(_00979_),
    .B(net309),
    .C(_13815_),
    .Y(_06800_));
 OAI21x1_ASAP7_75t_R _25126_ (.A1(_13817_),
    .A2(_18429_),
    .B(_06800_),
    .Y(_16750_));
 OA21x2_ASAP7_75t_R _25127_ (.A1(_00915_),
    .A2(_16747_),
    .B(_00948_),
    .Y(_06801_));
 OAI21x1_ASAP7_75t_R _25128_ (.A1(_00947_),
    .A2(_06801_),
    .B(_02277_),
    .Y(_16749_));
 XOR2x1_ASAP7_75t_R _25129_ (.A(_13620_),
    .Y(_06802_),
    .B(_18434_));
 AOI22x1_ASAP7_75t_R _25130_ (.A1(_13775_),
    .A2(_01011_),
    .B1(_02211_),
    .B2(_13778_),
    .Y(_06803_));
 OA21x2_ASAP7_75t_R _25131_ (.A1(_00284_),
    .A2(_05877_),
    .B(_06803_),
    .Y(_06804_));
 OA211x2_ASAP7_75t_R _25132_ (.A1(_13986_),
    .A2(_06148_),
    .B(_06804_),
    .C(_13817_),
    .Y(_06805_));
 AOI21x1_ASAP7_75t_R _25133_ (.A1(net309),
    .A2(_06802_),
    .B(_06805_),
    .Y(_17792_));
 AOI22x1_ASAP7_75t_R _25134_ (.A1(_13775_),
    .A2(_01077_),
    .B1(_02209_),
    .B2(_13778_),
    .Y(_06806_));
 OA211x2_ASAP7_75t_R _25135_ (.A1(_13986_),
    .A2(_04697_),
    .B(_06806_),
    .C(_13817_),
    .Y(_06807_));
 OA21x2_ASAP7_75t_R _25136_ (.A1(_00284_),
    .A2(_05892_),
    .B(_06807_),
    .Y(_06808_));
 AOI21x1_ASAP7_75t_R _25137_ (.A1(_14002_),
    .A2(_04700_),
    .B(_06808_),
    .Y(_06809_));
 OA21x2_ASAP7_75t_R _25138_ (.A1(_13620_),
    .A2(_04700_),
    .B(_06809_),
    .Y(_17796_));
 OR3x1_ASAP7_75t_R _25139_ (.A(_01110_),
    .B(net309),
    .C(_13815_),
    .Y(_06810_));
 OAI21x1_ASAP7_75t_R _25140_ (.A1(_13817_),
    .A2(_18449_),
    .B(_06810_),
    .Y(_16756_));
 OR3x1_ASAP7_75t_R _25141_ (.A(_01078_),
    .B(_01046_),
    .C(_16752_),
    .Y(_06811_));
 NAND2x1_ASAP7_75t_R _25142_ (.A(_05520_),
    .B(_06811_),
    .Y(_16755_));
 AO221x1_ASAP7_75t_R _25143_ (.A1(_13775_),
    .A2(_01142_),
    .B1(_02207_),
    .B2(_13778_),
    .C(net308),
    .Y(_06812_));
 OAI22x1_ASAP7_75t_R _25144_ (.A1(_13986_),
    .A2(_04916_),
    .B1(_04965_),
    .B2(_00284_),
    .Y(_06813_));
 OAI21x1_ASAP7_75t_R _25145_ (.A1(_13620_),
    .A2(_04919_),
    .B(net308),
    .Y(_06814_));
 OA21x2_ASAP7_75t_R _25146_ (.A1(_06812_),
    .A2(_06813_),
    .B(_06814_),
    .Y(_06815_));
 AO21x1_ASAP7_75t_R _25147_ (.A1(_14002_),
    .A2(_04919_),
    .B(_06815_),
    .Y(_17798_));
 AO221x1_ASAP7_75t_R _25148_ (.A1(_13775_),
    .A2(_01176_),
    .B1(_02206_),
    .B2(_13778_),
    .C(net309),
    .Y(_06816_));
 AOI21x1_ASAP7_75t_R _25149_ (.A1(_13772_),
    .A2(_05028_),
    .B(_06816_),
    .Y(_06817_));
 OA21x2_ASAP7_75t_R _25150_ (.A1(_00284_),
    .A2(_05075_),
    .B(_06817_),
    .Y(_06818_));
 AOI21x1_ASAP7_75t_R _25151_ (.A1(_14002_),
    .A2(_05030_),
    .B(_06818_),
    .Y(_06819_));
 OA21x2_ASAP7_75t_R _25152_ (.A1(_13620_),
    .A2(_05030_),
    .B(_06819_),
    .Y(_16758_));
 NOR2x1_ASAP7_75t_R _25153_ (.A(_00284_),
    .B(_05924_),
    .Y(_06820_));
 AO221x1_ASAP7_75t_R _25154_ (.A1(_13775_),
    .A2(_01208_),
    .B1(_02205_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_06821_));
 OA22x2_ASAP7_75t_R _25155_ (.A1(_13986_),
    .A2(_05136_),
    .B1(_06820_),
    .B2(_06821_),
    .Y(_06822_));
 OAI22x1_ASAP7_75t_R _25156_ (.A1(_13620_),
    .A2(_05138_),
    .B1(_06822_),
    .B2(net309),
    .Y(_06823_));
 AOI21x1_ASAP7_75t_R _25157_ (.A1(_14002_),
    .A2(_05138_),
    .B(_06823_),
    .Y(_17800_));
 AOI22x1_ASAP7_75t_R _25158_ (.A1(_13775_),
    .A2(_01242_),
    .B1(_02204_),
    .B2(_13778_),
    .Y(_06824_));
 OA211x2_ASAP7_75t_R _25159_ (.A1(_13986_),
    .A2(_05244_),
    .B(_06824_),
    .C(_13817_),
    .Y(_06825_));
 OA21x2_ASAP7_75t_R _25160_ (.A1(_00284_),
    .A2(_05936_),
    .B(_06825_),
    .Y(_06826_));
 AOI21x1_ASAP7_75t_R _25161_ (.A1(_14002_),
    .A2(_05247_),
    .B(_06826_),
    .Y(_06827_));
 OA21x2_ASAP7_75t_R _25162_ (.A1(_13620_),
    .A2(_05247_),
    .B(_06827_),
    .Y(_16761_));
 NOR2x1_ASAP7_75t_R _25163_ (.A(_00284_),
    .B(_05400_),
    .Y(_06828_));
 AO221x1_ASAP7_75t_R _25164_ (.A1(_13775_),
    .A2(_01274_),
    .B1(_02203_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_06829_));
 OA22x2_ASAP7_75t_R _25165_ (.A1(_13986_),
    .A2(_05355_),
    .B1(_06828_),
    .B2(_06829_),
    .Y(_06830_));
 OAI22x1_ASAP7_75t_R _25166_ (.A1(_13620_),
    .A2(_05357_),
    .B1(_06830_),
    .B2(net309),
    .Y(_06831_));
 AOI21x1_ASAP7_75t_R _25167_ (.A1(_14002_),
    .A2(_05357_),
    .B(_06831_),
    .Y(_17802_));
 TAPCELL_ASAP7_75t_R TAP_852 ();
 AND2x2_ASAP7_75t_R _25169_ (.A(_14599_),
    .B(_05570_),
    .Y(_17809_));
 NAND2x1_ASAP7_75t_R _25170_ (.A(_18363_),
    .B(_05570_),
    .Y(_17811_));
 AND2x2_ASAP7_75t_R _25171_ (.A(_05827_),
    .B(net2243),
    .Y(_17829_));
 AND2x2_ASAP7_75t_R _25172_ (.A(_05827_),
    .B(_05852_),
    .Y(_17856_));
 INVx1_ASAP7_75t_R _25173_ (.A(_01379_),
    .Y(_16796_));
 INVx1_ASAP7_75t_R _25174_ (.A(_01382_),
    .Y(_16801_));
 AND2x2_ASAP7_75t_R _25175_ (.A(_05827_),
    .B(_05972_),
    .Y(_17912_));
 INVx1_ASAP7_75t_R _25176_ (.A(_01438_),
    .Y(_17944_));
 INVx1_ASAP7_75t_R _25177_ (.A(_05982_),
    .Y(_16992_));
 AND2x2_ASAP7_75t_R _25178_ (.A(_05827_),
    .B(_05933_),
    .Y(_17960_));
 INVx1_ASAP7_75t_R _25179_ (.A(_00020_),
    .Y(_17997_));
 INVx1_ASAP7_75t_R _25180_ (.A(_00042_),
    .Y(_17405_));
 INVx2_ASAP7_75t_R _25181_ (.A(net2129),
    .Y(_17265_));
 INVx2_ASAP7_75t_R _25182_ (.A(_17313_),
    .Y(_17264_));
 INVx1_ASAP7_75t_R _25183_ (.A(_00046_),
    .Y(_17444_));
 INVx3_ASAP7_75t_R _25184_ (.A(net2133),
    .Y(_17396_));
 INVx2_ASAP7_75t_R _25185_ (.A(net2239),
    .Y(_17616_));
 INVx2_ASAP7_75t_R _25186_ (.A(_17642_),
    .Y(_17615_));
 INVx2_ASAP7_75t_R _25187_ (.A(_17689_),
    .Y(_17688_));
 INVx1_ASAP7_75t_R _25188_ (.A(_18390_),
    .Y(_18388_));
 INVx1_ASAP7_75t_R _25189_ (.A(_18405_),
    .Y(_18403_));
 INVx1_ASAP7_75t_R _25190_ (.A(_18410_),
    .Y(_18408_));
 INVx1_ASAP7_75t_R _25191_ (.A(_18415_),
    .Y(_18413_));
 INVx1_ASAP7_75t_R _25192_ (.A(_16386_),
    .Y(_18418_));
 INVx1_ASAP7_75t_R _25193_ (.A(_18425_),
    .Y(_18423_));
 INVx1_ASAP7_75t_R _25194_ (.A(_06722_),
    .Y(_06833_));
 NOR2x1_ASAP7_75t_R _25195_ (.A(_17752_),
    .B(_06833_),
    .Y(_17751_));
 INVx1_ASAP7_75t_R _25196_ (.A(_00243_),
    .Y(_18574_));
 OR2x6_ASAP7_75t_R _25197_ (.A(_06354_),
    .B(_06565_),
    .Y(_06834_));
 TAPCELL_ASAP7_75t_R TAP_851 ();
 TAPCELL_ASAP7_75t_R TAP_850 ();
 INVx1_ASAP7_75t_R _25200_ (.A(_06834_),
    .Y(_18604_));
 XNOR2x1_ASAP7_75t_R _25201_ (.B(_14179_),
    .Y(_06837_),
    .A(_13620_));
 NOR3x2_ASAP7_75t_R _25202_ (.B(_14139_),
    .C(_14168_),
    .Y(_06838_),
    .A(_14122_));
 AO221x1_ASAP7_75t_R _25203_ (.A1(_13775_),
    .A2(_00663_),
    .B1(_01450_),
    .B2(_13778_),
    .C(_13538_),
    .Y(_06839_));
 AOI21x1_ASAP7_75t_R _25204_ (.A1(_13772_),
    .A2(_06838_),
    .B(_06839_),
    .Y(_06840_));
 OAI21x1_ASAP7_75t_R _25205_ (.A1(_00284_),
    .A2(_14921_),
    .B(_06840_),
    .Y(_06841_));
 OA21x2_ASAP7_75t_R _25206_ (.A1(_13817_),
    .A2(_06837_),
    .B(_06841_),
    .Y(_17759_));
 INVx1_ASAP7_75t_R _25207_ (.A(_18344_),
    .Y(_18346_));
 AND3x1_ASAP7_75t_R _25208_ (.A(_06760_),
    .B(_13817_),
    .C(_13778_),
    .Y(_06842_));
 AO21x1_ASAP7_75t_R _25209_ (.A1(net309),
    .A2(_18346_),
    .B(_06842_),
    .Y(_17763_));
 AND3x1_ASAP7_75t_R _25210_ (.A(_06765_),
    .B(_13817_),
    .C(_13778_),
    .Y(_06843_));
 AO21x1_ASAP7_75t_R _25211_ (.A1(net309),
    .A2(_15172_),
    .B(_06843_),
    .Y(_17767_));
 OR3x1_ASAP7_75t_R _25212_ (.A(_00674_),
    .B(net309),
    .C(_13815_),
    .Y(_06844_));
 OAI21x1_ASAP7_75t_R _25213_ (.A1(_13817_),
    .A2(_18361_),
    .B(_06844_),
    .Y(_16729_));
 INVx1_ASAP7_75t_R _25214_ (.A(_00677_),
    .Y(_06845_));
 AND3x1_ASAP7_75t_R _25215_ (.A(_06845_),
    .B(_13817_),
    .C(_13778_),
    .Y(_06846_));
 AO21x1_ASAP7_75t_R _25216_ (.A1(net309),
    .A2(_15280_),
    .B(_06846_),
    .Y(_17769_));
 NOR2x1_ASAP7_75t_R _25217_ (.A(_00284_),
    .B(net2310),
    .Y(_06847_));
 AO221x1_ASAP7_75t_R _25218_ (.A1(_13775_),
    .A2(_00682_),
    .B1(_01442_),
    .B2(_13778_),
    .C(net309),
    .Y(_06848_));
 AO21x1_ASAP7_75t_R _25219_ (.A1(_13772_),
    .A2(_14651_),
    .B(_06848_),
    .Y(_06849_));
 OAI22x1_ASAP7_75t_R _25220_ (.A1(_13620_),
    .A2(_18375_),
    .B1(_06847_),
    .B2(_06849_),
    .Y(_06850_));
 AOI21x1_ASAP7_75t_R _25221_ (.A1(_14002_),
    .A2(_18375_),
    .B(_06850_),
    .Y(_17773_));
 OR3x1_ASAP7_75t_R _25222_ (.A(_00686_),
    .B(net309),
    .C(_13815_),
    .Y(_06851_));
 OAI21x1_ASAP7_75t_R _25223_ (.A1(_13817_),
    .A2(_18385_),
    .B(_06851_),
    .Y(_17777_));
 OR3x1_ASAP7_75t_R _25224_ (.A(_00750_),
    .B(net308),
    .C(_13815_),
    .Y(_06852_));
 OAI21x1_ASAP7_75t_R _25225_ (.A1(_13817_),
    .A2(_18394_),
    .B(_06852_),
    .Y(_17781_));
 INVx1_ASAP7_75t_R _25226_ (.A(_00783_),
    .Y(_06853_));
 AND3x1_ASAP7_75t_R _25227_ (.A(_06853_),
    .B(_13817_),
    .C(_13778_),
    .Y(_06854_));
 AO21x1_ASAP7_75t_R _25228_ (.A1(net308),
    .A2(_15887_),
    .B(_06854_),
    .Y(_16742_));
 XNOR2x1_ASAP7_75t_R _25229_ (.B(_18405_),
    .Y(_06855_),
    .A(_13620_));
 NOR2x1_ASAP7_75t_R _25230_ (.A(_00284_),
    .B(_05823_),
    .Y(_06856_));
 AO22x1_ASAP7_75t_R _25231_ (.A1(_13775_),
    .A2(_00816_),
    .B1(_02217_),
    .B2(_13778_),
    .Y(_06857_));
 OR3x1_ASAP7_75t_R _25232_ (.A(_13772_),
    .B(_06856_),
    .C(_06857_),
    .Y(_06858_));
 OA211x2_ASAP7_75t_R _25233_ (.A1(_13986_),
    .A2(_15972_),
    .B(_06858_),
    .C(_13817_),
    .Y(_06859_));
 AO21x1_ASAP7_75t_R _25234_ (.A1(net308),
    .A2(_06855_),
    .B(_06859_),
    .Y(_17783_));
 OR3x1_ASAP7_75t_R _25235_ (.A(_00881_),
    .B(net308),
    .C(_13815_),
    .Y(_06860_));
 OAI21x1_ASAP7_75t_R _25236_ (.A1(_13817_),
    .A2(_16262_),
    .B(_06860_),
    .Y(_17787_));
 XNOR2x1_ASAP7_75t_R _25237_ (.B(_18425_),
    .Y(_06861_),
    .A(_13620_));
 OAI22x1_ASAP7_75t_R _25238_ (.A1(_13986_),
    .A2(_16456_),
    .B1(_05861_),
    .B2(_00284_),
    .Y(_06862_));
 AO221x1_ASAP7_75t_R _25239_ (.A1(_13775_),
    .A2(_00946_),
    .B1(_02213_),
    .B2(_13778_),
    .C(net309),
    .Y(_06863_));
 OA22x2_ASAP7_75t_R _25240_ (.A1(_13817_),
    .A2(_06861_),
    .B1(_06862_),
    .B2(_06863_),
    .Y(_17791_));
 AO221x1_ASAP7_75t_R _25241_ (.A1(_13775_),
    .A2(_00979_),
    .B1(_02212_),
    .B2(_13778_),
    .C(net308),
    .Y(_06864_));
 AOI21x1_ASAP7_75t_R _25242_ (.A1(_13772_),
    .A2(net2181),
    .B(_06864_),
    .Y(_06865_));
 OA21x2_ASAP7_75t_R _25243_ (.A1(_00284_),
    .A2(_16617_),
    .B(_06865_),
    .Y(_06866_));
 AOI21x1_ASAP7_75t_R _25244_ (.A1(_14002_),
    .A2(_16571_),
    .B(_06866_),
    .Y(_06867_));
 OA21x2_ASAP7_75t_R _25245_ (.A1(_13620_),
    .A2(_16571_),
    .B(_06867_),
    .Y(_16751_));
 OR3x1_ASAP7_75t_R _25246_ (.A(_01011_),
    .B(net309),
    .C(_13815_),
    .Y(_06868_));
 OAI21x1_ASAP7_75t_R _25247_ (.A1(_13817_),
    .A2(_18435_),
    .B(_06868_),
    .Y(_17793_));
 OR3x1_ASAP7_75t_R _25248_ (.A(_01077_),
    .B(net309),
    .C(_13815_),
    .Y(_06869_));
 OAI21x1_ASAP7_75t_R _25249_ (.A1(_13817_),
    .A2(_18444_),
    .B(_06869_),
    .Y(_17797_));
 NOR2x1_ASAP7_75t_R _25250_ (.A(_00284_),
    .B(_04854_),
    .Y(_06870_));
 AO221x1_ASAP7_75t_R _25251_ (.A1(_13775_),
    .A2(_01110_),
    .B1(_02208_),
    .B2(_13778_),
    .C(_13772_),
    .Y(_06871_));
 OA22x2_ASAP7_75t_R _25252_ (.A1(_13986_),
    .A2(_04808_),
    .B1(_06870_),
    .B2(_06871_),
    .Y(_06872_));
 OAI22x1_ASAP7_75t_R _25253_ (.A1(_13620_),
    .A2(_04810_),
    .B1(_06872_),
    .B2(net309),
    .Y(_06873_));
 AOI21x1_ASAP7_75t_R _25254_ (.A1(_14002_),
    .A2(_04810_),
    .B(_06873_),
    .Y(_16757_));
 OR3x1_ASAP7_75t_R _25255_ (.A(_01142_),
    .B(net309),
    .C(_13815_),
    .Y(_06874_));
 OAI21x1_ASAP7_75t_R _25256_ (.A1(_13817_),
    .A2(_18455_),
    .B(_06874_),
    .Y(_17799_));
 OR3x1_ASAP7_75t_R _25257_ (.A(_01176_),
    .B(net309),
    .C(_13815_),
    .Y(_06875_));
 OAI21x1_ASAP7_75t_R _25258_ (.A1(_13817_),
    .A2(_18460_),
    .B(_06875_),
    .Y(_16760_));
 OA21x2_ASAP7_75t_R _25259_ (.A1(_16752_),
    .A2(_05523_),
    .B(_05522_),
    .Y(_06876_));
 INVx1_ASAP7_75t_R _25260_ (.A(_06876_),
    .Y(_16759_));
 OR3x1_ASAP7_75t_R _25261_ (.A(_01208_),
    .B(net309),
    .C(_13815_),
    .Y(_06877_));
 OAI21x1_ASAP7_75t_R _25262_ (.A1(_13817_),
    .A2(_05184_),
    .B(_06877_),
    .Y(_17801_));
 OR3x1_ASAP7_75t_R _25263_ (.A(_01242_),
    .B(net309),
    .C(_13815_),
    .Y(_06878_));
 OAI21x1_ASAP7_75t_R _25264_ (.A1(_13817_),
    .A2(_18469_),
    .B(_06878_),
    .Y(_16762_));
 OA21x2_ASAP7_75t_R _25265_ (.A1(_01177_),
    .A2(_06876_),
    .B(_01210_),
    .Y(_06879_));
 OAI21x1_ASAP7_75t_R _25266_ (.A1(_01209_),
    .A2(_06879_),
    .B(_02281_),
    .Y(_16763_));
 OR3x1_ASAP7_75t_R _25267_ (.A(_01274_),
    .B(net309),
    .C(_13815_),
    .Y(_06880_));
 OAI21x1_ASAP7_75t_R _25268_ (.A1(_13817_),
    .A2(_18474_),
    .B(_06880_),
    .Y(_17803_));
 TAPCELL_ASAP7_75t_R TAP_849 ();
 TAPCELL_ASAP7_75t_R TAP_848 ();
 AND2x2_ASAP7_75t_R _25271_ (.A(_05821_),
    .B(_05840_),
    .Y(_17830_));
 AND2x2_ASAP7_75t_R _25272_ (.A(net2370),
    .B(_05840_),
    .Y(_17857_));
 INVx1_ASAP7_75t_R _25273_ (.A(_01395_),
    .Y(_16800_));
 INVx1_ASAP7_75t_R _25274_ (.A(_05975_),
    .Y(_16823_));
 OA21x2_ASAP7_75t_R _25275_ (.A1(_01398_),
    .A2(_05975_),
    .B(_01411_),
    .Y(_06882_));
 OAI21x1_ASAP7_75t_R _25276_ (.A1(net2334),
    .A2(_06882_),
    .B(_02322_),
    .Y(_16871_));
 AND2x2_ASAP7_75t_R _25277_ (.A(_05840_),
    .B(_05883_),
    .Y(_17913_));
 AOI21x1_ASAP7_75t_R _25278_ (.A1(_02326_),
    .A2(_05979_),
    .B(_05977_),
    .Y(_16925_));
 INVx1_ASAP7_75t_R _25279_ (.A(_01433_),
    .Y(_17927_));
 INVx1_ASAP7_75t_R _25280_ (.A(_01439_),
    .Y(_17947_));
 AND2x2_ASAP7_75t_R _25281_ (.A(_05840_),
    .B(_05908_),
    .Y(_17961_));
 OA21x2_ASAP7_75t_R _25282_ (.A1(_00009_),
    .A2(_05982_),
    .B(_00016_),
    .Y(_06883_));
 OAI21x1_ASAP7_75t_R _25283_ (.A1(net2145),
    .A2(_06883_),
    .B(_02336_),
    .Y(_17075_));
 INVx1_ASAP7_75t_R _25284_ (.A(_00026_),
    .Y(_17128_));
 INVx1_ASAP7_75t_R _25285_ (.A(_00028_),
    .Y(_17167_));
 OR3x1_ASAP7_75t_R _25286_ (.A(_00031_),
    .B(_05987_),
    .C(_05989_),
    .Y(_06884_));
 NAND2x1_ASAP7_75t_R _25287_ (.A(_02344_),
    .B(_06884_),
    .Y(_17276_));
 NAND2x1_ASAP7_75t_R _25288_ (.A(_02347_),
    .B(_05993_),
    .Y(_17364_));
 INVx1_ASAP7_75t_R _25289_ (.A(_17445_),
    .Y(_17395_));
 INVx1_ASAP7_75t_R _25290_ (.A(_00047_),
    .Y(_17404_));
 INVx1_ASAP7_75t_R _25291_ (.A(_05997_),
    .Y(_17455_));
 INVx1_ASAP7_75t_R _25292_ (.A(_00050_),
    .Y(_17443_));
 OA21x2_ASAP7_75t_R _25293_ (.A1(_00049_),
    .A2(_05997_),
    .B(_00053_),
    .Y(_06885_));
 OAI21x1_ASAP7_75t_R _25294_ (.A1(net2134),
    .A2(_06885_),
    .B(_02353_),
    .Y(_17533_));
 AO21x1_ASAP7_75t_R _25295_ (.A1(_00056_),
    .A2(_06001_),
    .B(_00055_),
    .Y(_06886_));
 NAND2x1_ASAP7_75t_R _25296_ (.A(_02354_),
    .B(_06886_),
    .Y(_17599_));
 INVx1_ASAP7_75t_R _25297_ (.A(_06005_),
    .Y(_17657_));
 INVx2_ASAP7_75t_R _25298_ (.A(_06007_),
    .Y(_17709_));
 INVx1_ASAP7_75t_R _25299_ (.A(_17718_),
    .Y(_17687_));
 INVx1_ASAP7_75t_R _25300_ (.A(_17725_),
    .Y(_17695_));
 INVx1_ASAP7_75t_R _25301_ (.A(_18379_),
    .Y(_18381_));
 INVx1_ASAP7_75t_R _25302_ (.A(_18389_),
    .Y(_18391_));
 INVx1_ASAP7_75t_R _25303_ (.A(_18394_),
    .Y(_18396_));
 INVx2_ASAP7_75t_R _25304_ (.A(_16262_),
    .Y(_18416_));
 INVx1_ASAP7_75t_R _25305_ (.A(_18419_),
    .Y(_18421_));
 INVx1_ASAP7_75t_R _25306_ (.A(_18424_),
    .Y(_18426_));
 INVx1_ASAP7_75t_R _25307_ (.A(_18434_),
    .Y(_18436_));
 INVx1_ASAP7_75t_R _25308_ (.A(_18439_),
    .Y(_18441_));
 INVx2_ASAP7_75t_R _25309_ (.A(_18444_),
    .Y(_18446_));
 INVx1_ASAP7_75t_R _25310_ (.A(_04919_),
    .Y(_18456_));
 INVx1_ASAP7_75t_R _25311_ (.A(_05184_),
    .Y(_18466_));
 INVx1_ASAP7_75t_R _25312_ (.A(_18474_),
    .Y(_18476_));
 INVx1_ASAP7_75t_R _25313_ (.A(_01718_),
    .Y(_06887_));
 AO32x1_ASAP7_75t_R _25314_ (.A1(net3131),
    .A2(_06235_),
    .A3(net3132),
    .B1(_06301_),
    .B2(_06887_),
    .Y(_02647_));
 OA21x2_ASAP7_75t_R _25315_ (.A1(_02032_),
    .A2(_06208_),
    .B(_06209_),
    .Y(_06888_));
 OR2x2_ASAP7_75t_R _25316_ (.A(_05744_),
    .B(_06216_),
    .Y(_06889_));
 OR3x1_ASAP7_75t_R _25317_ (.A(_14803_),
    .B(_06888_),
    .C(_06889_),
    .Y(_06890_));
 NAND2x1_ASAP7_75t_R _25318_ (.A(net3104),
    .B(_06890_),
    .Y(_06891_));
 OA211x2_ASAP7_75t_R _25319_ (.A1(_06609_),
    .A2(_06318_),
    .B(_06891_),
    .C(_05557_),
    .Y(_06892_));
 INVx1_ASAP7_75t_R _25320_ (.A(_06671_),
    .Y(_06893_));
 AND3x1_ASAP7_75t_R _25321_ (.A(_01716_),
    .B(_01717_),
    .C(_06893_),
    .Y(_06894_));
 AO21x1_ASAP7_75t_R _25322_ (.A1(_14793_),
    .A2(_06234_),
    .B(_06894_),
    .Y(_06895_));
 AO21x1_ASAP7_75t_R _25323_ (.A1(_06225_),
    .A2(_01716_),
    .B(_06562_),
    .Y(_06896_));
 AND3x1_ASAP7_75t_R _25324_ (.A(_14791_),
    .B(_06664_),
    .C(net3303),
    .Y(_06897_));
 AO221x1_ASAP7_75t_R _25325_ (.A1(_01714_),
    .A2(_06895_),
    .B1(_06896_),
    .B2(_01715_),
    .C(net3304),
    .Y(_06898_));
 NAND2x1_ASAP7_75t_R _25326_ (.A(_06655_),
    .B(net3104),
    .Y(_06899_));
 OA21x2_ASAP7_75t_R _25327_ (.A1(_05557_),
    .A2(_05748_),
    .B(_06616_),
    .Y(_06900_));
 AND3x1_ASAP7_75t_R _25328_ (.A(_14796_),
    .B(_06899_),
    .C(_06900_),
    .Y(_06901_));
 NAND2x1_ASAP7_75t_R _25329_ (.A(_01717_),
    .B(_14794_),
    .Y(_06902_));
 OA33x2_ASAP7_75t_R _25330_ (.A1(_06892_),
    .A2(_06898_),
    .A3(_06901_),
    .B1(_06902_),
    .B2(_06668_),
    .B3(net3134),
    .Y(_02648_));
 AND2x2_ASAP7_75t_R _25331_ (.A(net3132),
    .B(net3358),
    .Y(_06903_));
 AO21x1_ASAP7_75t_R _25332_ (.A1(_06655_),
    .A2(_06903_),
    .B(_05556_),
    .Y(_06904_));
 OAI21x1_ASAP7_75t_R _25333_ (.A1(_05557_),
    .A2(_05748_),
    .B(_06616_),
    .Y(_06905_));
 AO21x1_ASAP7_75t_R _25334_ (.A1(_06899_),
    .A2(_06904_),
    .B(_06905_),
    .Y(_06906_));
 AND2x2_ASAP7_75t_R _25335_ (.A(_06339_),
    .B(_06891_),
    .Y(_06907_));
 INVx1_ASAP7_75t_R _25336_ (.A(_06903_),
    .Y(_06908_));
 OAI21x1_ASAP7_75t_R _25337_ (.A1(_06615_),
    .A2(_06908_),
    .B(_06609_),
    .Y(_06909_));
 AND3x1_ASAP7_75t_R _25338_ (.A(_14793_),
    .B(_01716_),
    .C(_06893_),
    .Y(_06910_));
 AO32x1_ASAP7_75t_R _25339_ (.A1(net3132),
    .A2(net3358),
    .A3(_06910_),
    .B1(_05556_),
    .B2(_01715_),
    .Y(_06911_));
 AO21x1_ASAP7_75t_R _25340_ (.A1(_06562_),
    .A2(_06911_),
    .B(net3304),
    .Y(_06912_));
 AO221x1_ASAP7_75t_R _25341_ (.A1(_14796_),
    .A2(_06906_),
    .B1(_06907_),
    .B2(_06909_),
    .C(net3305),
    .Y(_02649_));
 AO21x1_ASAP7_75t_R _25342_ (.A1(_01717_),
    .A2(_06910_),
    .B(_06234_),
    .Y(_06913_));
 AND2x2_ASAP7_75t_R _25343_ (.A(_01714_),
    .B(_14791_),
    .Y(_06914_));
 AO21x1_ASAP7_75t_R _25344_ (.A1(_06225_),
    .A2(_01716_),
    .B(_06914_),
    .Y(_06915_));
 AO222x2_ASAP7_75t_R _25345_ (.A1(_01714_),
    .A2(_06913_),
    .B1(_06915_),
    .B2(_01715_),
    .C1(_06217_),
    .C2(_06892_),
    .Y(_06916_));
 OA21x2_ASAP7_75t_R _25346_ (.A1(_06899_),
    .A2(_06905_),
    .B(_14796_),
    .Y(_06917_));
 INVx1_ASAP7_75t_R _25347_ (.A(net3304),
    .Y(_06918_));
 OA21x2_ASAP7_75t_R _25348_ (.A1(_06916_),
    .A2(_06917_),
    .B(_06918_),
    .Y(_02650_));
 AND3x1_ASAP7_75t_R _25349_ (.A(_14794_),
    .B(_06655_),
    .C(net3104),
    .Y(_06919_));
 NAND2x1_ASAP7_75t_R _25350_ (.A(_06217_),
    .B(_06891_),
    .Y(_06920_));
 AO32x1_ASAP7_75t_R _25351_ (.A1(_01717_),
    .A2(_14794_),
    .A3(net3104),
    .B1(_06920_),
    .B2(_05557_),
    .Y(_06921_));
 AO21x1_ASAP7_75t_R _25352_ (.A1(_06900_),
    .A2(_06919_),
    .B(_06921_),
    .Y(_02651_));
 OR3x1_ASAP7_75t_R _25353_ (.A(_14828_),
    .B(_06202_),
    .C(_06692_),
    .Y(_06922_));
 AO21x1_ASAP7_75t_R _25354_ (.A1(_14828_),
    .A2(net3056),
    .B(_06621_),
    .Y(_06923_));
 AO21x1_ASAP7_75t_R _25355_ (.A1(_01713_),
    .A2(_06922_),
    .B(_06923_),
    .Y(_06924_));
 INVx1_ASAP7_75t_R _25356_ (.A(_06621_),
    .Y(_06925_));
 AOI21x1_ASAP7_75t_R _25357_ (.A1(_14797_),
    .A2(_06925_),
    .B(_01713_),
    .Y(_06926_));
 AO21x1_ASAP7_75t_R _25358_ (.A1(_05752_),
    .A2(_06924_),
    .B(_06926_),
    .Y(_02652_));
 OR3x4_ASAP7_75t_R _25359_ (.A(_01714_),
    .B(_14791_),
    .C(_06227_),
    .Y(_06927_));
 INVx1_ASAP7_75t_R _25360_ (.A(_06927_),
    .Y(_06928_));
 TAPCELL_ASAP7_75t_R TAP_847 ();
 OR3x1_ASAP7_75t_R _25362_ (.A(_05724_),
    .B(_01717_),
    .C(_06888_),
    .Y(_06930_));
 OAI21x1_ASAP7_75t_R _25363_ (.A1(_14791_),
    .A2(_06229_),
    .B(_06930_),
    .Y(_06931_));
 NAND2x2_ASAP7_75t_R _25364_ (.A(_06230_),
    .B(_06931_),
    .Y(_06932_));
 TAPCELL_ASAP7_75t_R TAP_846 ();
 AOI22x1_ASAP7_75t_R _25366_ (.A1(_06669_),
    .A2(_06928_),
    .B1(_06932_),
    .B2(_01712_),
    .Y(_02653_));
 INVx1_ASAP7_75t_R _25367_ (.A(_01711_),
    .Y(_06934_));
 AO32x1_ASAP7_75t_R _25368_ (.A1(net3102),
    .A2(_02034_),
    .A3(_06928_),
    .B1(_06932_),
    .B2(_06934_),
    .Y(_02654_));
 AND2x4_ASAP7_75t_R _25369_ (.A(_06230_),
    .B(_06931_),
    .Y(_06935_));
 OAI22x1_ASAP7_75t_R _25370_ (.A1(_02034_),
    .A2(_06927_),
    .B1(_06935_),
    .B2(_01726_),
    .Y(_02655_));
 NAND2x2_ASAP7_75t_R _25371_ (.A(_00187_),
    .B(_00191_),
    .Y(_06936_));
 AO21x2_ASAP7_75t_R _25372_ (.A1(_13495_),
    .A2(_14236_),
    .B(_05563_),
    .Y(_06937_));
 OR4x2_ASAP7_75t_R _25373_ (.A(_13525_),
    .B(net305),
    .C(_14179_),
    .D(_06937_),
    .Y(_06938_));
 AND3x1_ASAP7_75t_R _25374_ (.A(_14359_),
    .B(_05568_),
    .C(_05616_),
    .Y(_06939_));
 OA21x2_ASAP7_75t_R _25375_ (.A1(_14297_),
    .A2(_06938_),
    .B(_06939_),
    .Y(_06940_));
 AND3x2_ASAP7_75t_R _25376_ (.A(_14424_),
    .B(_14709_),
    .C(_05573_),
    .Y(_06941_));
 AND4x2_ASAP7_75t_R _25377_ (.A(_13523_),
    .B(net305),
    .C(_14179_),
    .D(_05564_),
    .Y(_06942_));
 AO31x2_ASAP7_75t_R _25378_ (.A1(_14296_),
    .A2(_14359_),
    .A3(_18360_),
    .B(_05563_),
    .Y(_06943_));
 AND3x1_ASAP7_75t_R _25379_ (.A(_06941_),
    .B(_06942_),
    .C(_06943_),
    .Y(_06944_));
 AND5x2_ASAP7_75t_R _25380_ (.A(_13523_),
    .B(net305),
    .C(_14179_),
    .D(_18380_),
    .E(_05564_),
    .Y(_06945_));
 AND4x2_ASAP7_75t_R _25381_ (.A(_14297_),
    .B(_14359_),
    .C(net310),
    .D(_05596_),
    .Y(_06946_));
 AND3x4_ASAP7_75t_R _25382_ (.A(_05586_),
    .B(_06945_),
    .C(_06946_),
    .Y(_06947_));
 TAPCELL_ASAP7_75t_R TAP_845 ();
 AO31x2_ASAP7_75t_R _25384_ (.A1(net302),
    .A2(_14359_),
    .A3(_05596_),
    .B(_05563_),
    .Y(_06949_));
 AO32x2_ASAP7_75t_R _25385_ (.A1(_05616_),
    .A2(_06938_),
    .A3(_06949_),
    .B1(_06946_),
    .B2(_05656_),
    .Y(_06950_));
 OR4x2_ASAP7_75t_R _25386_ (.A(_06940_),
    .B(_06944_),
    .C(_06947_),
    .D(_06950_),
    .Y(_06951_));
 OR3x2_ASAP7_75t_R _25387_ (.A(_05659_),
    .B(_13513_),
    .C(_13512_),
    .Y(_06952_));
 OA21x2_ASAP7_75t_R _25388_ (.A1(net2362),
    .A2(_13520_),
    .B(_14173_),
    .Y(_06953_));
 AND3x4_ASAP7_75t_R _25389_ (.A(_06952_),
    .B(_06953_),
    .C(_05564_),
    .Y(_06954_));
 AO31x2_ASAP7_75t_R _25390_ (.A1(_13523_),
    .A2(_13894_),
    .A3(_06954_),
    .B(_14358_),
    .Y(_06955_));
 AND4x2_ASAP7_75t_R _25391_ (.A(_13531_),
    .B(_14424_),
    .C(_14709_),
    .D(_05573_),
    .Y(_06956_));
 AND2x2_ASAP7_75t_R _25392_ (.A(_14296_),
    .B(_06956_),
    .Y(_06957_));
 OA211x2_ASAP7_75t_R _25393_ (.A1(_14359_),
    .A2(_05693_),
    .B(_06955_),
    .C(_06957_),
    .Y(_06958_));
 AND5x1_ASAP7_75t_R _25394_ (.A(_13523_),
    .B(_13894_),
    .C(_14179_),
    .D(_14238_),
    .E(_05570_),
    .Y(_06959_));
 AO21x2_ASAP7_75t_R _25395_ (.A1(net302),
    .A2(_14359_),
    .B(_05563_),
    .Y(_06960_));
 OA211x2_ASAP7_75t_R _25396_ (.A1(_05693_),
    .A2(_06959_),
    .B(_06960_),
    .C(_06956_),
    .Y(_06961_));
 OR3x1_ASAP7_75t_R _25397_ (.A(_14179_),
    .B(_14239_),
    .C(_14297_),
    .Y(_06962_));
 OA211x2_ASAP7_75t_R _25398_ (.A1(_05667_),
    .A2(_06962_),
    .B(_06956_),
    .C(_14358_),
    .Y(_06963_));
 AND5x2_ASAP7_75t_R _25399_ (.A(_05626_),
    .B(_14424_),
    .C(_14709_),
    .D(_05570_),
    .E(_05572_),
    .Y(_06964_));
 AND3x4_ASAP7_75t_R _25400_ (.A(_01743_),
    .B(_05630_),
    .C(_06964_),
    .Y(_06965_));
 TAPCELL_ASAP7_75t_R TAP_844 ();
 AND4x1_ASAP7_75t_R _25402_ (.A(_05724_),
    .B(_05568_),
    .C(_05584_),
    .D(_05588_),
    .Y(_06967_));
 AO21x2_ASAP7_75t_R _25403_ (.A1(_14180_),
    .A2(_14238_),
    .B(_05563_),
    .Y(_06968_));
 OA21x2_ASAP7_75t_R _25404_ (.A1(_06965_),
    .A2(_06967_),
    .B(_06968_),
    .Y(_06969_));
 AND2x2_ASAP7_75t_R _25405_ (.A(_05626_),
    .B(_05570_),
    .Y(_06970_));
 OAI21x1_ASAP7_75t_R _25406_ (.A1(_14179_),
    .A2(_14239_),
    .B(_06970_),
    .Y(_06971_));
 OA211x2_ASAP7_75t_R _25407_ (.A1(_13521_),
    .A2(_14703_),
    .B(_05568_),
    .C(_14358_),
    .Y(_06972_));
 NAND2x1_ASAP7_75t_R _25408_ (.A(_14357_),
    .B(_05570_),
    .Y(_06973_));
 AND4x1_ASAP7_75t_R _25409_ (.A(_14296_),
    .B(_06973_),
    .C(_05588_),
    .D(_05678_),
    .Y(_06974_));
 AO32x1_ASAP7_75t_R _25410_ (.A1(_06941_),
    .A2(_06971_),
    .A3(_06972_),
    .B1(_06974_),
    .B2(_05663_),
    .Y(_06975_));
 OR5x2_ASAP7_75t_R _25411_ (.A(_06958_),
    .B(_06961_),
    .C(_06963_),
    .D(_06969_),
    .E(_06975_),
    .Y(_06976_));
 OAI21x1_ASAP7_75t_R _25412_ (.A1(_06951_),
    .A2(_06976_),
    .B(_05739_),
    .Y(_06977_));
 AO221x1_ASAP7_75t_R _25413_ (.A1(_00172_),
    .A2(_13492_),
    .B1(_13802_),
    .B2(_13803_),
    .C(_13552_),
    .Y(_06978_));
 AND3x4_ASAP7_75t_R _25414_ (.A(_05752_),
    .B(_06925_),
    .C(_06978_),
    .Y(_06979_));
 INVx1_ASAP7_75t_R _25415_ (.A(_06979_),
    .Y(_06980_));
 AOI21x1_ASAP7_75t_R _25416_ (.A1(net310),
    .A2(_06977_),
    .B(_06980_),
    .Y(_06981_));
 TAPCELL_ASAP7_75t_R TAP_843 ();
 AND5x1_ASAP7_75t_R _25418_ (.A(net2804),
    .B(_05551_),
    .C(_01316_),
    .D(_01607_),
    .E(_05552_),
    .Y(_06983_));
 OAI21x1_ASAP7_75t_R _25419_ (.A1(_06981_),
    .A2(_06983_),
    .B(_13890_),
    .Y(_06984_));
 OR3x4_ASAP7_75t_R _25420_ (.A(_05658_),
    .B(_14293_),
    .C(_06984_),
    .Y(_06985_));
 TAPCELL_ASAP7_75t_R TAP_842 ();
 NOR2x2_ASAP7_75t_R _25422_ (.A(_06936_),
    .B(_06985_),
    .Y(_06987_));
 TAPCELL_ASAP7_75t_R TAP_841 ();
 TAPCELL_ASAP7_75t_R TAP_840 ();
 NAND3x2_ASAP7_75t_R _25425_ (.B(_05630_),
    .C(_06964_),
    .Y(_06990_),
    .A(_01743_));
 TAPCELL_ASAP7_75t_R TAP_839 ();
 OA31x2_ASAP7_75t_R _25427_ (.A1(_14179_),
    .A2(_14239_),
    .A3(_05662_),
    .B1(net310),
    .Y(_06992_));
 TAPCELL_ASAP7_75t_R TAP_838 ();
 OR4x2_ASAP7_75t_R _25429_ (.A(_13523_),
    .B(_13894_),
    .C(_14179_),
    .D(_06937_),
    .Y(_06994_));
 TAPCELL_ASAP7_75t_R TAP_837 ();
 OA22x2_ASAP7_75t_R _25431_ (.A1(_02139_),
    .A2(_06992_),
    .B1(_06994_),
    .B2(_01913_),
    .Y(_06996_));
 NAND2x1_ASAP7_75t_R _25432_ (.A(_13523_),
    .B(_13894_),
    .Y(_06997_));
 OR4x2_ASAP7_75t_R _25433_ (.A(_14179_),
    .B(_06937_),
    .C(_06997_),
    .D(_06990_),
    .Y(_06998_));
 TAPCELL_ASAP7_75t_R TAP_836 ();
 OR2x6_ASAP7_75t_R _25435_ (.A(_05589_),
    .B(_06992_),
    .Y(_07000_));
 TAPCELL_ASAP7_75t_R TAP_835 ();
 OA22x2_ASAP7_75t_R _25437_ (.A1(_01945_),
    .A2(_06998_),
    .B1(_07000_),
    .B2(_01577_),
    .Y(_07002_));
 OR4x2_ASAP7_75t_R _25438_ (.A(_05594_),
    .B(_05622_),
    .C(_05598_),
    .D(_05600_),
    .Y(_07003_));
 OR4x2_ASAP7_75t_R _25439_ (.A(_14297_),
    .B(_14359_),
    .C(_06992_),
    .D(_07003_),
    .Y(_07004_));
 TAPCELL_ASAP7_75t_R TAP_834 ();
 OA21x2_ASAP7_75t_R _25441_ (.A1(_14297_),
    .A2(_14358_),
    .B(net310),
    .Y(_07006_));
 OR4x1_ASAP7_75t_R _25442_ (.A(_13525_),
    .B(net305),
    .C(_14180_),
    .D(_06937_),
    .Y(_07007_));
 OR3x4_ASAP7_75t_R _25443_ (.A(_07003_),
    .B(_07006_),
    .C(_07007_),
    .Y(_07008_));
 OA21x2_ASAP7_75t_R _25444_ (.A1(_00661_),
    .A2(_07004_),
    .B(_07008_),
    .Y(_07009_));
 OA211x2_ASAP7_75t_R _25445_ (.A1(_06990_),
    .A2(_06996_),
    .B(_07002_),
    .C(_07009_),
    .Y(_07010_));
 TAPCELL_ASAP7_75t_R TAP_833 ();
 NAND2x1_ASAP7_75t_R _25447_ (.A(net3516),
    .B(_06947_),
    .Y(_07012_));
 OR4x1_ASAP7_75t_R _25448_ (.A(_14179_),
    .B(_14239_),
    .C(_14297_),
    .D(_05662_),
    .Y(_07013_));
 AND2x6_ASAP7_75t_R _25449_ (.A(net310),
    .B(_07013_),
    .Y(_07014_));
 TAPCELL_ASAP7_75t_R TAP_832 ();
 OR2x6_ASAP7_75t_R _25451_ (.A(_14297_),
    .B(_06994_),
    .Y(_07016_));
 TAPCELL_ASAP7_75t_R TAP_831 ();
 TAPCELL_ASAP7_75t_R TAP_830 ();
 OAI22x1_ASAP7_75t_R _25454_ (.A1(_00659_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_00660_),
    .Y(_07019_));
 NAND2x1_ASAP7_75t_R _25455_ (.A(_06950_),
    .B(_07019_),
    .Y(_07020_));
 OAI21x1_ASAP7_75t_R _25456_ (.A1(_14297_),
    .A2(_06938_),
    .B(_06939_),
    .Y(_07021_));
 OA22x2_ASAP7_75t_R _25457_ (.A1(_02172_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02066_),
    .Y(_07022_));
 OR4x2_ASAP7_75t_R _25458_ (.A(_13523_),
    .B(net305),
    .C(_14179_),
    .D(_06937_),
    .Y(_07023_));
 OR2x6_ASAP7_75t_R _25459_ (.A(_05589_),
    .B(_07023_),
    .Y(_07024_));
 TAPCELL_ASAP7_75t_R TAP_829 ();
 OR2x6_ASAP7_75t_R _25461_ (.A(_05589_),
    .B(_06994_),
    .Y(_07026_));
 TAPCELL_ASAP7_75t_R TAP_828 ();
 OR2x6_ASAP7_75t_R _25463_ (.A(_06990_),
    .B(_07023_),
    .Y(_07028_));
 TAPCELL_ASAP7_75t_R TAP_827 ();
 OA222x2_ASAP7_75t_R _25465_ (.A1(_01995_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02098_),
    .C1(_07028_),
    .C2(_02029_),
    .Y(_07030_));
 OA21x2_ASAP7_75t_R _25466_ (.A1(_07021_),
    .A2(_07022_),
    .B(_07030_),
    .Y(_07031_));
 AND4x2_ASAP7_75t_R _25467_ (.A(_07010_),
    .B(_07012_),
    .C(_07020_),
    .D(_07031_),
    .Y(_07032_));
 AND4x1_ASAP7_75t_R _25468_ (.A(_13802_),
    .B(_13803_),
    .C(_06981_),
    .D(_07032_),
    .Y(_07033_));
 NAND2x2_ASAP7_75t_R _25469_ (.A(_01730_),
    .B(_01731_),
    .Y(_07034_));
 INVx1_ASAP7_75t_R _25470_ (.A(_01863_),
    .Y(_07035_));
 AND2x6_ASAP7_75t_R _25471_ (.A(_01730_),
    .B(_01731_),
    .Y(_07036_));
 AND2x2_ASAP7_75t_R _25472_ (.A(_07035_),
    .B(_07036_),
    .Y(_07037_));
 AO21x1_ASAP7_75t_R _25473_ (.A1(net34),
    .A2(_07034_),
    .B(_07037_),
    .Y(_07038_));
 CKINVDCx8_ASAP7_75t_R _25474_ (.A(_01642_),
    .Y(_07039_));
 TAPCELL_ASAP7_75t_R TAP_826 ();
 AND2x6_ASAP7_75t_R _25476_ (.A(_07039_),
    .B(net433),
    .Y(_07041_));
 TAPCELL_ASAP7_75t_R TAP_825 ();
 TAPCELL_ASAP7_75t_R TAP_824 ();
 NOR2x2_ASAP7_75t_R _25479_ (.A(net432),
    .B(net433),
    .Y(_07044_));
 INVx1_ASAP7_75t_R _25480_ (.A(net2392),
    .Y(_07045_));
 AND2x6_ASAP7_75t_R _25481_ (.A(_05762_),
    .B(_01731_),
    .Y(_07046_));
 TAPCELL_ASAP7_75t_R TAP_823 ();
 OAI22x1_ASAP7_75t_R _25483_ (.A1(_07045_),
    .A2(_01730_),
    .B1(_01855_),
    .B2(_07046_),
    .Y(_07048_));
 AND2x2_ASAP7_75t_R _25484_ (.A(net27),
    .B(net433),
    .Y(_07049_));
 NAND2x1_ASAP7_75t_R _25485_ (.A(_01871_),
    .B(_07036_),
    .Y(_07050_));
 CKINVDCx8_ASAP7_75t_R _25486_ (.A(_01643_),
    .Y(_07051_));
 OA211x2_ASAP7_75t_R _25487_ (.A1(net57),
    .A2(_07036_),
    .B(_07050_),
    .C(_07051_),
    .Y(_07052_));
 TAPCELL_ASAP7_75t_R TAP_822 ();
 OA21x2_ASAP7_75t_R _25489_ (.A1(_07049_),
    .A2(_07052_),
    .B(net432),
    .Y(_07054_));
 AO221x2_ASAP7_75t_R _25490_ (.A1(_07038_),
    .A2(_07041_),
    .B1(_07044_),
    .B2(_07048_),
    .C(_07054_),
    .Y(_07055_));
 NOR2x2_ASAP7_75t_R _25491_ (.A(net290),
    .B(_07055_),
    .Y(_07056_));
 TAPCELL_ASAP7_75t_R TAP_821 ();
 TAPCELL_ASAP7_75t_R TAP_820 ();
 AND2x6_ASAP7_75t_R _25494_ (.A(_13570_),
    .B(_13534_),
    .Y(_07059_));
 NAND2x2_ASAP7_75t_R _25495_ (.A(_13537_),
    .B(_07059_),
    .Y(_07060_));
 NAND2x2_ASAP7_75t_R _25496_ (.A(_01314_),
    .B(_01732_),
    .Y(_07061_));
 OR2x6_ASAP7_75t_R _25497_ (.A(_05815_),
    .B(_07061_),
    .Y(_07062_));
 TAPCELL_ASAP7_75t_R TAP_819 ();
 NOR2x2_ASAP7_75t_R _25499_ (.A(_05815_),
    .B(_07061_),
    .Y(_07064_));
 OR2x6_ASAP7_75t_R _25500_ (.A(_07059_),
    .B(_07064_),
    .Y(_07065_));
 TAPCELL_ASAP7_75t_R TAP_818 ();
 AO32x2_ASAP7_75t_R _25502_ (.A1(_01356_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00324_),
    .Y(_07067_));
 AND3x1_ASAP7_75t_R _25503_ (.A(_13817_),
    .B(_06979_),
    .C(_07067_),
    .Y(_07068_));
 TAPCELL_ASAP7_75t_R TAP_817 ();
 TAPCELL_ASAP7_75t_R TAP_816 ();
 NAND2x2_ASAP7_75t_R _25506_ (.A(_01713_),
    .B(_13459_),
    .Y(_07071_));
 OA31x2_ASAP7_75t_R _25507_ (.A1(_02357_),
    .A2(_14179_),
    .A3(_14239_),
    .B1(_07071_),
    .Y(_07072_));
 XNOR2x2_ASAP7_75t_R _25508_ (.A(net302),
    .B(_07072_),
    .Y(_07073_));
 TAPCELL_ASAP7_75t_R TAP_815 ();
 NAND2x1_ASAP7_75t_R _25510_ (.A(_13548_),
    .B(_13553_),
    .Y(_07075_));
 OR3x1_ASAP7_75t_R _25511_ (.A(_13564_),
    .B(_13569_),
    .C(_13575_),
    .Y(_07076_));
 OA211x2_ASAP7_75t_R _25512_ (.A1(_07075_),
    .A2(_07076_),
    .B(_06634_),
    .C(_06632_),
    .Y(_07077_));
 TAPCELL_ASAP7_75t_R TAP_814 ();
 TAPCELL_ASAP7_75t_R TAP_813 ();
 AO211x2_ASAP7_75t_R _25515_ (.A1(_13554_),
    .A2(_13576_),
    .B(_13606_),
    .C(_13584_),
    .Y(_07080_));
 TAPCELL_ASAP7_75t_R TAP_812 ();
 OA21x2_ASAP7_75t_R _25517_ (.A1(_01613_),
    .A2(_13807_),
    .B(_07080_),
    .Y(_07082_));
 AO32x2_ASAP7_75t_R _25518_ (.A1(_14987_),
    .A2(_14992_),
    .A3(_07077_),
    .B1(_07082_),
    .B2(_05183_),
    .Y(_07083_));
 TAPCELL_ASAP7_75t_R TAP_811 ();
 OA211x2_ASAP7_75t_R _25520_ (.A1(_01612_),
    .A2(_13807_),
    .B(_05293_),
    .C(_07080_),
    .Y(_07085_));
 AO32x2_ASAP7_75t_R _25521_ (.A1(_14854_),
    .A2(_14923_),
    .A3(_07077_),
    .B1(_07085_),
    .B2(_05292_),
    .Y(_07086_));
 AND2x2_ASAP7_75t_R _25522_ (.A(_13894_),
    .B(_07086_),
    .Y(_07087_));
 AO21x2_ASAP7_75t_R _25523_ (.A1(net304),
    .A2(_07083_),
    .B(_07087_),
    .Y(_07088_));
 NAND2x1_ASAP7_75t_R _25524_ (.A(_00073_),
    .B(_07071_),
    .Y(_07089_));
 OA21x2_ASAP7_75t_R _25525_ (.A1(_07071_),
    .A2(_14179_),
    .B(_07089_),
    .Y(_07090_));
 TAPCELL_ASAP7_75t_R TAP_810 ();
 AO21x2_ASAP7_75t_R _25527_ (.A1(_01713_),
    .A2(_13459_),
    .B(_00072_),
    .Y(_07092_));
 AO221x2_ASAP7_75t_R _25528_ (.A1(_13442_),
    .A2(_13474_),
    .B1(_13514_),
    .B2(_13522_),
    .C(_07071_),
    .Y(_07093_));
 AND2x6_ASAP7_75t_R _25529_ (.A(_07092_),
    .B(_07093_),
    .Y(_07094_));
 NAND2x2_ASAP7_75t_R _25530_ (.A(_07090_),
    .B(_07094_),
    .Y(_07095_));
 NAND2x2_ASAP7_75t_R _25531_ (.A(_07092_),
    .B(_07093_),
    .Y(_07096_));
 NAND2x2_ASAP7_75t_R _25532_ (.A(_07090_),
    .B(_07096_),
    .Y(_07097_));
 OA21x2_ASAP7_75t_R _25533_ (.A1(_13997_),
    .A2(_13998_),
    .B(_07077_),
    .Y(_07098_));
 AND3x4_ASAP7_75t_R _25534_ (.A(_05457_),
    .B(_05511_),
    .C(_07080_),
    .Y(_07099_));
 OA21x2_ASAP7_75t_R _25535_ (.A1(_07098_),
    .A2(_07099_),
    .B(_13894_),
    .Y(_07100_));
 AO211x2_ASAP7_75t_R _25536_ (.A1(_13810_),
    .A2(_05400_),
    .B(_05403_),
    .C(_07077_),
    .Y(_07101_));
 OA31x2_ASAP7_75t_R _25537_ (.A1(_13809_),
    .A2(_13814_),
    .A3(_07080_),
    .B1(_07101_),
    .Y(_07102_));
 AND2x4_ASAP7_75t_R _25538_ (.A(net303),
    .B(_07102_),
    .Y(_07103_));
 NOR2x2_ASAP7_75t_R _25539_ (.A(_07100_),
    .B(_07103_),
    .Y(_07104_));
 OA22x2_ASAP7_75t_R _25540_ (.A1(_07088_),
    .A2(_07095_),
    .B1(_07097_),
    .B2(_07104_),
    .Y(_07105_));
 TAPCELL_ASAP7_75t_R TAP_809 ();
 OR3x4_ASAP7_75t_R _25542_ (.A(_15223_),
    .B(_15225_),
    .C(_07080_),
    .Y(_07107_));
 OR3x4_ASAP7_75t_R _25543_ (.A(_04745_),
    .B(_04746_),
    .C(_07077_),
    .Y(_07108_));
 AND3x1_ASAP7_75t_R _25544_ (.A(_07094_),
    .B(_07107_),
    .C(_07108_),
    .Y(_07109_));
 TAPCELL_ASAP7_75t_R TAP_808 ();
 NAND2x1_ASAP7_75t_R _25546_ (.A(_18351_),
    .B(_07077_),
    .Y(_07111_));
 OA211x2_ASAP7_75t_R _25547_ (.A1(_04967_),
    .A2(_07077_),
    .B(_07111_),
    .C(_07096_),
    .Y(_07112_));
 OA21x2_ASAP7_75t_R _25548_ (.A1(_07109_),
    .A2(_07112_),
    .B(net304),
    .Y(_07113_));
 NAND2x1_ASAP7_75t_R _25549_ (.A(_18344_),
    .B(_07077_),
    .Y(_07114_));
 OA21x2_ASAP7_75t_R _25550_ (.A1(_05077_),
    .A2(_07077_),
    .B(_07114_),
    .Y(_07115_));
 OA211x2_ASAP7_75t_R _25551_ (.A1(_15112_),
    .A2(_04854_),
    .B(_07080_),
    .C(_04856_),
    .Y(_07116_));
 AO21x2_ASAP7_75t_R _25552_ (.A1(_15172_),
    .A2(_07077_),
    .B(_07116_),
    .Y(_07117_));
 OR2x2_ASAP7_75t_R _25553_ (.A(_07096_),
    .B(_07117_),
    .Y(_07118_));
 TAPCELL_ASAP7_75t_R TAP_807 ();
 OA211x2_ASAP7_75t_R _25555_ (.A1(_07094_),
    .A2(_07115_),
    .B(_07118_),
    .C(_13894_),
    .Y(_07120_));
 OAI21x1_ASAP7_75t_R _25556_ (.A1(_07071_),
    .A2(_14179_),
    .B(_07089_),
    .Y(_07121_));
 TAPCELL_ASAP7_75t_R TAP_806 ();
 OAI21x1_ASAP7_75t_R _25558_ (.A1(_07113_),
    .A2(_07120_),
    .B(_07121_),
    .Y(_07123_));
 AND2x2_ASAP7_75t_R _25559_ (.A(_02358_),
    .B(_07071_),
    .Y(_07124_));
 XNOR2x2_ASAP7_75t_R _25560_ (.A(_14238_),
    .B(_07124_),
    .Y(_07125_));
 AO211x2_ASAP7_75t_R _25561_ (.A1(_13810_),
    .A2(_14783_),
    .B(_14787_),
    .C(_07080_),
    .Y(_07126_));
 OA31x2_ASAP7_75t_R _25562_ (.A1(_16507_),
    .A2(_16508_),
    .A3(_07077_),
    .B1(_07126_),
    .Y(_07127_));
 OA211x2_ASAP7_75t_R _25563_ (.A1(_15112_),
    .A2(_16617_),
    .B(_07080_),
    .C(_16619_),
    .Y(_07128_));
 AO211x2_ASAP7_75t_R _25564_ (.A1(_15401_),
    .A2(_07077_),
    .B(_07128_),
    .C(net305),
    .Y(_07129_));
 OA21x2_ASAP7_75t_R _25565_ (.A1(_13894_),
    .A2(_07127_),
    .B(_07129_),
    .Y(_07130_));
 OR2x2_ASAP7_75t_R _25566_ (.A(_15280_),
    .B(_07080_),
    .Y(_07131_));
 OR3x1_ASAP7_75t_R _25567_ (.A(_04630_),
    .B(_04631_),
    .C(_07077_),
    .Y(_07132_));
 OR2x2_ASAP7_75t_R _25568_ (.A(_04516_),
    .B(_07077_),
    .Y(_07133_));
 TAPCELL_ASAP7_75t_R TAP_805 ();
 OA21x2_ASAP7_75t_R _25570_ (.A1(_15337_),
    .A2(_07080_),
    .B(net304),
    .Y(_07135_));
 AO32x2_ASAP7_75t_R _25571_ (.A1(_13894_),
    .A2(_07131_),
    .A3(_07132_),
    .B1(_07133_),
    .B2(_07135_),
    .Y(_07136_));
 OAI22x1_ASAP7_75t_R _25572_ (.A1(_07095_),
    .A2(_07130_),
    .B1(_07136_),
    .B2(_07097_),
    .Y(_07137_));
 OR2x2_ASAP7_75t_R _25573_ (.A(_15887_),
    .B(_07080_),
    .Y(_07138_));
 OA31x2_ASAP7_75t_R _25574_ (.A1(_16018_),
    .A2(_16019_),
    .A3(_07077_),
    .B1(net304),
    .Y(_07139_));
 AO211x2_ASAP7_75t_R _25575_ (.A1(_13810_),
    .A2(_15773_),
    .B(_15777_),
    .C(_07080_),
    .Y(_07140_));
 AO211x2_ASAP7_75t_R _25576_ (.A1(_13810_),
    .A2(_16138_),
    .B(_16144_),
    .C(_07077_),
    .Y(_07141_));
 AND3x1_ASAP7_75t_R _25577_ (.A(_13894_),
    .B(_07140_),
    .C(_07141_),
    .Y(_07142_));
 AOI21x1_ASAP7_75t_R _25578_ (.A1(_07138_),
    .A2(_07139_),
    .B(_07142_),
    .Y(_07143_));
 AND3x1_ASAP7_75t_R _25579_ (.A(_07121_),
    .B(_07094_),
    .C(_07143_),
    .Y(_07144_));
 TAPCELL_ASAP7_75t_R TAP_804 ();
 AND2x2_ASAP7_75t_R _25581_ (.A(_18390_),
    .B(_07077_),
    .Y(_07146_));
 AOI211x1_ASAP7_75t_R _25582_ (.A1(_16262_),
    .A2(_07080_),
    .B(_07146_),
    .C(_13894_),
    .Y(_07147_));
 AND2x2_ASAP7_75t_R _25583_ (.A(_16386_),
    .B(_07080_),
    .Y(_07148_));
 AOI211x1_ASAP7_75t_R _25584_ (.A1(_18385_),
    .A2(_07077_),
    .B(_07148_),
    .C(net303),
    .Y(_07149_));
 NAND2x2_ASAP7_75t_R _25585_ (.A(_07121_),
    .B(_07096_),
    .Y(_07150_));
 NOR3x2_ASAP7_75t_R _25586_ (.B(_07149_),
    .C(_07150_),
    .Y(_07151_),
    .A(_07147_));
 XNOR2x2_ASAP7_75t_R _25587_ (.A(_14239_),
    .B(_07124_),
    .Y(_07152_));
 OA31x2_ASAP7_75t_R _25588_ (.A1(_07137_),
    .A2(_07144_),
    .A3(_07151_),
    .B1(_07152_),
    .Y(_07153_));
 AO31x2_ASAP7_75t_R _25589_ (.A1(_07105_),
    .A2(_07123_),
    .A3(_07125_),
    .B(_07153_),
    .Y(_07154_));
 NAND2x1_ASAP7_75t_R _25590_ (.A(_18409_),
    .B(_07077_),
    .Y(_07155_));
 NAND2x1_ASAP7_75t_R _25591_ (.A(_18394_),
    .B(_07080_),
    .Y(_07156_));
 OR2x2_ASAP7_75t_R _25592_ (.A(_15887_),
    .B(_07077_),
    .Y(_07157_));
 OA31x2_ASAP7_75t_R _25593_ (.A1(_16018_),
    .A2(_16019_),
    .A3(_07080_),
    .B1(_13894_),
    .Y(_07158_));
 AO32x2_ASAP7_75t_R _25594_ (.A1(net305),
    .A2(_07155_),
    .A3(_07156_),
    .B1(_07157_),
    .B2(_07158_),
    .Y(_07159_));
 AND2x2_ASAP7_75t_R _25595_ (.A(_16386_),
    .B(_07077_),
    .Y(_07160_));
 AOI211x1_ASAP7_75t_R _25596_ (.A1(_18385_),
    .A2(_07080_),
    .B(_07160_),
    .C(_13894_),
    .Y(_07161_));
 TAPCELL_ASAP7_75t_R TAP_803 ();
 AND2x2_ASAP7_75t_R _25598_ (.A(_18390_),
    .B(_07080_),
    .Y(_07163_));
 AOI211x1_ASAP7_75t_R _25599_ (.A1(_16262_),
    .A2(_07077_),
    .B(_07163_),
    .C(net303),
    .Y(_07164_));
 OR3x1_ASAP7_75t_R _25600_ (.A(_07095_),
    .B(_07161_),
    .C(_07164_),
    .Y(_07165_));
 NAND2x2_ASAP7_75t_R _25601_ (.A(_07121_),
    .B(_07094_),
    .Y(_07166_));
 OR2x2_ASAP7_75t_R _25602_ (.A(_15280_),
    .B(_07077_),
    .Y(_07167_));
 OR3x1_ASAP7_75t_R _25603_ (.A(_04630_),
    .B(_04631_),
    .C(_07080_),
    .Y(_07168_));
 OR2x2_ASAP7_75t_R _25604_ (.A(_04516_),
    .B(_07080_),
    .Y(_07169_));
 OA21x2_ASAP7_75t_R _25605_ (.A1(_15337_),
    .A2(_07077_),
    .B(_13894_),
    .Y(_07170_));
 AO32x2_ASAP7_75t_R _25606_ (.A1(net304),
    .A2(_07167_),
    .A3(_07168_),
    .B1(_07169_),
    .B2(_07170_),
    .Y(_07171_));
 AO211x2_ASAP7_75t_R _25607_ (.A1(_13810_),
    .A2(_14783_),
    .B(_14787_),
    .C(_07077_),
    .Y(_07172_));
 OA31x2_ASAP7_75t_R _25608_ (.A1(_16507_),
    .A2(_16508_),
    .A3(_07080_),
    .B1(_07172_),
    .Y(_07173_));
 AO211x2_ASAP7_75t_R _25609_ (.A1(_13810_),
    .A2(net2310),
    .B(_15400_),
    .C(_07077_),
    .Y(_07174_));
 OA211x2_ASAP7_75t_R _25610_ (.A1(_16620_),
    .A2(_07080_),
    .B(_07174_),
    .C(net305),
    .Y(_07175_));
 AO21x1_ASAP7_75t_R _25611_ (.A1(_13894_),
    .A2(_07173_),
    .B(_07175_),
    .Y(_07176_));
 OA22x2_ASAP7_75t_R _25612_ (.A1(_07166_),
    .A2(_07171_),
    .B1(_07176_),
    .B2(_07150_),
    .Y(_07177_));
 OA211x2_ASAP7_75t_R _25613_ (.A1(_07097_),
    .A2(_07159_),
    .B(_07165_),
    .C(_07177_),
    .Y(_07178_));
 TAPCELL_ASAP7_75t_R TAP_802 ();
 TAPCELL_ASAP7_75t_R TAP_801 ();
 NAND2x1_ASAP7_75t_R _25616_ (.A(_18351_),
    .B(_07080_),
    .Y(_07181_));
 OA21x2_ASAP7_75t_R _25617_ (.A1(_04967_),
    .A2(_07080_),
    .B(_07181_),
    .Y(_07182_));
 NAND2x1_ASAP7_75t_R _25618_ (.A(_18344_),
    .B(_07080_),
    .Y(_07183_));
 OA211x2_ASAP7_75t_R _25619_ (.A1(_05077_),
    .A2(_07080_),
    .B(_07183_),
    .C(net304),
    .Y(_07184_));
 AOI21x1_ASAP7_75t_R _25620_ (.A1(_13894_),
    .A2(_07182_),
    .B(_07184_),
    .Y(_07185_));
 TAPCELL_ASAP7_75t_R TAP_800 ();
 OR3x1_ASAP7_75t_R _25622_ (.A(_04745_),
    .B(_04746_),
    .C(_07080_),
    .Y(_07187_));
 OR3x1_ASAP7_75t_R _25623_ (.A(_15223_),
    .B(_15225_),
    .C(_07077_),
    .Y(_07188_));
 AO211x2_ASAP7_75t_R _25624_ (.A1(_13810_),
    .A2(_15167_),
    .B(_15171_),
    .C(_07077_),
    .Y(_07189_));
 OA211x2_ASAP7_75t_R _25625_ (.A1(_04857_),
    .A2(_07080_),
    .B(_07189_),
    .C(net305),
    .Y(_07190_));
 AO31x2_ASAP7_75t_R _25626_ (.A1(_13894_),
    .A2(_07187_),
    .A3(_07188_),
    .B(_07190_),
    .Y(_07191_));
 NOR2x1_ASAP7_75t_R _25627_ (.A(_07094_),
    .B(_07191_),
    .Y(_07192_));
 AOI21x1_ASAP7_75t_R _25628_ (.A1(_07094_),
    .A2(_07185_),
    .B(_07192_),
    .Y(_07193_));
 TAPCELL_ASAP7_75t_R TAP_799 ();
 AND2x2_ASAP7_75t_R _25630_ (.A(_07090_),
    .B(_07152_),
    .Y(_07195_));
 AOI22x1_ASAP7_75t_R _25631_ (.A1(_07125_),
    .A2(_07178_),
    .B1(_07193_),
    .B2(_07195_),
    .Y(_07196_));
 AND2x2_ASAP7_75t_R _25632_ (.A(_07121_),
    .B(_07152_),
    .Y(_07197_));
 TAPCELL_ASAP7_75t_R TAP_798 ();
 TAPCELL_ASAP7_75t_R TAP_797 ();
 AND3x2_ASAP7_75t_R _25635_ (.A(_14854_),
    .B(_14923_),
    .C(_07080_),
    .Y(_07200_));
 AOI21x1_ASAP7_75t_R _25636_ (.A1(_18469_),
    .A2(_07077_),
    .B(_07200_),
    .Y(_07201_));
 OA21x2_ASAP7_75t_R _25637_ (.A1(_01613_),
    .A2(_13807_),
    .B(_07077_),
    .Y(_07202_));
 AOI22x1_ASAP7_75t_R _25638_ (.A1(_18339_),
    .A2(_07080_),
    .B1(_07202_),
    .B2(_05183_),
    .Y(_07203_));
 AND2x2_ASAP7_75t_R _25639_ (.A(_13894_),
    .B(_07203_),
    .Y(_07204_));
 AO21x2_ASAP7_75t_R _25640_ (.A1(_13893_),
    .A2(_07201_),
    .B(_07204_),
    .Y(_07205_));
 AND2x2_ASAP7_75t_R _25641_ (.A(_18474_),
    .B(_07077_),
    .Y(_07206_));
 AO21x1_ASAP7_75t_R _25642_ (.A1(_18332_),
    .A2(_07080_),
    .B(_07206_),
    .Y(_07207_));
 NAND2x1_ASAP7_75t_R _25643_ (.A(_17807_),
    .B(_07077_),
    .Y(_07208_));
 OA211x2_ASAP7_75t_R _25644_ (.A1(_18326_),
    .A2(_07077_),
    .B(_07208_),
    .C(_13893_),
    .Y(_07209_));
 TAPCELL_ASAP7_75t_R TAP_796 ();
 AOI211x1_ASAP7_75t_R _25646_ (.A1(_13894_),
    .A2(_07207_),
    .B(_07209_),
    .C(_07096_),
    .Y(_07211_));
 AO21x1_ASAP7_75t_R _25647_ (.A1(_07096_),
    .A2(_07205_),
    .B(_07211_),
    .Y(_07212_));
 AOI21x1_ASAP7_75t_R _25648_ (.A1(_07197_),
    .A2(_07212_),
    .B(_07073_),
    .Y(_07213_));
 AND2x2_ASAP7_75t_R _25649_ (.A(_13578_),
    .B(_13582_),
    .Y(_07214_));
 OA21x2_ASAP7_75t_R _25650_ (.A1(_06633_),
    .A2(_13606_),
    .B(_07214_),
    .Y(_07215_));
 INVx2_ASAP7_75t_R _25651_ (.A(_07215_),
    .Y(_07216_));
 AO221x2_ASAP7_75t_R _25652_ (.A1(_07073_),
    .A2(_07154_),
    .B1(_07196_),
    .B2(_07213_),
    .C(_07216_),
    .Y(_07217_));
 XNOR2x2_ASAP7_75t_R _25653_ (.A(_14297_),
    .B(_07072_),
    .Y(_07218_));
 NAND2x2_ASAP7_75t_R _25654_ (.A(_07218_),
    .B(_07152_),
    .Y(_07219_));
 AND3x4_ASAP7_75t_R _25655_ (.A(_07214_),
    .B(_06633_),
    .C(_06634_),
    .Y(_07220_));
 AND3x1_ASAP7_75t_R _25656_ (.A(net304),
    .B(_07092_),
    .C(_07093_),
    .Y(_07221_));
 OA22x2_ASAP7_75t_R _25657_ (.A1(_07098_),
    .A2(_07099_),
    .B1(_07220_),
    .B2(_07221_),
    .Y(_07222_));
 AND2x6_ASAP7_75t_R _25658_ (.A(_17807_),
    .B(_07220_),
    .Y(_07223_));
 AND2x2_ASAP7_75t_R _25659_ (.A(_07090_),
    .B(_07223_),
    .Y(_07224_));
 AO21x1_ASAP7_75t_R _25660_ (.A1(_07121_),
    .A2(_07222_),
    .B(_07224_),
    .Y(_07225_));
 TAPCELL_ASAP7_75t_R TAP_795 ();
 AO21x1_ASAP7_75t_R _25662_ (.A1(_07218_),
    .A2(_07152_),
    .B(_07223_),
    .Y(_07227_));
 TAPCELL_ASAP7_75t_R TAP_794 ();
 OA211x2_ASAP7_75t_R _25664_ (.A1(_07219_),
    .A2(_07225_),
    .B(_07227_),
    .C(_07077_),
    .Y(_07229_));
 TAPCELL_ASAP7_75t_R TAP_793 ();
 OA211x2_ASAP7_75t_R _25666_ (.A1(_13577_),
    .A2(_06635_),
    .B(_13618_),
    .C(_13584_),
    .Y(_07231_));
 AND3x1_ASAP7_75t_R _25667_ (.A(_13584_),
    .B(_13606_),
    .C(_06630_),
    .Y(_07232_));
 AND2x2_ASAP7_75t_R _25668_ (.A(_06634_),
    .B(_06635_),
    .Y(_07233_));
 OA211x2_ASAP7_75t_R _25669_ (.A1(_07232_),
    .A2(_07233_),
    .B(_13618_),
    .C(_13577_),
    .Y(_07234_));
 TAPCELL_ASAP7_75t_R TAP_792 ();
 TAPCELL_ASAP7_75t_R TAP_791 ();
 AND2x2_ASAP7_75t_R _25672_ (.A(_13618_),
    .B(_06635_),
    .Y(_07237_));
 NAND2x2_ASAP7_75t_R _25673_ (.A(_13618_),
    .B(_06635_),
    .Y(_07238_));
 AND2x2_ASAP7_75t_R _25674_ (.A(_02359_),
    .B(_07238_),
    .Y(_07239_));
 AOI211x1_ASAP7_75t_R _25675_ (.A1(_02360_),
    .A2(_07237_),
    .B(_07239_),
    .C(_07234_),
    .Y(_07240_));
 AO21x1_ASAP7_75t_R _25676_ (.A1(_00074_),
    .A2(_07234_),
    .B(_07240_),
    .Y(_07241_));
 AND3x4_ASAP7_75t_R _25677_ (.A(_13584_),
    .B(_06633_),
    .C(_06630_),
    .Y(_07242_));
 OA21x2_ASAP7_75t_R _25678_ (.A1(_13538_),
    .A2(_07067_),
    .B(_13804_),
    .Y(_07243_));
 NAND2x1_ASAP7_75t_R _25679_ (.A(_06979_),
    .B(_07243_),
    .Y(_07244_));
 AO221x1_ASAP7_75t_R _25680_ (.A1(_07231_),
    .A2(_07241_),
    .B1(_07242_),
    .B2(\ex_block_i.alu_adder_result_ex_o[0] ),
    .C(_07244_),
    .Y(_07245_));
 NOR2x1_ASAP7_75t_R _25681_ (.A(_07229_),
    .B(_07245_),
    .Y(_07246_));
 OA211x2_ASAP7_75t_R _25682_ (.A1(_13618_),
    .A2(_06691_),
    .B(_07217_),
    .C(_07246_),
    .Y(_07247_));
 OR4x2_ASAP7_75t_R _25683_ (.A(_07033_),
    .B(_07056_),
    .C(_07068_),
    .D(_07247_),
    .Y(_07248_));
 TAPCELL_ASAP7_75t_R TAP_790 ();
 NAND2x1_ASAP7_75t_R _25685_ (.A(_06987_),
    .B(_07248_),
    .Y(_07250_));
 OA21x2_ASAP7_75t_R _25686_ (.A1(_13848_),
    .A2(_06987_),
    .B(_07250_),
    .Y(_02656_));
 TAPCELL_ASAP7_75t_R TAP_789 ();
 TAPCELL_ASAP7_75t_R TAP_788 ();
 AND2x6_ASAP7_75t_R _25689_ (.A(net432),
    .B(_07051_),
    .Y(_07253_));
 TAPCELL_ASAP7_75t_R TAP_787 ();
 TAPCELL_ASAP7_75t_R TAP_786 ();
 AO221x1_ASAP7_75t_R _25692_ (.A1(net35),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net58),
    .C(_07036_),
    .Y(_07256_));
 INVx1_ASAP7_75t_R _25693_ (.A(_01862_),
    .Y(_07257_));
 INVx1_ASAP7_75t_R _25694_ (.A(_01870_),
    .Y(_07258_));
 TAPCELL_ASAP7_75t_R TAP_785 ();
 AO221x1_ASAP7_75t_R _25696_ (.A1(_07257_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07258_),
    .C(_07034_),
    .Y(_07260_));
 INVx1_ASAP7_75t_R _25697_ (.A(net44),
    .Y(_07261_));
 OAI22x1_ASAP7_75t_R _25698_ (.A1(_07261_),
    .A2(_01730_),
    .B1(_01854_),
    .B2(_07046_),
    .Y(_07262_));
 TAPCELL_ASAP7_75t_R TAP_784 ();
 AND2x4_ASAP7_75t_R _25700_ (.A(net432),
    .B(net433),
    .Y(_07264_));
 AO222x2_ASAP7_75t_R _25701_ (.A1(_07256_),
    .A2(_07260_),
    .B1(_07262_),
    .B2(_07044_),
    .C1(net38),
    .C2(_07264_),
    .Y(_07265_));
 TAPCELL_ASAP7_75t_R TAP_783 ();
 NAND2x1_ASAP7_75t_R _25703_ (.A(_00279_),
    .B(_07062_),
    .Y(_07267_));
 TAPCELL_ASAP7_75t_R TAP_782 ();
 AND3x1_ASAP7_75t_R _25705_ (.A(_00279_),
    .B(_01360_),
    .C(_07062_),
    .Y(_07269_));
 AO21x1_ASAP7_75t_R _25706_ (.A1(_00291_),
    .A2(_07267_),
    .B(_07269_),
    .Y(_07270_));
 NAND2x1_ASAP7_75t_R _25707_ (.A(_13817_),
    .B(_07270_),
    .Y(_07271_));
 TAPCELL_ASAP7_75t_R TAP_781 ();
 AND2x6_ASAP7_75t_R _25709_ (.A(_07218_),
    .B(_07152_),
    .Y(_07273_));
 NAND2x1_ASAP7_75t_R _25710_ (.A(_07166_),
    .B(_07223_),
    .Y(_07274_));
 OAI21x1_ASAP7_75t_R _25711_ (.A1(_07104_),
    .A2(_07166_),
    .B(_07274_),
    .Y(_07275_));
 AND2x2_ASAP7_75t_R _25712_ (.A(_07219_),
    .B(_07223_),
    .Y(_07276_));
 AO21x1_ASAP7_75t_R _25713_ (.A1(_07273_),
    .A2(_07275_),
    .B(_07276_),
    .Y(_07277_));
 OA211x2_ASAP7_75t_R _25714_ (.A1(_05077_),
    .A2(_07080_),
    .B(_07183_),
    .C(_13894_),
    .Y(_07278_));
 AOI21x1_ASAP7_75t_R _25715_ (.A1(net304),
    .A2(_07203_),
    .B(_07278_),
    .Y(_07279_));
 AO211x2_ASAP7_75t_R _25716_ (.A1(_18469_),
    .A2(_07077_),
    .B(_07200_),
    .C(_13893_),
    .Y(_07280_));
 OA211x2_ASAP7_75t_R _25717_ (.A1(_13894_),
    .A2(_07207_),
    .B(_07280_),
    .C(_07094_),
    .Y(_07281_));
 TAPCELL_ASAP7_75t_R TAP_780 ();
 AOI211x1_ASAP7_75t_R _25719_ (.A1(_07096_),
    .A2(_07279_),
    .B(_07281_),
    .C(_07090_),
    .Y(_07283_));
 TAPCELL_ASAP7_75t_R TAP_779 ();
 OA211x2_ASAP7_75t_R _25721_ (.A1(_04857_),
    .A2(_07080_),
    .B(_07189_),
    .C(_13894_),
    .Y(_07285_));
 OA211x2_ASAP7_75t_R _25722_ (.A1(_04967_),
    .A2(_07080_),
    .B(_07181_),
    .C(net304),
    .Y(_07286_));
 OR3x1_ASAP7_75t_R _25723_ (.A(_07096_),
    .B(_07285_),
    .C(_07286_),
    .Y(_07287_));
 AND3x2_ASAP7_75t_R _25724_ (.A(net305),
    .B(_07187_),
    .C(_07188_),
    .Y(_07288_));
 AND3x1_ASAP7_75t_R _25725_ (.A(_13894_),
    .B(_07167_),
    .C(_07168_),
    .Y(_07289_));
 OR3x1_ASAP7_75t_R _25726_ (.A(_07094_),
    .B(_07288_),
    .C(_07289_),
    .Y(_07290_));
 AND3x1_ASAP7_75t_R _25727_ (.A(_07090_),
    .B(_07287_),
    .C(_07290_),
    .Y(_07291_));
 TAPCELL_ASAP7_75t_R TAP_778 ();
 OA21x2_ASAP7_75t_R _25729_ (.A1(_07283_),
    .A2(_07291_),
    .B(_07273_),
    .Y(_07293_));
 AOI211x1_ASAP7_75t_R _25730_ (.A1(_16262_),
    .A2(_07077_),
    .B(_07163_),
    .C(_13894_),
    .Y(_07294_));
 AND3x2_ASAP7_75t_R _25731_ (.A(_13894_),
    .B(_07155_),
    .C(_07156_),
    .Y(_07295_));
 OA21x2_ASAP7_75t_R _25732_ (.A1(_07294_),
    .A2(_07295_),
    .B(_07094_),
    .Y(_07296_));
 XNOR2x1_ASAP7_75t_R _25733_ (.B(_07077_),
    .Y(_07297_),
    .A(_13894_));
 NAND2x1_ASAP7_75t_R _25734_ (.A(_18400_),
    .B(_07297_),
    .Y(_07298_));
 OR2x2_ASAP7_75t_R _25735_ (.A(_16020_),
    .B(_07297_),
    .Y(_07299_));
 AND3x1_ASAP7_75t_R _25736_ (.A(_07096_),
    .B(_07298_),
    .C(_07299_),
    .Y(_07300_));
 OA21x2_ASAP7_75t_R _25737_ (.A1(_07296_),
    .A2(_07300_),
    .B(_07090_),
    .Y(_07301_));
 TAPCELL_ASAP7_75t_R TAP_777 ();
 AND2x2_ASAP7_75t_R _25739_ (.A(net303),
    .B(_07173_),
    .Y(_07303_));
 AOI211x1_ASAP7_75t_R _25740_ (.A1(_18385_),
    .A2(_07080_),
    .B(_07160_),
    .C(net303),
    .Y(_07304_));
 OA21x2_ASAP7_75t_R _25741_ (.A1(_16620_),
    .A2(_07080_),
    .B(_07174_),
    .Y(_07305_));
 OA21x2_ASAP7_75t_R _25742_ (.A1(_15337_),
    .A2(_07077_),
    .B(net304),
    .Y(_07306_));
 AO221x1_ASAP7_75t_R _25743_ (.A1(_13894_),
    .A2(_07305_),
    .B1(_07306_),
    .B2(_07169_),
    .C(_07096_),
    .Y(_07307_));
 OA31x2_ASAP7_75t_R _25744_ (.A1(_07094_),
    .A2(_07303_),
    .A3(_07304_),
    .B1(_07307_),
    .Y(_07308_));
 AND2x2_ASAP7_75t_R _25745_ (.A(_07121_),
    .B(_07308_),
    .Y(_07309_));
 AND2x4_ASAP7_75t_R _25746_ (.A(_07218_),
    .B(_07125_),
    .Y(_07310_));
 OA21x2_ASAP7_75t_R _25747_ (.A1(_07301_),
    .A2(_07309_),
    .B(_07310_),
    .Y(_07311_));
 AOI211x1_ASAP7_75t_R _25748_ (.A1(_18385_),
    .A2(_07077_),
    .B(_07148_),
    .C(_13894_),
    .Y(_07312_));
 AND2x2_ASAP7_75t_R _25749_ (.A(_13894_),
    .B(_07127_),
    .Y(_07313_));
 NOR2x1_ASAP7_75t_R _25750_ (.A(_07312_),
    .B(_07313_),
    .Y(_07314_));
 AO21x1_ASAP7_75t_R _25751_ (.A1(_16262_),
    .A2(_07080_),
    .B(_07146_),
    .Y(_07315_));
 NAND3x2_ASAP7_75t_R _25752_ (.B(_07140_),
    .C(_07141_),
    .Y(_07316_),
    .A(net305));
 OA211x2_ASAP7_75t_R _25753_ (.A1(net303),
    .A2(_07315_),
    .B(_07316_),
    .C(_07094_),
    .Y(_07317_));
 AOI211x1_ASAP7_75t_R _25754_ (.A1(_07096_),
    .A2(_07314_),
    .B(_07317_),
    .C(_07090_),
    .Y(_07318_));
 AND3x1_ASAP7_75t_R _25755_ (.A(net304),
    .B(_07131_),
    .C(_07132_),
    .Y(_07319_));
 AND3x1_ASAP7_75t_R _25756_ (.A(_13894_),
    .B(_07107_),
    .C(_07108_),
    .Y(_07320_));
 AO21x1_ASAP7_75t_R _25757_ (.A1(_15401_),
    .A2(_07077_),
    .B(_07128_),
    .Y(_07321_));
 OA21x2_ASAP7_75t_R _25758_ (.A1(_15337_),
    .A2(_07080_),
    .B(_13894_),
    .Y(_07322_));
 AO221x1_ASAP7_75t_R _25759_ (.A1(net304),
    .A2(_07321_),
    .B1(_07133_),
    .B2(_07322_),
    .C(_07096_),
    .Y(_07323_));
 OA31x2_ASAP7_75t_R _25760_ (.A1(_07094_),
    .A2(_07319_),
    .A3(_07320_),
    .B1(_07323_),
    .Y(_07324_));
 AND2x2_ASAP7_75t_R _25761_ (.A(_07090_),
    .B(_07324_),
    .Y(_07325_));
 AND2x2_ASAP7_75t_R _25762_ (.A(_07073_),
    .B(_07152_),
    .Y(_07326_));
 OA21x2_ASAP7_75t_R _25763_ (.A1(_07318_),
    .A2(_07325_),
    .B(_07326_),
    .Y(_07327_));
 TAPCELL_ASAP7_75t_R TAP_776 ();
 AND2x2_ASAP7_75t_R _25765_ (.A(net303),
    .B(_07117_),
    .Y(_07329_));
 OA211x2_ASAP7_75t_R _25766_ (.A1(_04967_),
    .A2(_07077_),
    .B(_07111_),
    .C(_13894_),
    .Y(_07330_));
 OR3x1_ASAP7_75t_R _25767_ (.A(_07096_),
    .B(_07329_),
    .C(_07330_),
    .Y(_07331_));
 NOR2x1_ASAP7_75t_R _25768_ (.A(net304),
    .B(_07083_),
    .Y(_07332_));
 AO221x1_ASAP7_75t_R _25769_ (.A1(_07092_),
    .A2(_07093_),
    .B1(_07115_),
    .B2(net304),
    .C(_07332_),
    .Y(_07333_));
 NAND2x1_ASAP7_75t_R _25770_ (.A(_07086_),
    .B(_07221_),
    .Y(_07334_));
 OR3x1_ASAP7_75t_R _25771_ (.A(_07094_),
    .B(_07098_),
    .C(_07099_),
    .Y(_07335_));
 NAND2x1_ASAP7_75t_R _25772_ (.A(_00072_),
    .B(_07071_),
    .Y(_07336_));
 OA211x2_ASAP7_75t_R _25773_ (.A1(_07071_),
    .A2(_13525_),
    .B(_07336_),
    .C(_07220_),
    .Y(_07337_));
 AO211x2_ASAP7_75t_R _25774_ (.A1(_07094_),
    .A2(_07102_),
    .B(_07337_),
    .C(net304),
    .Y(_07338_));
 AND4x1_ASAP7_75t_R _25775_ (.A(_07090_),
    .B(_07334_),
    .C(_07335_),
    .D(_07338_),
    .Y(_07339_));
 AO31x2_ASAP7_75t_R _25776_ (.A1(_07121_),
    .A2(_07331_),
    .A3(_07333_),
    .B(_07339_),
    .Y(_07340_));
 AND3x1_ASAP7_75t_R _25777_ (.A(_07073_),
    .B(_07125_),
    .C(_07340_),
    .Y(_07341_));
 OR4x2_ASAP7_75t_R _25778_ (.A(_07293_),
    .B(_07311_),
    .C(_07327_),
    .D(_07341_),
    .Y(_07342_));
 TAPCELL_ASAP7_75t_R TAP_775 ();
 TAPCELL_ASAP7_75t_R TAP_774 ();
 TAPCELL_ASAP7_75t_R TAP_773 ();
 TAPCELL_ASAP7_75t_R TAP_772 ();
 TAPCELL_ASAP7_75t_R TAP_771 ();
 TAPCELL_ASAP7_75t_R TAP_770 ();
 TAPCELL_ASAP7_75t_R TAP_769 ();
 AND3x1_ASAP7_75t_R _25786_ (.A(_00076_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07350_));
 TAPCELL_ASAP7_75t_R TAP_768 ();
 AOI211x1_ASAP7_75t_R _25788_ (.A1(_00075_),
    .A2(_07238_),
    .B(_07350_),
    .C(_07234_),
    .Y(_07352_));
 AO21x1_ASAP7_75t_R _25789_ (.A1(_02361_),
    .A2(_07234_),
    .B(_07352_),
    .Y(_07353_));
 TAPCELL_ASAP7_75t_R TAP_767 ();
 AO221x1_ASAP7_75t_R _25791_ (.A1(net297),
    .A2(_07242_),
    .B1(_07353_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07355_));
 AO221x1_ASAP7_75t_R _25792_ (.A1(_07077_),
    .A2(_07277_),
    .B1(_07342_),
    .B2(_07215_),
    .C(_07355_),
    .Y(_07356_));
 TAPCELL_ASAP7_75t_R TAP_766 ();
 TAPCELL_ASAP7_75t_R TAP_765 ();
 AND2x4_ASAP7_75t_R _25795_ (.A(_05616_),
    .B(_06949_),
    .Y(_07359_));
 AOI22x1_ASAP7_75t_R _25796_ (.A1(_06938_),
    .A2(_07359_),
    .B1(_06946_),
    .B2(_05656_),
    .Y(_07360_));
 TAPCELL_ASAP7_75t_R TAP_764 ();
 TAPCELL_ASAP7_75t_R TAP_763 ();
 OA22x2_ASAP7_75t_R _25799_ (.A1(_01518_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01487_),
    .Y(_07363_));
 OA22x2_ASAP7_75t_R _25800_ (.A1(_01944_),
    .A2(_06938_),
    .B1(_06994_),
    .B2(_01912_),
    .Y(_07364_));
 TAPCELL_ASAP7_75t_R TAP_762 ();
 NAND2x1_ASAP7_75t_R _25802_ (.A(net3646),
    .B(_06947_),
    .Y(_07366_));
 NAND2x2_ASAP7_75t_R _25803_ (.A(_05693_),
    .B(_06965_),
    .Y(_07367_));
 TAPCELL_ASAP7_75t_R TAP_761 ();
 OR2x6_ASAP7_75t_R _25805_ (.A(_05589_),
    .B(_06938_),
    .Y(_07369_));
 TAPCELL_ASAP7_75t_R TAP_760 ();
 OA222x2_ASAP7_75t_R _25807_ (.A1(_01576_),
    .A2(_07000_),
    .B1(_07367_),
    .B2(_02138_),
    .C1(_07369_),
    .C2(_00658_),
    .Y(_07371_));
 OA211x2_ASAP7_75t_R _25808_ (.A1(_06990_),
    .A2(_07364_),
    .B(_07366_),
    .C(_07371_),
    .Y(_07372_));
 TAPCELL_ASAP7_75t_R TAP_759 ();
 TAPCELL_ASAP7_75t_R TAP_758 ();
 TAPCELL_ASAP7_75t_R TAP_757 ();
 OA22x2_ASAP7_75t_R _25812_ (.A1(_02171_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02065_),
    .Y(_07376_));
 TAPCELL_ASAP7_75t_R TAP_756 ();
 TAPCELL_ASAP7_75t_R TAP_755 ();
 OA222x2_ASAP7_75t_R _25815_ (.A1(_01994_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02097_),
    .C1(_07028_),
    .C2(_02028_),
    .Y(_07379_));
 OA21x2_ASAP7_75t_R _25816_ (.A1(_07021_),
    .A2(_07376_),
    .B(_07379_),
    .Y(_07380_));
 OA211x2_ASAP7_75t_R _25817_ (.A1(_07360_),
    .A2(_07363_),
    .B(_07372_),
    .C(_07380_),
    .Y(_07381_));
 NAND2x1_ASAP7_75t_R _25818_ (.A(_06981_),
    .B(_07381_),
    .Y(_07382_));
 AO21x1_ASAP7_75t_R _25819_ (.A1(_07271_),
    .A2(_07356_),
    .B(_07382_),
    .Y(_07383_));
 OA21x2_ASAP7_75t_R _25820_ (.A1(_06981_),
    .A2(_07265_),
    .B(_07383_),
    .Y(_07384_));
 NOR2x1_ASAP7_75t_R _25821_ (.A(_01708_),
    .B(_06987_),
    .Y(_07385_));
 AO21x1_ASAP7_75t_R _25822_ (.A1(_06987_),
    .A2(_07384_),
    .B(_07385_),
    .Y(_02657_));
 AO21x1_ASAP7_75t_R _25823_ (.A1(_07107_),
    .A2(_07108_),
    .B(_13894_),
    .Y(_07386_));
 OA211x2_ASAP7_75t_R _25824_ (.A1(net303),
    .A2(_07117_),
    .B(_07386_),
    .C(_07096_),
    .Y(_07387_));
 AND2x2_ASAP7_75t_R _25825_ (.A(_07094_),
    .B(_07136_),
    .Y(_07388_));
 OR3x1_ASAP7_75t_R _25826_ (.A(_07121_),
    .B(_07387_),
    .C(_07388_),
    .Y(_07389_));
 OA21x2_ASAP7_75t_R _25827_ (.A1(_07147_),
    .A2(_07149_),
    .B(_07094_),
    .Y(_07390_));
 AND2x2_ASAP7_75t_R _25828_ (.A(_07096_),
    .B(_07130_),
    .Y(_07391_));
 OR3x1_ASAP7_75t_R _25829_ (.A(_07090_),
    .B(_07390_),
    .C(_07391_),
    .Y(_07392_));
 NAND2x1_ASAP7_75t_R _25830_ (.A(_07389_),
    .B(_07392_),
    .Y(_07393_));
 TAPCELL_ASAP7_75t_R TAP_754 ();
 OA211x2_ASAP7_75t_R _25832_ (.A1(_05077_),
    .A2(_07077_),
    .B(_07114_),
    .C(_07094_),
    .Y(_07395_));
 NOR2x1_ASAP7_75t_R _25833_ (.A(_07094_),
    .B(_07086_),
    .Y(_07396_));
 OR2x2_ASAP7_75t_R _25834_ (.A(_07395_),
    .B(_07396_),
    .Y(_07397_));
 NOR2x1_ASAP7_75t_R _25835_ (.A(_07094_),
    .B(_07083_),
    .Y(_07398_));
 OA211x2_ASAP7_75t_R _25836_ (.A1(_04967_),
    .A2(_07077_),
    .B(_07111_),
    .C(_07094_),
    .Y(_07399_));
 OR3x1_ASAP7_75t_R _25837_ (.A(_13894_),
    .B(_07398_),
    .C(_07399_),
    .Y(_07400_));
 OA21x2_ASAP7_75t_R _25838_ (.A1(net304),
    .A2(_07397_),
    .B(_07400_),
    .Y(_07401_));
 OR3x1_ASAP7_75t_R _25839_ (.A(_07096_),
    .B(_07100_),
    .C(_07103_),
    .Y(_07402_));
 OA211x2_ASAP7_75t_R _25840_ (.A1(_07094_),
    .A2(_07223_),
    .B(_07402_),
    .C(_07090_),
    .Y(_07403_));
 NAND2x1_ASAP7_75t_R _25841_ (.A(_07073_),
    .B(_07125_),
    .Y(_07404_));
 AOI211x1_ASAP7_75t_R _25842_ (.A1(_07121_),
    .A2(_07401_),
    .B(_07403_),
    .C(_07404_),
    .Y(_07405_));
 AO21x1_ASAP7_75t_R _25843_ (.A1(_07326_),
    .A2(_07393_),
    .B(_07405_),
    .Y(_07406_));
 NOR2x1_ASAP7_75t_R _25844_ (.A(_07096_),
    .B(_07191_),
    .Y(_07407_));
 NOR2x1_ASAP7_75t_R _25845_ (.A(_07094_),
    .B(_07171_),
    .Y(_07408_));
 OR3x1_ASAP7_75t_R _25846_ (.A(_07121_),
    .B(_07407_),
    .C(_07408_),
    .Y(_07409_));
 NOR2x1_ASAP7_75t_R _25847_ (.A(_07096_),
    .B(_07205_),
    .Y(_07410_));
 AO211x2_ASAP7_75t_R _25848_ (.A1(_07096_),
    .A2(_07185_),
    .B(_07410_),
    .C(_07090_),
    .Y(_07411_));
 AO221x2_ASAP7_75t_R _25849_ (.A1(_07092_),
    .A2(_07093_),
    .B1(_07138_),
    .B2(_07139_),
    .C(_07142_),
    .Y(_07412_));
 OAI21x1_ASAP7_75t_R _25850_ (.A1(_07096_),
    .A2(_07159_),
    .B(_07412_),
    .Y(_07413_));
 AO211x2_ASAP7_75t_R _25851_ (.A1(_13894_),
    .A2(_07173_),
    .B(_07175_),
    .C(_07096_),
    .Y(_07414_));
 OA31x2_ASAP7_75t_R _25852_ (.A1(_07094_),
    .A2(_07161_),
    .A3(_07164_),
    .B1(_07414_),
    .Y(_07415_));
 NAND2x1_ASAP7_75t_R _25853_ (.A(_07121_),
    .B(_07415_),
    .Y(_07416_));
 OA21x2_ASAP7_75t_R _25854_ (.A1(_07121_),
    .A2(_07413_),
    .B(_07416_),
    .Y(_07417_));
 AO32x1_ASAP7_75t_R _25855_ (.A1(_07273_),
    .A2(_07409_),
    .A3(_07411_),
    .B1(_07310_),
    .B2(_07417_),
    .Y(_07418_));
 OR3x1_ASAP7_75t_R _25856_ (.A(_07216_),
    .B(_07406_),
    .C(_07418_),
    .Y(_07419_));
 TAPCELL_ASAP7_75t_R TAP_753 ();
 AO32x1_ASAP7_75t_R _25858_ (.A1(_01364_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00663_),
    .Y(_07421_));
 TAPCELL_ASAP7_75t_R TAP_752 ();
 AND3x1_ASAP7_75t_R _25860_ (.A(_07334_),
    .B(_07335_),
    .C(_07338_),
    .Y(_07423_));
 OA21x2_ASAP7_75t_R _25861_ (.A1(_07090_),
    .A2(_07125_),
    .B(_07223_),
    .Y(_07424_));
 AO21x1_ASAP7_75t_R _25862_ (.A1(_07197_),
    .A2(_07423_),
    .B(_07424_),
    .Y(_07425_));
 AND2x6_ASAP7_75t_R _25863_ (.A(_07218_),
    .B(_07077_),
    .Y(_07426_));
 TAPCELL_ASAP7_75t_R TAP_751 ();
 AND3x1_ASAP7_75t_R _25865_ (.A(_00078_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07428_));
 AOI211x1_ASAP7_75t_R _25866_ (.A1(_00077_),
    .A2(_07238_),
    .B(_07428_),
    .C(_07234_),
    .Y(_07429_));
 AO21x2_ASAP7_75t_R _25867_ (.A1(_02362_),
    .A2(_07234_),
    .B(_07429_),
    .Y(_07430_));
 TAPCELL_ASAP7_75t_R TAP_750 ();
 AO222x2_ASAP7_75t_R _25869_ (.A1(net171),
    .A2(_07242_),
    .B1(_07425_),
    .B2(_07426_),
    .C1(_07430_),
    .C2(_07231_),
    .Y(_07432_));
 NOR2x1_ASAP7_75t_R _25870_ (.A(_13817_),
    .B(_07432_),
    .Y(_07433_));
 AO21x1_ASAP7_75t_R _25871_ (.A1(_13817_),
    .A2(_07421_),
    .B(_07433_),
    .Y(_07434_));
 TAPCELL_ASAP7_75t_R TAP_749 ();
 TAPCELL_ASAP7_75t_R TAP_748 ();
 OAI22x1_ASAP7_75t_R _25874_ (.A1(_01517_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01486_),
    .Y(_07437_));
 AO32x2_ASAP7_75t_R _25875_ (.A1(_05681_),
    .A2(_05676_),
    .A3(_06938_),
    .B1(_05644_),
    .B2(_05656_),
    .Y(_07438_));
 OAI22x1_ASAP7_75t_R _25876_ (.A1(_02170_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02064_),
    .Y(_07439_));
 AND2x4_ASAP7_75t_R _25877_ (.A(_13894_),
    .B(_05663_),
    .Y(_07440_));
 AOI211x1_ASAP7_75t_R _25878_ (.A1(net302),
    .A2(_07440_),
    .B(_05621_),
    .C(_05623_),
    .Y(_07441_));
 AOI22x1_ASAP7_75t_R _25879_ (.A1(_07437_),
    .A2(_07438_),
    .B1(_07439_),
    .B2(_07441_),
    .Y(_07442_));
 AND3x2_ASAP7_75t_R _25880_ (.A(_05586_),
    .B(_05644_),
    .C(_06945_),
    .Y(_07443_));
 NAND2x1_ASAP7_75t_R _25881_ (.A(net3523),
    .B(_07443_),
    .Y(_07444_));
 TAPCELL_ASAP7_75t_R TAP_747 ();
 TAPCELL_ASAP7_75t_R TAP_746 ();
 NAND3x2_ASAP7_75t_R _25884_ (.B(_05627_),
    .C(_05630_),
    .Y(_07447_),
    .A(_05601_));
 OAI22x1_ASAP7_75t_R _25885_ (.A1(_02034_),
    .A2(_05589_),
    .B1(_07447_),
    .B2(_02137_),
    .Y(_07448_));
 INVx1_ASAP7_75t_R _25886_ (.A(_01943_),
    .Y(_07449_));
 AND2x2_ASAP7_75t_R _25887_ (.A(_05602_),
    .B(_06960_),
    .Y(_07450_));
 AO21x1_ASAP7_75t_R _25888_ (.A1(_07449_),
    .A2(_05632_),
    .B(_07450_),
    .Y(_07451_));
 AOI22x1_ASAP7_75t_R _25889_ (.A1(_05693_),
    .A2(_07448_),
    .B1(_07451_),
    .B2(_07440_),
    .Y(_07452_));
 TAPCELL_ASAP7_75t_R TAP_745 ();
 TAPCELL_ASAP7_75t_R TAP_744 ();
 TAPCELL_ASAP7_75t_R PHY_743 ();
 OA222x2_ASAP7_75t_R _25893_ (.A1(_01993_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02096_),
    .C1(_07369_),
    .C2(_01575_),
    .Y(_07456_));
 INVx1_ASAP7_75t_R _25894_ (.A(_05641_),
    .Y(_07457_));
 OR3x1_ASAP7_75t_R _25895_ (.A(_13523_),
    .B(_14179_),
    .C(_06937_),
    .Y(_07458_));
 AND2x2_ASAP7_75t_R _25896_ (.A(_02027_),
    .B(_13894_),
    .Y(_07459_));
 AO21x1_ASAP7_75t_R _25897_ (.A1(_01911_),
    .A2(_13893_),
    .B(_07459_),
    .Y(_07460_));
 OA33x2_ASAP7_75t_R _25898_ (.A1(_01315_),
    .A2(_07457_),
    .A3(_06992_),
    .B1(_07458_),
    .B2(_07460_),
    .B3(_07447_),
    .Y(_07461_));
 AND5x2_ASAP7_75t_R _25899_ (.A(_07442_),
    .B(net3524),
    .C(_07452_),
    .D(_07456_),
    .E(_07461_),
    .Y(_07462_));
 AND4x2_ASAP7_75t_R _25900_ (.A(_06981_),
    .B(_07419_),
    .C(_07434_),
    .D(_07462_),
    .Y(_07463_));
 AO221x1_ASAP7_75t_R _25901_ (.A1(net36),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net28),
    .C(_07036_),
    .Y(_07464_));
 INVx1_ASAP7_75t_R _25902_ (.A(_01861_),
    .Y(_07465_));
 INVx1_ASAP7_75t_R _25903_ (.A(_01869_),
    .Y(_07466_));
 AO221x1_ASAP7_75t_R _25904_ (.A1(_07465_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07466_),
    .C(_07034_),
    .Y(_07467_));
 INVx1_ASAP7_75t_R _25905_ (.A(net2395),
    .Y(_07468_));
 OAI22x1_ASAP7_75t_R _25906_ (.A1(_07468_),
    .A2(_01730_),
    .B1(_01853_),
    .B2(_07046_),
    .Y(_07469_));
 AO222x2_ASAP7_75t_R _25907_ (.A1(net3772),
    .A2(_07264_),
    .B1(_07464_),
    .B2(_07467_),
    .C1(_07469_),
    .C2(_07044_),
    .Y(_07470_));
 NOR2x2_ASAP7_75t_R _25908_ (.A(net290),
    .B(net3773),
    .Y(_07471_));
 NOR2x2_ASAP7_75t_R _25909_ (.A(_07463_),
    .B(_07471_),
    .Y(_07472_));
 NOR2x1_ASAP7_75t_R _25910_ (.A(_01707_),
    .B(net288),
    .Y(_07473_));
 AO21x1_ASAP7_75t_R _25911_ (.A1(net288),
    .A2(_07472_),
    .B(_07473_),
    .Y(_02658_));
 AO21x2_ASAP7_75t_R _25912_ (.A1(net310),
    .A2(_06977_),
    .B(_06980_),
    .Y(_07474_));
 TAPCELL_ASAP7_75t_R PHY_742 ();
 TAPCELL_ASAP7_75t_R PHY_741 ();
 TAPCELL_ASAP7_75t_R PHY_740 ();
 TAPCELL_ASAP7_75t_R PHY_739 ();
 OR3x2_ASAP7_75t_R _25917_ (.A(_13894_),
    .B(_07395_),
    .C(_07396_),
    .Y(_07479_));
 NOR2x1_ASAP7_75t_R _25918_ (.A(_07096_),
    .B(_07083_),
    .Y(_07480_));
 AND2x2_ASAP7_75t_R _25919_ (.A(_07096_),
    .B(_07102_),
    .Y(_07481_));
 OR3x2_ASAP7_75t_R _25920_ (.A(net303),
    .B(_07480_),
    .C(_07481_),
    .Y(_07482_));
 AND2x2_ASAP7_75t_R _25921_ (.A(_07090_),
    .B(_07222_),
    .Y(_07483_));
 AO31x2_ASAP7_75t_R _25922_ (.A1(_07121_),
    .A2(_07479_),
    .A3(_07482_),
    .B(_07483_),
    .Y(_07484_));
 AO221x1_ASAP7_75t_R _25923_ (.A1(net304),
    .A2(_07321_),
    .B1(_07133_),
    .B2(_07322_),
    .C(_07094_),
    .Y(_07485_));
 OA31x2_ASAP7_75t_R _25924_ (.A1(_07096_),
    .A2(_07312_),
    .A3(_07313_),
    .B1(_07485_),
    .Y(_07486_));
 AND2x2_ASAP7_75t_R _25925_ (.A(_07121_),
    .B(_07486_),
    .Y(_07487_));
 OR2x2_ASAP7_75t_R _25926_ (.A(_07319_),
    .B(_07320_),
    .Y(_07488_));
 OR3x1_ASAP7_75t_R _25927_ (.A(_07094_),
    .B(_07329_),
    .C(_07330_),
    .Y(_07489_));
 OA211x2_ASAP7_75t_R _25928_ (.A1(_07096_),
    .A2(_07488_),
    .B(_07489_),
    .C(_07090_),
    .Y(_07490_));
 TAPCELL_ASAP7_75t_R PHY_738 ();
 OA21x2_ASAP7_75t_R _25930_ (.A1(_07487_),
    .A2(_07490_),
    .B(_07152_),
    .Y(_07492_));
 AO21x1_ASAP7_75t_R _25931_ (.A1(_07125_),
    .A2(_07484_),
    .B(_07492_),
    .Y(_07493_));
 AOI21x1_ASAP7_75t_R _25932_ (.A1(_07298_),
    .A2(_07299_),
    .B(_07096_),
    .Y(_07494_));
 OA211x2_ASAP7_75t_R _25933_ (.A1(net303),
    .A2(_07315_),
    .B(_07316_),
    .C(_07096_),
    .Y(_07495_));
 NOR2x1_ASAP7_75t_R _25934_ (.A(_07494_),
    .B(_07495_),
    .Y(_07496_));
 OR3x1_ASAP7_75t_R _25935_ (.A(_07096_),
    .B(_07303_),
    .C(_07304_),
    .Y(_07497_));
 OR3x1_ASAP7_75t_R _25936_ (.A(_07094_),
    .B(_07294_),
    .C(_07295_),
    .Y(_07498_));
 AND3x1_ASAP7_75t_R _25937_ (.A(_07121_),
    .B(_07497_),
    .C(_07498_),
    .Y(_07499_));
 AO21x1_ASAP7_75t_R _25938_ (.A1(_07090_),
    .A2(_07496_),
    .B(_07499_),
    .Y(_07500_));
 AO22x1_ASAP7_75t_R _25939_ (.A1(_13894_),
    .A2(_07305_),
    .B1(_07306_),
    .B2(_07169_),
    .Y(_07501_));
 OR3x1_ASAP7_75t_R _25940_ (.A(_07096_),
    .B(_07288_),
    .C(_07289_),
    .Y(_07502_));
 OA21x2_ASAP7_75t_R _25941_ (.A1(_07094_),
    .A2(_07501_),
    .B(_07502_),
    .Y(_07503_));
 AOI211x1_ASAP7_75t_R _25942_ (.A1(net304),
    .A2(_07182_),
    .B(_07285_),
    .C(_07094_),
    .Y(_07504_));
 AOI211x1_ASAP7_75t_R _25943_ (.A1(_07094_),
    .A2(_07279_),
    .B(_07504_),
    .C(_07090_),
    .Y(_07505_));
 AO21x1_ASAP7_75t_R _25944_ (.A1(_07090_),
    .A2(_07503_),
    .B(_07505_),
    .Y(_07506_));
 AO22x1_ASAP7_75t_R _25945_ (.A1(_07310_),
    .A2(_07500_),
    .B1(_07506_),
    .B2(_07273_),
    .Y(_07507_));
 AO21x1_ASAP7_75t_R _25946_ (.A1(_07073_),
    .A2(_07493_),
    .B(_07507_),
    .Y(_07508_));
 TAPCELL_ASAP7_75t_R PHY_737 ();
 INVx1_ASAP7_75t_R _25948_ (.A(_07197_),
    .Y(_07510_));
 NOR3x2_ASAP7_75t_R _25949_ (.B(_07100_),
    .C(_07103_),
    .Y(_07511_),
    .A(_07094_));
 AOI211x1_ASAP7_75t_R _25950_ (.A1(_07094_),
    .A2(_07088_),
    .B(_07510_),
    .C(_07511_),
    .Y(_07512_));
 OR2x2_ASAP7_75t_R _25951_ (.A(_07424_),
    .B(_07512_),
    .Y(_07513_));
 AND3x1_ASAP7_75t_R _25952_ (.A(_00080_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07514_));
 AOI211x1_ASAP7_75t_R _25953_ (.A1(_00079_),
    .A2(_07238_),
    .B(_07514_),
    .C(_07234_),
    .Y(_07515_));
 AO21x1_ASAP7_75t_R _25954_ (.A1(_02363_),
    .A2(_07234_),
    .B(_07515_),
    .Y(_07516_));
 AO222x2_ASAP7_75t_R _25955_ (.A1(net174),
    .A2(_07242_),
    .B1(_07426_),
    .B2(_07513_),
    .C1(_07516_),
    .C2(_07231_),
    .Y(_07517_));
 NAND2x1_ASAP7_75t_R _25956_ (.A(_00665_),
    .B(_07065_),
    .Y(_07518_));
 AND2x4_ASAP7_75t_R _25957_ (.A(_07060_),
    .B(_07062_),
    .Y(_07519_));
 INVx1_ASAP7_75t_R _25958_ (.A(_07519_),
    .Y(_07520_));
 OA21x2_ASAP7_75t_R _25959_ (.A1(_02231_),
    .A2(_07520_),
    .B(_13817_),
    .Y(_07521_));
 NAND3x2_ASAP7_75t_R _25960_ (.B(_06942_),
    .C(_06960_),
    .Y(_07522_),
    .A(_06956_));
 TAPCELL_ASAP7_75t_R PHY_736 ();
 OAI22x1_ASAP7_75t_R _25962_ (.A1(_00081_),
    .A2(_07369_),
    .B1(_07522_),
    .B2(_01946_),
    .Y(_07524_));
 TAPCELL_ASAP7_75t_R PHY_735 ();
 OA22x2_ASAP7_75t_R _25964_ (.A1(_01992_),
    .A2(_05589_),
    .B1(_06990_),
    .B2(_02026_),
    .Y(_07526_));
 TAPCELL_ASAP7_75t_R PHY_734 ();
 OAI21x1_ASAP7_75t_R _25966_ (.A1(_07023_),
    .A2(_07526_),
    .B(_07004_),
    .Y(_07528_));
 AND2x2_ASAP7_75t_R _25967_ (.A(net3543),
    .B(_06947_),
    .Y(_07529_));
 INVx2_ASAP7_75t_R _25968_ (.A(_06994_),
    .Y(_07530_));
 OAI22x1_ASAP7_75t_R _25969_ (.A1(_02095_),
    .A2(_05589_),
    .B1(_06990_),
    .B2(_01910_),
    .Y(_07531_));
 AND4x1_ASAP7_75t_R _25970_ (.A(_06236_),
    .B(_05693_),
    .C(_06949_),
    .D(_06941_),
    .Y(_07532_));
 AO21x1_ASAP7_75t_R _25971_ (.A1(_07530_),
    .A2(_07531_),
    .B(_07532_),
    .Y(_07533_));
 TAPCELL_ASAP7_75t_R PHY_733 ();
 OAI22x1_ASAP7_75t_R _25973_ (.A1(_02136_),
    .A2(_06992_),
    .B1(_06938_),
    .B2(_01942_),
    .Y(_07535_));
 AO21x1_ASAP7_75t_R _25974_ (.A1(net3513),
    .A2(_06942_),
    .B(_07535_),
    .Y(_07536_));
 OAI22x1_ASAP7_75t_R _25975_ (.A1(_01516_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01485_),
    .Y(_07537_));
 OAI22x1_ASAP7_75t_R _25976_ (.A1(_02169_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02063_),
    .Y(_07538_));
 AO222x2_ASAP7_75t_R _25977_ (.A1(_06965_),
    .A2(_07536_),
    .B1(_07537_),
    .B2(_06950_),
    .C1(_07538_),
    .C2(_06940_),
    .Y(_07539_));
 OR5x2_ASAP7_75t_R _25978_ (.A(_07524_),
    .B(_07528_),
    .C(_07529_),
    .D(_07533_),
    .E(_07539_),
    .Y(_07540_));
 AO221x1_ASAP7_75t_R _25979_ (.A1(net308),
    .A2(_07517_),
    .B1(_07518_),
    .B2(_07521_),
    .C(_07540_),
    .Y(_07541_));
 AO21x1_ASAP7_75t_R _25980_ (.A1(_07215_),
    .A2(_07508_),
    .B(_07541_),
    .Y(_07542_));
 NAND2x2_ASAP7_75t_R _25981_ (.A(net310),
    .B(_06977_),
    .Y(_07543_));
 AO221x1_ASAP7_75t_R _25982_ (.A1(net37),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net29),
    .C(_07036_),
    .Y(_07544_));
 INVx1_ASAP7_75t_R _25983_ (.A(_01860_),
    .Y(_07545_));
 INVx1_ASAP7_75t_R _25984_ (.A(_01868_),
    .Y(_07546_));
 AO221x1_ASAP7_75t_R _25985_ (.A1(_07545_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07546_),
    .C(_07034_),
    .Y(_07547_));
 INVx1_ASAP7_75t_R _25986_ (.A(net46),
    .Y(_07548_));
 OAI22x1_ASAP7_75t_R _25987_ (.A1(_07548_),
    .A2(_01730_),
    .B1(_01852_),
    .B2(_07046_),
    .Y(_07549_));
 AO22x1_ASAP7_75t_R _25988_ (.A1(net52),
    .A2(_07264_),
    .B1(_07549_),
    .B2(_07044_),
    .Y(_07550_));
 AO221x2_ASAP7_75t_R _25989_ (.A1(_06979_),
    .A2(_07543_),
    .B1(_07544_),
    .B2(_07547_),
    .C(_07550_),
    .Y(_07551_));
 OA21x2_ASAP7_75t_R _25990_ (.A1(_07474_),
    .A2(_07542_),
    .B(_07551_),
    .Y(_07552_));
 NOR2x1_ASAP7_75t_R _25991_ (.A(_01706_),
    .B(_06987_),
    .Y(_07553_));
 AO21x1_ASAP7_75t_R _25992_ (.A1(_06987_),
    .A2(_07552_),
    .B(_07553_),
    .Y(_02659_));
 TAPCELL_ASAP7_75t_R PHY_732 ();
 TAPCELL_ASAP7_75t_R PHY_731 ();
 TAPCELL_ASAP7_75t_R PHY_730 ();
 AND3x1_ASAP7_75t_R _25996_ (.A(_00083_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07557_));
 AOI211x1_ASAP7_75t_R _25997_ (.A1(_00082_),
    .A2(_07238_),
    .B(_07557_),
    .C(_07234_),
    .Y(_07558_));
 AO21x1_ASAP7_75t_R _25998_ (.A1(_02364_),
    .A2(_07234_),
    .B(_07558_),
    .Y(_07559_));
 TAPCELL_ASAP7_75t_R PHY_729 ();
 AO21x2_ASAP7_75t_R _26000_ (.A1(_07273_),
    .A2(_07484_),
    .B(_07276_),
    .Y(_07561_));
 AO222x2_ASAP7_75t_R _26001_ (.A1(net175),
    .A2(_07242_),
    .B1(_07559_),
    .B2(_07231_),
    .C1(_07561_),
    .C2(_07077_),
    .Y(_07562_));
 AO32x1_ASAP7_75t_R _26002_ (.A1(_01376_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00668_),
    .Y(_07563_));
 NAND2x1_ASAP7_75t_R _26003_ (.A(_13817_),
    .B(_07563_),
    .Y(_07564_));
 OAI21x1_ASAP7_75t_R _26004_ (.A1(_13817_),
    .A2(_07562_),
    .B(_07564_),
    .Y(_07565_));
 OA211x2_ASAP7_75t_R _26005_ (.A1(_13894_),
    .A2(_07127_),
    .B(_07129_),
    .C(_07094_),
    .Y(_07566_));
 AO211x2_ASAP7_75t_R _26006_ (.A1(_07096_),
    .A2(_07136_),
    .B(_07566_),
    .C(_07090_),
    .Y(_07567_));
 OA31x2_ASAP7_75t_R _26007_ (.A1(_07121_),
    .A2(_07113_),
    .A3(_07120_),
    .B1(_07567_),
    .Y(_07568_));
 AOI211x1_ASAP7_75t_R _26008_ (.A1(_07094_),
    .A2(_07088_),
    .B(_07511_),
    .C(_07090_),
    .Y(_07569_));
 AO21x1_ASAP7_75t_R _26009_ (.A1(_07090_),
    .A2(_07223_),
    .B(_07152_),
    .Y(_07570_));
 OA22x2_ASAP7_75t_R _26010_ (.A1(_07125_),
    .A2(_07568_),
    .B1(_07569_),
    .B2(_07570_),
    .Y(_07571_));
 OR3x1_ASAP7_75t_R _26011_ (.A(_07121_),
    .B(_07147_),
    .C(_07149_),
    .Y(_07572_));
 OA21x2_ASAP7_75t_R _26012_ (.A1(_07090_),
    .A2(_07159_),
    .B(_07572_),
    .Y(_07573_));
 OR3x1_ASAP7_75t_R _26013_ (.A(_07090_),
    .B(_07161_),
    .C(_07164_),
    .Y(_07574_));
 NAND2x1_ASAP7_75t_R _26014_ (.A(_07090_),
    .B(_07143_),
    .Y(_07575_));
 AND3x1_ASAP7_75t_R _26015_ (.A(_07094_),
    .B(_07574_),
    .C(_07575_),
    .Y(_07576_));
 AO21x1_ASAP7_75t_R _26016_ (.A1(_07096_),
    .A2(_07573_),
    .B(_07576_),
    .Y(_07577_));
 TAPCELL_ASAP7_75t_R PHY_728 ();
 OR2x2_ASAP7_75t_R _26018_ (.A(_07096_),
    .B(_07171_),
    .Y(_07579_));
 OA21x2_ASAP7_75t_R _26019_ (.A1(_07094_),
    .A2(_07176_),
    .B(_07579_),
    .Y(_07580_));
 AO33x2_ASAP7_75t_R _26020_ (.A1(_07218_),
    .A2(_07197_),
    .A3(_07193_),
    .B1(_07273_),
    .B2(_07580_),
    .B3(_07090_),
    .Y(_07581_));
 AO221x1_ASAP7_75t_R _26021_ (.A1(_07073_),
    .A2(_07571_),
    .B1(_07577_),
    .B2(_07310_),
    .C(_07581_),
    .Y(_07582_));
 NAND2x1_ASAP7_75t_R _26022_ (.A(_07215_),
    .B(_07582_),
    .Y(_07583_));
 OAI22x1_ASAP7_75t_R _26023_ (.A1(_01941_),
    .A2(_06938_),
    .B1(_06994_),
    .B2(_01909_),
    .Y(_07584_));
 TAPCELL_ASAP7_75t_R PHY_727 ();
 OA21x2_ASAP7_75t_R _26025_ (.A1(_02135_),
    .A2(_07367_),
    .B(_07004_),
    .Y(_07586_));
 OAI21x1_ASAP7_75t_R _26026_ (.A1(_01991_),
    .A2(_07024_),
    .B(_07586_),
    .Y(_07587_));
 AO21x2_ASAP7_75t_R _26027_ (.A1(_06965_),
    .A2(_07584_),
    .B(_07587_),
    .Y(_07588_));
 TAPCELL_ASAP7_75t_R PHY_726 ();
 OAI22x1_ASAP7_75t_R _26029_ (.A1(_02168_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02062_),
    .Y(_07590_));
 OAI22x1_ASAP7_75t_R _26030_ (.A1(_01515_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01484_),
    .Y(_07591_));
 TAPCELL_ASAP7_75t_R PHY_725 ();
 TAPCELL_ASAP7_75t_R PHY_724 ();
 TAPCELL_ASAP7_75t_R PHY_723 ();
 OA222x2_ASAP7_75t_R _26034_ (.A1(_02094_),
    .A2(_07026_),
    .B1(_07028_),
    .B2(_02025_),
    .C1(_00084_),
    .C2(_07369_),
    .Y(_07595_));
 INVx1_ASAP7_75t_R _26035_ (.A(_07595_),
    .Y(_07596_));
 AO221x1_ASAP7_75t_R _26036_ (.A1(_06940_),
    .A2(_07590_),
    .B1(_07591_),
    .B2(_06950_),
    .C(_07596_),
    .Y(_07597_));
 AOI211x1_ASAP7_75t_R _26037_ (.A1(net3384),
    .A2(_06947_),
    .B(_07588_),
    .C(_07597_),
    .Y(_07598_));
 AND4x2_ASAP7_75t_R _26038_ (.A(net290),
    .B(_07565_),
    .C(_07583_),
    .D(_07598_),
    .Y(_07599_));
 AO221x1_ASAP7_75t_R _26039_ (.A1(net39),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net30),
    .C(_07036_),
    .Y(_07600_));
 INVx1_ASAP7_75t_R _26040_ (.A(_01859_),
    .Y(_07601_));
 INVx1_ASAP7_75t_R _26041_ (.A(_01867_),
    .Y(_07602_));
 AO221x1_ASAP7_75t_R _26042_ (.A1(_07601_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07602_),
    .C(_07034_),
    .Y(_07603_));
 INVx1_ASAP7_75t_R _26043_ (.A(net47),
    .Y(_07604_));
 OAI22x1_ASAP7_75t_R _26044_ (.A1(_07604_),
    .A2(_01730_),
    .B1(_01851_),
    .B2(_07046_),
    .Y(_07605_));
 AO222x2_ASAP7_75t_R _26045_ (.A1(net53),
    .A2(_07264_),
    .B1(_07600_),
    .B2(_07603_),
    .C1(_07605_),
    .C2(_07044_),
    .Y(_07606_));
 NOR2x1_ASAP7_75t_R _26046_ (.A(net290),
    .B(_07606_),
    .Y(_07607_));
 NOR2x2_ASAP7_75t_R _26047_ (.A(_07599_),
    .B(_07607_),
    .Y(_07608_));
 NOR2x1_ASAP7_75t_R _26048_ (.A(_01705_),
    .B(net288),
    .Y(_07609_));
 AO21x1_ASAP7_75t_R _26049_ (.A1(net288),
    .A2(_07608_),
    .B(_07609_),
    .Y(_02660_));
 TAPCELL_ASAP7_75t_R PHY_722 ();
 TAPCELL_ASAP7_75t_R PHY_721 ();
 AND2x2_ASAP7_75t_R _26052_ (.A(_07121_),
    .B(_07401_),
    .Y(_07612_));
 INVx1_ASAP7_75t_R _26053_ (.A(_07104_),
    .Y(_07613_));
 INVx1_ASAP7_75t_R _26054_ (.A(_07095_),
    .Y(_07614_));
 AO21x1_ASAP7_75t_R _26055_ (.A1(_07090_),
    .A2(_07096_),
    .B(_07125_),
    .Y(_07615_));
 AO32x1_ASAP7_75t_R _26056_ (.A1(_07613_),
    .A2(_07614_),
    .A3(_07152_),
    .B1(_07223_),
    .B2(_07615_),
    .Y(_07616_));
 AO21x2_ASAP7_75t_R _26057_ (.A1(_07152_),
    .A2(_07612_),
    .B(_07616_),
    .Y(_07617_));
 NAND2x1_ASAP7_75t_R _26058_ (.A(_07426_),
    .B(_07617_),
    .Y(_07618_));
 TAPCELL_ASAP7_75t_R PHY_720 ();
 OR2x2_ASAP7_75t_R _26060_ (.A(_07090_),
    .B(_07324_),
    .Y(_07620_));
 AO21x1_ASAP7_75t_R _26061_ (.A1(_07331_),
    .A2(_07333_),
    .B(_07121_),
    .Y(_07621_));
 AND3x1_ASAP7_75t_R _26062_ (.A(_07152_),
    .B(_07620_),
    .C(_07621_),
    .Y(_07622_));
 AO21x1_ASAP7_75t_R _26063_ (.A1(_07121_),
    .A2(_07423_),
    .B(_07224_),
    .Y(_07623_));
 AND2x2_ASAP7_75t_R _26064_ (.A(_07125_),
    .B(_07623_),
    .Y(_07624_));
 NAND2x2_ASAP7_75t_R _26065_ (.A(_07218_),
    .B(_07125_),
    .Y(_07625_));
 OA21x2_ASAP7_75t_R _26066_ (.A1(_07296_),
    .A2(_07300_),
    .B(_07121_),
    .Y(_07626_));
 AOI211x1_ASAP7_75t_R _26067_ (.A1(_07096_),
    .A2(_07314_),
    .B(_07317_),
    .C(_07121_),
    .Y(_07627_));
 AND3x1_ASAP7_75t_R _26068_ (.A(_07121_),
    .B(_07287_),
    .C(_07290_),
    .Y(_07628_));
 AND2x2_ASAP7_75t_R _26069_ (.A(_07090_),
    .B(_07308_),
    .Y(_07629_));
 OA33x2_ASAP7_75t_R _26070_ (.A1(_07625_),
    .A2(_07626_),
    .A3(_07627_),
    .B1(_07628_),
    .B2(_07629_),
    .B3(_07219_),
    .Y(_07630_));
 OA31x2_ASAP7_75t_R _26071_ (.A1(_07218_),
    .A2(_07622_),
    .A3(_07624_),
    .B1(_07630_),
    .Y(_07631_));
 NAND2x1_ASAP7_75t_R _26072_ (.A(_07215_),
    .B(_07631_),
    .Y(_07632_));
 TAPCELL_ASAP7_75t_R PHY_719 ();
 AND3x1_ASAP7_75t_R _26074_ (.A(_00086_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07634_));
 TAPCELL_ASAP7_75t_R PHY_718 ();
 AOI211x1_ASAP7_75t_R _26076_ (.A1(_00085_),
    .A2(_07238_),
    .B(_07634_),
    .C(_07234_),
    .Y(_07636_));
 AO21x1_ASAP7_75t_R _26077_ (.A1(_02365_),
    .A2(_07234_),
    .B(_07636_),
    .Y(_07637_));
 AOI22x1_ASAP7_75t_R _26078_ (.A1(net176),
    .A2(_07242_),
    .B1(_07637_),
    .B2(_07231_),
    .Y(_07638_));
 XNOR2x2_ASAP7_75t_R _26079_ (.A(_01387_),
    .B(_01385_),
    .Y(_07639_));
 INVx1_ASAP7_75t_R _26080_ (.A(_07639_),
    .Y(_07640_));
 AO221x1_ASAP7_75t_R _26081_ (.A1(_00670_),
    .A2(_07065_),
    .B1(_07640_),
    .B2(_07519_),
    .C(net308),
    .Y(_07641_));
 OA22x2_ASAP7_75t_R _26082_ (.A1(_01514_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01483_),
    .Y(_07642_));
 TAPCELL_ASAP7_75t_R PHY_717 ();
 OA22x2_ASAP7_75t_R _26084_ (.A1(_02167_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02061_),
    .Y(_07644_));
 OA22x2_ASAP7_75t_R _26085_ (.A1(_01990_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_00087_),
    .Y(_07645_));
 OR3x1_ASAP7_75t_R _26086_ (.A(_02024_),
    .B(_06990_),
    .C(_07023_),
    .Y(_07646_));
 OA211x2_ASAP7_75t_R _26087_ (.A1(_02093_),
    .A2(_07026_),
    .B(_07645_),
    .C(_07646_),
    .Y(_07647_));
 NAND2x1_ASAP7_75t_R _26088_ (.A(net3630),
    .B(_06947_),
    .Y(_07648_));
 OA21x2_ASAP7_75t_R _26089_ (.A1(_01940_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_07649_));
 OA211x2_ASAP7_75t_R _26090_ (.A1(_02134_),
    .A2(_07367_),
    .B(_07648_),
    .C(_07649_),
    .Y(_07650_));
 OA211x2_ASAP7_75t_R _26091_ (.A1(_07021_),
    .A2(_07644_),
    .B(_07647_),
    .C(_07650_),
    .Y(_07651_));
 OA21x2_ASAP7_75t_R _26092_ (.A1(_07360_),
    .A2(_07642_),
    .B(_07651_),
    .Y(_07652_));
 OA211x2_ASAP7_75t_R _26093_ (.A1(_13817_),
    .A2(_07638_),
    .B(_07641_),
    .C(_07652_),
    .Y(_07653_));
 AND4x2_ASAP7_75t_R _26094_ (.A(net290),
    .B(_07618_),
    .C(_07632_),
    .D(_07653_),
    .Y(_07654_));
 AO221x1_ASAP7_75t_R _26095_ (.A1(net40),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net31),
    .C(_07036_),
    .Y(_07655_));
 INVx1_ASAP7_75t_R _26096_ (.A(_01858_),
    .Y(_07656_));
 INVx1_ASAP7_75t_R _26097_ (.A(_01866_),
    .Y(_07657_));
 AO221x1_ASAP7_75t_R _26098_ (.A1(_07656_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07657_),
    .C(_07034_),
    .Y(_07658_));
 NOR2x1_ASAP7_75t_R _26099_ (.A(_01850_),
    .B(_07046_),
    .Y(_07659_));
 AO21x1_ASAP7_75t_R _26100_ (.A1(net48),
    .A2(_05762_),
    .B(_07659_),
    .Y(_07660_));
 AO222x2_ASAP7_75t_R _26101_ (.A1(net54),
    .A2(_07264_),
    .B1(_07655_),
    .B2(_07658_),
    .C1(_07660_),
    .C2(_07044_),
    .Y(_07661_));
 NOR2x1_ASAP7_75t_R _26102_ (.A(net290),
    .B(_07661_),
    .Y(_07662_));
 NOR2x2_ASAP7_75t_R _26103_ (.A(_07654_),
    .B(_07662_),
    .Y(_07663_));
 NOR2x1_ASAP7_75t_R _26104_ (.A(_01704_),
    .B(net288),
    .Y(_07664_));
 AO21x1_ASAP7_75t_R _26105_ (.A1(net288),
    .A2(_07663_),
    .B(_07664_),
    .Y(_02661_));
 AO221x1_ASAP7_75t_R _26106_ (.A1(net2563),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net2440),
    .C(_07036_),
    .Y(_07665_));
 INVx1_ASAP7_75t_R _26107_ (.A(_01857_),
    .Y(_07666_));
 INVx1_ASAP7_75t_R _26108_ (.A(_01865_),
    .Y(_07667_));
 AO221x1_ASAP7_75t_R _26109_ (.A1(_07666_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07667_),
    .C(_07034_),
    .Y(_07668_));
 INVx1_ASAP7_75t_R _26110_ (.A(net2419),
    .Y(_07669_));
 OAI22x1_ASAP7_75t_R _26111_ (.A1(_07669_),
    .A2(_01730_),
    .B1(_01849_),
    .B2(_07046_),
    .Y(_07670_));
 AO222x2_ASAP7_75t_R _26112_ (.A1(net3769),
    .A2(_07264_),
    .B1(_07665_),
    .B2(_07668_),
    .C1(_07670_),
    .C2(_07044_),
    .Y(_07671_));
 TAPCELL_ASAP7_75t_R PHY_716 ();
 OA21x2_ASAP7_75t_R _26114_ (.A1(_07387_),
    .A2(_07388_),
    .B(_07121_),
    .Y(_07673_));
 AO21x2_ASAP7_75t_R _26115_ (.A1(_07090_),
    .A2(_07401_),
    .B(_07673_),
    .Y(_07674_));
 OR2x2_ASAP7_75t_R _26116_ (.A(_07152_),
    .B(_07275_),
    .Y(_07675_));
 OA21x2_ASAP7_75t_R _26117_ (.A1(_07125_),
    .A2(_07674_),
    .B(_07675_),
    .Y(_07676_));
 NAND2x1_ASAP7_75t_R _26118_ (.A(_07121_),
    .B(_07413_),
    .Y(_07677_));
 OR3x1_ASAP7_75t_R _26119_ (.A(_07121_),
    .B(_07390_),
    .C(_07391_),
    .Y(_07678_));
 AND2x2_ASAP7_75t_R _26120_ (.A(_07677_),
    .B(_07678_),
    .Y(_07679_));
 NOR3x1_ASAP7_75t_R _26121_ (.A(_07090_),
    .B(_07407_),
    .C(_07408_),
    .Y(_07680_));
 AO21x1_ASAP7_75t_R _26122_ (.A1(_07090_),
    .A2(_07415_),
    .B(_07680_),
    .Y(_07681_));
 OA22x2_ASAP7_75t_R _26123_ (.A1(_07625_),
    .A2(_07679_),
    .B1(_07681_),
    .B2(_07219_),
    .Y(_07682_));
 OA211x2_ASAP7_75t_R _26124_ (.A1(_07218_),
    .A2(_07676_),
    .B(_07682_),
    .C(_07215_),
    .Y(_07683_));
 INVx1_ASAP7_75t_R _26125_ (.A(_02233_),
    .Y(_07684_));
 TAPCELL_ASAP7_75t_R PHY_715 ();
 AO32x1_ASAP7_75t_R _26127_ (.A1(_07684_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00672_),
    .Y(_07686_));
 NAND2x1_ASAP7_75t_R _26128_ (.A(_13817_),
    .B(_07686_),
    .Y(_07687_));
 AND3x1_ASAP7_75t_R _26129_ (.A(_00089_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07688_));
 AOI211x1_ASAP7_75t_R _26130_ (.A1(_00088_),
    .A2(_07238_),
    .B(_07688_),
    .C(_07234_),
    .Y(_07689_));
 AO21x1_ASAP7_75t_R _26131_ (.A1(_02366_),
    .A2(_07234_),
    .B(_07689_),
    .Y(_07690_));
 AO221x2_ASAP7_75t_R _26132_ (.A1(net177),
    .A2(_07242_),
    .B1(_07690_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07691_));
 AO32x1_ASAP7_75t_R _26133_ (.A1(_07077_),
    .A2(_07273_),
    .A3(_07340_),
    .B1(_07687_),
    .B2(_07691_),
    .Y(_07692_));
 OA22x2_ASAP7_75t_R _26134_ (.A1(_02166_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02060_),
    .Y(_07693_));
 OA22x2_ASAP7_75t_R _26135_ (.A1(_02092_),
    .A2(_07026_),
    .B1(_07369_),
    .B2(_00090_),
    .Y(_07694_));
 OA22x2_ASAP7_75t_R _26136_ (.A1(_01989_),
    .A2(_07024_),
    .B1(_07028_),
    .B2(_02023_),
    .Y(_07695_));
 TAPCELL_ASAP7_75t_R PHY_714 ();
 OA22x2_ASAP7_75t_R _26138_ (.A1(_01939_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02133_),
    .Y(_07697_));
 OA21x2_ASAP7_75t_R _26139_ (.A1(_01712_),
    .A2(_07000_),
    .B(_07004_),
    .Y(_07698_));
 AND4x1_ASAP7_75t_R _26140_ (.A(_14297_),
    .B(_14359_),
    .C(net310),
    .D(_05596_),
    .Y(_07699_));
 AND3x4_ASAP7_75t_R _26141_ (.A(_05586_),
    .B(_07699_),
    .C(_06945_),
    .Y(_07700_));
 TAPCELL_ASAP7_75t_R PHY_713 ();
 NAND2x2_ASAP7_75t_R _26143_ (.A(net3744),
    .B(_07700_),
    .Y(_07702_));
 AND5x2_ASAP7_75t_R _26144_ (.A(_07694_),
    .B(_07695_),
    .C(_07697_),
    .D(_07698_),
    .E(_07702_),
    .Y(_07703_));
 OAI22x1_ASAP7_75t_R _26145_ (.A1(_01513_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01482_),
    .Y(_07704_));
 NAND2x1_ASAP7_75t_R _26146_ (.A(_06950_),
    .B(_07704_),
    .Y(_07705_));
 OA211x2_ASAP7_75t_R _26147_ (.A1(_07021_),
    .A2(_07693_),
    .B(_07703_),
    .C(_07705_),
    .Y(_07706_));
 INVx1_ASAP7_75t_R _26148_ (.A(_07706_),
    .Y(_07707_));
 OR4x2_ASAP7_75t_R _26149_ (.A(_07474_),
    .B(_07683_),
    .C(_07692_),
    .D(_07707_),
    .Y(_07708_));
 OA21x2_ASAP7_75t_R _26150_ (.A1(net290),
    .A2(net3770),
    .B(_07708_),
    .Y(_07709_));
 NOR2x1_ASAP7_75t_R _26151_ (.A(_01703_),
    .B(net288),
    .Y(_07710_));
 AO21x1_ASAP7_75t_R _26152_ (.A1(net288),
    .A2(_07709_),
    .B(_07710_),
    .Y(_02662_));
 OA211x2_ASAP7_75t_R _26153_ (.A1(_07096_),
    .A2(_07488_),
    .B(_07489_),
    .C(_07121_),
    .Y(_07711_));
 AO31x2_ASAP7_75t_R _26154_ (.A1(_07090_),
    .A2(_07479_),
    .A3(_07482_),
    .B(_07711_),
    .Y(_07712_));
 OR2x2_ASAP7_75t_R _26155_ (.A(_07152_),
    .B(_07225_),
    .Y(_07713_));
 OA21x2_ASAP7_75t_R _26156_ (.A1(_07125_),
    .A2(_07712_),
    .B(_07713_),
    .Y(_07714_));
 AND2x2_ASAP7_75t_R _26157_ (.A(_07090_),
    .B(_07486_),
    .Y(_07715_));
 AO21x1_ASAP7_75t_R _26158_ (.A1(_07121_),
    .A2(_07496_),
    .B(_07715_),
    .Y(_07716_));
 AND3x1_ASAP7_75t_R _26159_ (.A(_07090_),
    .B(_07497_),
    .C(_07498_),
    .Y(_07717_));
 AO21x1_ASAP7_75t_R _26160_ (.A1(_07121_),
    .A2(_07503_),
    .B(_07717_),
    .Y(_07718_));
 OA222x2_ASAP7_75t_R _26161_ (.A1(_07218_),
    .A2(_07714_),
    .B1(_07716_),
    .B2(_07625_),
    .C1(_07718_),
    .C2(_07219_),
    .Y(_07719_));
 AND3x1_ASAP7_75t_R _26162_ (.A(_00092_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07720_));
 AOI211x1_ASAP7_75t_R _26163_ (.A1(_00091_),
    .A2(_07238_),
    .B(_07720_),
    .C(_07234_),
    .Y(_07721_));
 AO21x1_ASAP7_75t_R _26164_ (.A1(_02367_),
    .A2(_07234_),
    .B(_07721_),
    .Y(_07722_));
 AO22x1_ASAP7_75t_R _26165_ (.A1(net178),
    .A2(_07242_),
    .B1(_07722_),
    .B2(_07231_),
    .Y(_07723_));
 TAPCELL_ASAP7_75t_R PHY_712 ();
 TAPCELL_ASAP7_75t_R PHY_711 ();
 TAPCELL_ASAP7_75t_R PHY_710 ();
 XNOR2x1_ASAP7_75t_R _26169_ (.B(_02232_),
    .Y(_07727_),
    .A(net2335));
 AND2x2_ASAP7_75t_R _26170_ (.A(_07062_),
    .B(_07727_),
    .Y(_07728_));
 AO21x1_ASAP7_75t_R _26171_ (.A1(_00674_),
    .A2(_07064_),
    .B(_07728_),
    .Y(_07729_));
 AO21x1_ASAP7_75t_R _26172_ (.A1(_07060_),
    .A2(_07729_),
    .B(net308),
    .Y(_07730_));
 AOI21x1_ASAP7_75t_R _26173_ (.A1(_00674_),
    .A2(_07059_),
    .B(_07730_),
    .Y(_07731_));
 AO21x1_ASAP7_75t_R _26174_ (.A1(net308),
    .A2(_07723_),
    .B(_07731_),
    .Y(_07732_));
 NAND2x2_ASAP7_75t_R _26175_ (.A(_07105_),
    .B(_07123_),
    .Y(_07733_));
 AND3x1_ASAP7_75t_R _26176_ (.A(_07733_),
    .B(_07152_),
    .C(_07426_),
    .Y(_07734_));
 OAI22x1_ASAP7_75t_R _26177_ (.A1(_01512_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01481_),
    .Y(_07735_));
 NAND2x1_ASAP7_75t_R _26178_ (.A(_06950_),
    .B(_07735_),
    .Y(_07736_));
 OA21x2_ASAP7_75t_R _26179_ (.A1(_01938_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_07737_));
 OA22x2_ASAP7_75t_R _26180_ (.A1(_02091_),
    .A2(_07026_),
    .B1(_07522_),
    .B2(_01947_),
    .Y(_07738_));
 OA211x2_ASAP7_75t_R _26181_ (.A1(_02022_),
    .A2(_07028_),
    .B(_07737_),
    .C(_07738_),
    .Y(_07739_));
 OR3x4_ASAP7_75t_R _26182_ (.A(_06992_),
    .B(_07003_),
    .C(_07006_),
    .Y(_07740_));
 OA222x2_ASAP7_75t_R _26183_ (.A1(_01711_),
    .A2(_07000_),
    .B1(_07367_),
    .B2(_02132_),
    .C1(_07740_),
    .C2(_01454_),
    .Y(_07741_));
 NAND2x1_ASAP7_75t_R _26184_ (.A(net3613),
    .B(_06947_),
    .Y(_07742_));
 OA22x2_ASAP7_75t_R _26185_ (.A1(_02165_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02059_),
    .Y(_07743_));
 INVx1_ASAP7_75t_R _26186_ (.A(net3207),
    .Y(_07744_));
 NAND2x2_ASAP7_75t_R _26187_ (.A(_06942_),
    .B(_06965_),
    .Y(_07745_));
 OA222x2_ASAP7_75t_R _26188_ (.A1(_01988_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01574_),
    .C1(_07744_),
    .C2(_07745_),
    .Y(_07746_));
 OA21x2_ASAP7_75t_R _26189_ (.A1(_07021_),
    .A2(_07743_),
    .B(_07746_),
    .Y(_07747_));
 AND5x2_ASAP7_75t_R _26190_ (.A(_07736_),
    .B(_07739_),
    .C(_07741_),
    .D(net3614),
    .E(_07747_),
    .Y(_07748_));
 INVx1_ASAP7_75t_R _26191_ (.A(_07748_),
    .Y(_07749_));
 OR3x1_ASAP7_75t_R _26192_ (.A(_07732_),
    .B(_07734_),
    .C(_07749_),
    .Y(_07750_));
 AOI21x1_ASAP7_75t_R _26193_ (.A1(_07215_),
    .A2(_07719_),
    .B(_07750_),
    .Y(_07751_));
 AO221x1_ASAP7_75t_R _26194_ (.A1(net2566),
    .A2(_07041_),
    .B1(_07253_),
    .B2(net2569),
    .C(_07036_),
    .Y(_07752_));
 INVx1_ASAP7_75t_R _26195_ (.A(_01856_),
    .Y(_07753_));
 INVx1_ASAP7_75t_R _26196_ (.A(_01864_),
    .Y(_07754_));
 AO221x1_ASAP7_75t_R _26197_ (.A1(_07753_),
    .A2(_07041_),
    .B1(_07253_),
    .B2(_07754_),
    .C(_07034_),
    .Y(_07755_));
 INVx1_ASAP7_75t_R _26198_ (.A(net2510),
    .Y(_07756_));
 OAI22x1_ASAP7_75t_R _26199_ (.A1(_07756_),
    .A2(_01730_),
    .B1(_01733_),
    .B2(_07046_),
    .Y(_07757_));
 AO222x2_ASAP7_75t_R _26200_ (.A1(net3763),
    .A2(_07264_),
    .B1(_07752_),
    .B2(_07755_),
    .C1(_07757_),
    .C2(_07044_),
    .Y(_07758_));
 NOR2x2_ASAP7_75t_R _26201_ (.A(net290),
    .B(net3764),
    .Y(_07759_));
 AOI21x1_ASAP7_75t_R _26202_ (.A1(_06981_),
    .A2(_07751_),
    .B(_07759_),
    .Y(_07760_));
 TAPCELL_ASAP7_75t_R PHY_709 ();
 NOR2x1_ASAP7_75t_R _26204_ (.A(_01702_),
    .B(_06987_),
    .Y(_07762_));
 AO21x1_ASAP7_75t_R _26205_ (.A1(_06987_),
    .A2(net252),
    .B(_07762_),
    .Y(_02663_));
 INVx1_ASAP7_75t_R _26206_ (.A(_02235_),
    .Y(_07763_));
 TAPCELL_ASAP7_75t_R PHY_708 ();
 AO32x1_ASAP7_75t_R _26208_ (.A1(_07763_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00677_),
    .Y(_07765_));
 AND2x2_ASAP7_75t_R _26209_ (.A(_07125_),
    .B(_07223_),
    .Y(_07766_));
 INVx1_ASAP7_75t_R _26210_ (.A(_07766_),
    .Y(_07767_));
 OAI21x1_ASAP7_75t_R _26211_ (.A1(_07105_),
    .A2(_07125_),
    .B(_07767_),
    .Y(_07768_));
 AND2x2_ASAP7_75t_R _26212_ (.A(_07073_),
    .B(_07121_),
    .Y(_07769_));
 OR2x2_ASAP7_75t_R _26213_ (.A(_07113_),
    .B(_07120_),
    .Y(_07770_));
 AO22x1_ASAP7_75t_R _26214_ (.A1(_07218_),
    .A2(_07178_),
    .B1(_07769_),
    .B2(_07770_),
    .Y(_07771_));
 OR3x1_ASAP7_75t_R _26215_ (.A(_07137_),
    .B(_07144_),
    .C(_07151_),
    .Y(_07772_));
 NOR2x1_ASAP7_75t_R _26216_ (.A(_07772_),
    .B(_07625_),
    .Y(_07773_));
 AO221x2_ASAP7_75t_R _26217_ (.A1(_07073_),
    .A2(_07768_),
    .B1(_07771_),
    .B2(_07152_),
    .C(_07773_),
    .Y(_07774_));
 AND3x1_ASAP7_75t_R _26218_ (.A(_00094_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07775_));
 AOI211x1_ASAP7_75t_R _26219_ (.A1(_00093_),
    .A2(_07238_),
    .B(_07775_),
    .C(_07234_),
    .Y(_07776_));
 AO21x1_ASAP7_75t_R _26220_ (.A1(_02368_),
    .A2(_07234_),
    .B(_07776_),
    .Y(_07777_));
 AO221x2_ASAP7_75t_R _26221_ (.A1(net179),
    .A2(_07242_),
    .B1(_07777_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07778_));
 AOI221x1_ASAP7_75t_R _26222_ (.A1(_07426_),
    .A2(_07714_),
    .B1(_07774_),
    .B2(_07215_),
    .C(_07778_),
    .Y(_07779_));
 AO21x1_ASAP7_75t_R _26223_ (.A1(_13817_),
    .A2(_07765_),
    .B(_07779_),
    .Y(_07780_));
 TAPCELL_ASAP7_75t_R PHY_707 ();
 TAPCELL_ASAP7_75t_R PHY_706 ();
 TAPCELL_ASAP7_75t_R PHY_705 ();
 OA22x2_ASAP7_75t_R _26227_ (.A1(_01511_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01480_),
    .Y(_07784_));
 OA22x2_ASAP7_75t_R _26228_ (.A1(_02164_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02058_),
    .Y(_07785_));
 TAPCELL_ASAP7_75t_R PHY_704 ();
 TAPCELL_ASAP7_75t_R PHY_703 ();
 OA222x2_ASAP7_75t_R _26231_ (.A1(_01987_),
    .A2(_07024_),
    .B1(_07028_),
    .B2(_02021_),
    .C1(_07008_),
    .C2(_00095_),
    .Y(_07788_));
 OA21x2_ASAP7_75t_R _26232_ (.A1(_07021_),
    .A2(_07785_),
    .B(_07788_),
    .Y(_07789_));
 OA21x2_ASAP7_75t_R _26233_ (.A1(_14359_),
    .A2(_05693_),
    .B(_06955_),
    .Y(_07790_));
 NAND2x2_ASAP7_75t_R _26234_ (.A(_07790_),
    .B(_06957_),
    .Y(_07791_));
 TAPCELL_ASAP7_75t_R PHY_702 ();
 OA222x2_ASAP7_75t_R _26236_ (.A1(_01937_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02131_),
    .C1(_07000_),
    .C2(_01726_),
    .Y(_07793_));
 OA22x2_ASAP7_75t_R _26237_ (.A1(_02090_),
    .A2(_07026_),
    .B1(_07369_),
    .B2(_01573_),
    .Y(_07794_));
 NAND2x1_ASAP7_75t_R _26238_ (.A(net3723),
    .B(_06947_),
    .Y(_07795_));
 AND4x1_ASAP7_75t_R _26239_ (.A(_07791_),
    .B(_07793_),
    .C(_07794_),
    .D(net3724),
    .Y(_07796_));
 OA211x2_ASAP7_75t_R _26240_ (.A1(_07360_),
    .A2(_07784_),
    .B(_07789_),
    .C(_07796_),
    .Y(_07797_));
 AND2x2_ASAP7_75t_R _26241_ (.A(_06981_),
    .B(_07797_),
    .Y(_07798_));
 TAPCELL_ASAP7_75t_R PHY_701 ();
 TAPCELL_ASAP7_75t_R PHY_700 ();
 TAPCELL_ASAP7_75t_R PHY_699 ();
 TAPCELL_ASAP7_75t_R PHY_698 ();
 NOR2x1_ASAP7_75t_R _26246_ (.A(net3780),
    .B(net433),
    .Y(_07803_));
 AOI21x1_ASAP7_75t_R _26247_ (.A1(_07045_),
    .A2(net433),
    .B(_07803_),
    .Y(_07804_));
 TAPCELL_ASAP7_75t_R PHY_697 ();
 TAPCELL_ASAP7_75t_R PHY_696 ();
 OR2x2_ASAP7_75t_R _26250_ (.A(net57),
    .B(_07051_),
    .Y(_07807_));
 TAPCELL_ASAP7_75t_R PHY_695 ();
 OA211x2_ASAP7_75t_R _26252_ (.A1(net2494),
    .A2(net433),
    .B(_07807_),
    .C(net432),
    .Y(_07809_));
 AOI21x1_ASAP7_75t_R _26253_ (.A1(_07039_),
    .A2(_07804_),
    .B(_07809_),
    .Y(_07810_));
 TAPCELL_ASAP7_75t_R PHY_694 ();
 AOI211x1_ASAP7_75t_R _26255_ (.A1(net433),
    .A2(_01855_),
    .B(_07803_),
    .C(net432),
    .Y(_07812_));
 OA211x2_ASAP7_75t_R _26256_ (.A1(net433),
    .A2(_07035_),
    .B(_07807_),
    .C(net432),
    .Y(_07813_));
 TAPCELL_ASAP7_75t_R PHY_693 ();
 OAI21x1_ASAP7_75t_R _26258_ (.A1(_07812_),
    .A2(_07813_),
    .B(_07036_),
    .Y(_07815_));
 INVx1_ASAP7_75t_R _26259_ (.A(_01644_),
    .Y(_07816_));
 AND2x2_ASAP7_75t_R _26260_ (.A(net56),
    .B(net434),
    .Y(_07817_));
 AO21x1_ASAP7_75t_R _26261_ (.A1(net33),
    .A2(_07051_),
    .B(_07817_),
    .Y(_07818_));
 OR2x2_ASAP7_75t_R _26262_ (.A(net42),
    .B(_07051_),
    .Y(_07819_));
 OA211x2_ASAP7_75t_R _26263_ (.A1(net51),
    .A2(net434),
    .B(_07819_),
    .C(_07039_),
    .Y(_07820_));
 AO21x1_ASAP7_75t_R _26264_ (.A1(net432),
    .A2(_07818_),
    .B(_07820_),
    .Y(_07821_));
 AND3x2_ASAP7_75t_R _26265_ (.A(_07816_),
    .B(_05762_),
    .C(_07821_),
    .Y(_07822_));
 NOR2x2_ASAP7_75t_R _26266_ (.A(net290),
    .B(_07822_),
    .Y(_07823_));
 OA211x2_ASAP7_75t_R _26267_ (.A1(_01731_),
    .A2(_07810_),
    .B(_07815_),
    .C(_07823_),
    .Y(_07824_));
 AOI21x1_ASAP7_75t_R _26268_ (.A1(_07780_),
    .A2(_07798_),
    .B(_07824_),
    .Y(_07825_));
 NOR2x1_ASAP7_75t_R _26269_ (.A(_01701_),
    .B(net288),
    .Y(_07826_));
 AO21x1_ASAP7_75t_R _26270_ (.A1(net288),
    .A2(net257),
    .B(_07826_),
    .Y(_02664_));
 TAPCELL_ASAP7_75t_R PHY_692 ();
 AO21x1_ASAP7_75t_R _26272_ (.A1(_07152_),
    .A2(_07340_),
    .B(_07766_),
    .Y(_07828_));
 OR2x2_ASAP7_75t_R _26273_ (.A(_07301_),
    .B(_07309_),
    .Y(_07829_));
 OR3x1_ASAP7_75t_R _26274_ (.A(_07152_),
    .B(_07318_),
    .C(_07325_),
    .Y(_07830_));
 OA211x2_ASAP7_75t_R _26275_ (.A1(_07125_),
    .A2(_07829_),
    .B(_07830_),
    .C(_07218_),
    .Y(_07831_));
 AO21x1_ASAP7_75t_R _26276_ (.A1(_07073_),
    .A2(_07828_),
    .B(_07831_),
    .Y(_07832_));
 NAND2x1_ASAP7_75t_R _26277_ (.A(_07215_),
    .B(_07832_),
    .Y(_07833_));
 AND2x2_ASAP7_75t_R _26278_ (.A(_07073_),
    .B(_07223_),
    .Y(_07834_));
 AO221x1_ASAP7_75t_R _26279_ (.A1(_07275_),
    .A2(_07310_),
    .B1(_07674_),
    .B2(_07273_),
    .C(_07834_),
    .Y(_07835_));
 NAND2x1_ASAP7_75t_R _26280_ (.A(_07077_),
    .B(_07835_),
    .Y(_07836_));
 XOR2x2_ASAP7_75t_R _26281_ (.A(_01426_),
    .B(_02234_),
    .Y(_07837_));
 AO21x1_ASAP7_75t_R _26282_ (.A1(_00279_),
    .A2(_07062_),
    .B(_15282_),
    .Y(_07838_));
 OA21x2_ASAP7_75t_R _26283_ (.A1(_07267_),
    .A2(_07837_),
    .B(_07838_),
    .Y(_07839_));
 AND3x1_ASAP7_75t_R _26284_ (.A(_00097_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07840_));
 AOI211x1_ASAP7_75t_R _26285_ (.A1(_00096_),
    .A2(_07238_),
    .B(_07840_),
    .C(_07234_),
    .Y(_07841_));
 AO21x1_ASAP7_75t_R _26286_ (.A1(_02369_),
    .A2(_07234_),
    .B(_07841_),
    .Y(_07842_));
 AO221x2_ASAP7_75t_R _26287_ (.A1(net2200),
    .A2(_07242_),
    .B1(_07842_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07843_));
 OAI21x1_ASAP7_75t_R _26288_ (.A1(net308),
    .A2(_07839_),
    .B(_07843_),
    .Y(_07844_));
 OA22x2_ASAP7_75t_R _26289_ (.A1(_01510_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01479_),
    .Y(_07845_));
 OA22x2_ASAP7_75t_R _26290_ (.A1(_02163_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02057_),
    .Y(_07846_));
 OA222x2_ASAP7_75t_R _26291_ (.A1(_00098_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01572_),
    .C1(_01986_),
    .C2(_07024_),
    .Y(_07847_));
 OA21x2_ASAP7_75t_R _26292_ (.A1(_07021_),
    .A2(_07846_),
    .B(_07847_),
    .Y(_07848_));
 OA33x2_ASAP7_75t_R _26293_ (.A1(_02089_),
    .A2(_05589_),
    .A3(_06994_),
    .B1(_07023_),
    .B2(_06990_),
    .B3(_02020_),
    .Y(_07849_));
 OA22x2_ASAP7_75t_R _26294_ (.A1(_01936_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02130_),
    .Y(_07850_));
 NAND2x1_ASAP7_75t_R _26295_ (.A(net3714),
    .B(_07700_),
    .Y(_07851_));
 AND4x1_ASAP7_75t_R _26296_ (.A(_07004_),
    .B(_07849_),
    .C(_07850_),
    .D(net3715),
    .Y(_07852_));
 OA211x2_ASAP7_75t_R _26297_ (.A1(_07360_),
    .A2(_07845_),
    .B(_07848_),
    .C(_07852_),
    .Y(_07853_));
 AND4x1_ASAP7_75t_R _26298_ (.A(_06981_),
    .B(_07836_),
    .C(_07844_),
    .D(_07853_),
    .Y(_07854_));
 NOR2x1_ASAP7_75t_R _26299_ (.A(net38),
    .B(net434),
    .Y(_07855_));
 AO21x1_ASAP7_75t_R _26300_ (.A1(_07261_),
    .A2(net434),
    .B(_07855_),
    .Y(_07856_));
 OR2x2_ASAP7_75t_R _26301_ (.A(net58),
    .B(_07051_),
    .Y(_07857_));
 OA21x2_ASAP7_75t_R _26302_ (.A1(net35),
    .A2(net434),
    .B(_07857_),
    .Y(_07858_));
 NAND2x1_ASAP7_75t_R _26303_ (.A(net432),
    .B(_07858_),
    .Y(_07859_));
 OA21x2_ASAP7_75t_R _26304_ (.A1(net432),
    .A2(_07856_),
    .B(_07859_),
    .Y(_07860_));
 AOI211x1_ASAP7_75t_R _26305_ (.A1(net434),
    .A2(_01854_),
    .B(_07855_),
    .C(net432),
    .Y(_07861_));
 TAPCELL_ASAP7_75t_R PHY_691 ();
 OA211x2_ASAP7_75t_R _26307_ (.A1(net434),
    .A2(_07257_),
    .B(_07857_),
    .C(net432),
    .Y(_07863_));
 OAI21x1_ASAP7_75t_R _26308_ (.A1(_07861_),
    .A2(_07863_),
    .B(_07036_),
    .Y(_07864_));
 OA211x2_ASAP7_75t_R _26309_ (.A1(_01731_),
    .A2(_07860_),
    .B(_07864_),
    .C(_07823_),
    .Y(_07865_));
 AOI21x1_ASAP7_75t_R _26310_ (.A1(_07833_),
    .A2(_07854_),
    .B(_07865_),
    .Y(_07866_));
 NOR2x1_ASAP7_75t_R _26311_ (.A(_01700_),
    .B(_06987_),
    .Y(_07867_));
 AO21x1_ASAP7_75t_R _26312_ (.A1(_06987_),
    .A2(net256),
    .B(_07867_),
    .Y(_02665_));
 INVx1_ASAP7_75t_R _26313_ (.A(_02237_),
    .Y(_07868_));
 OAI21x1_ASAP7_75t_R _26314_ (.A1(_07868_),
    .A2(_07065_),
    .B(_00682_),
    .Y(_07869_));
 OA21x2_ASAP7_75t_R _26315_ (.A1(_02237_),
    .A2(_07520_),
    .B(_07869_),
    .Y(_07870_));
 AND3x1_ASAP7_75t_R _26316_ (.A(_00100_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07871_));
 AOI211x1_ASAP7_75t_R _26317_ (.A1(_00099_),
    .A2(_07238_),
    .B(_07871_),
    .C(_07234_),
    .Y(_07872_));
 AO21x1_ASAP7_75t_R _26318_ (.A1(_02370_),
    .A2(_07234_),
    .B(_07872_),
    .Y(_07873_));
 AO221x2_ASAP7_75t_R _26319_ (.A1(net151),
    .A2(_07242_),
    .B1(_07873_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07874_));
 OA21x2_ASAP7_75t_R _26320_ (.A1(net308),
    .A2(_07870_),
    .B(_07874_),
    .Y(_07875_));
 OA22x2_ASAP7_75t_R _26321_ (.A1(_01509_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01478_),
    .Y(_07876_));
 OA22x2_ASAP7_75t_R _26322_ (.A1(_02162_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02056_),
    .Y(_07877_));
 OA222x2_ASAP7_75t_R _26323_ (.A1(_00101_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01571_),
    .C1(_01985_),
    .C2(_07024_),
    .Y(_07878_));
 OA21x2_ASAP7_75t_R _26324_ (.A1(_07021_),
    .A2(_07877_),
    .B(_07878_),
    .Y(_07879_));
 OA33x2_ASAP7_75t_R _26325_ (.A1(_02088_),
    .A2(_05589_),
    .A3(_06994_),
    .B1(_07023_),
    .B2(_06990_),
    .B3(_02019_),
    .Y(_07880_));
 OA22x2_ASAP7_75t_R _26326_ (.A1(_01935_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02129_),
    .Y(_07881_));
 NAND2x1_ASAP7_75t_R _26327_ (.A(net3734),
    .B(_07700_),
    .Y(_07882_));
 AND4x1_ASAP7_75t_R _26328_ (.A(_07004_),
    .B(_07880_),
    .C(_07881_),
    .D(net3735),
    .Y(_07883_));
 OA211x2_ASAP7_75t_R _26329_ (.A1(_07360_),
    .A2(_07876_),
    .B(_07879_),
    .C(_07883_),
    .Y(_07884_));
 INVx1_ASAP7_75t_R _26330_ (.A(_07884_),
    .Y(_07885_));
 OR2x2_ASAP7_75t_R _26331_ (.A(_07622_),
    .B(_07624_),
    .Y(_07886_));
 AO21x1_ASAP7_75t_R _26332_ (.A1(_07426_),
    .A2(_07886_),
    .B(_07474_),
    .Y(_07887_));
 AOI22x1_ASAP7_75t_R _26333_ (.A1(_07310_),
    .A2(_07393_),
    .B1(_07417_),
    .B2(_07273_),
    .Y(_07888_));
 OA211x2_ASAP7_75t_R _26334_ (.A1(_07218_),
    .A2(_07617_),
    .B(_07888_),
    .C(_07215_),
    .Y(_07889_));
 OR4x2_ASAP7_75t_R _26335_ (.A(_07875_),
    .B(_07885_),
    .C(_07887_),
    .D(_07889_),
    .Y(_07890_));
 NOR2x1_ASAP7_75t_R _26336_ (.A(net49),
    .B(net433),
    .Y(_07891_));
 AO21x1_ASAP7_75t_R _26337_ (.A1(net433),
    .A2(_01853_),
    .B(_07891_),
    .Y(_07892_));
 OR2x2_ASAP7_75t_R _26338_ (.A(net28),
    .B(_07051_),
    .Y(_07893_));
 OA211x2_ASAP7_75t_R _26339_ (.A1(net433),
    .A2(_07465_),
    .B(_07893_),
    .C(net432),
    .Y(_07894_));
 INVx1_ASAP7_75t_R _26340_ (.A(_07894_),
    .Y(_07895_));
 OA21x2_ASAP7_75t_R _26341_ (.A1(net432),
    .A2(_07892_),
    .B(_07895_),
    .Y(_07896_));
 AO21x1_ASAP7_75t_R _26342_ (.A1(_07468_),
    .A2(net433),
    .B(_07891_),
    .Y(_07897_));
 OA211x2_ASAP7_75t_R _26343_ (.A1(net36),
    .A2(net433),
    .B(_07893_),
    .C(net432),
    .Y(_07898_));
 INVx1_ASAP7_75t_R _26344_ (.A(_07898_),
    .Y(_07899_));
 OA21x2_ASAP7_75t_R _26345_ (.A1(net432),
    .A2(_07897_),
    .B(_07899_),
    .Y(_07900_));
 OAI22x1_ASAP7_75t_R _26346_ (.A1(_07034_),
    .A2(_07896_),
    .B1(_07900_),
    .B2(_01731_),
    .Y(_07901_));
 OR3x1_ASAP7_75t_R _26347_ (.A(net290),
    .B(_07822_),
    .C(_07901_),
    .Y(_07902_));
 AND2x6_ASAP7_75t_R _26348_ (.A(_07890_),
    .B(_07902_),
    .Y(_07903_));
 NOR2x1_ASAP7_75t_R _26349_ (.A(_01699_),
    .B(net288),
    .Y(_07904_));
 AO21x1_ASAP7_75t_R _26350_ (.A1(net288),
    .A2(_07903_),
    .B(_07904_),
    .Y(_02666_));
 AO21x1_ASAP7_75t_R _26351_ (.A1(_07152_),
    .A2(_07484_),
    .B(_07766_),
    .Y(_07905_));
 AO22x1_ASAP7_75t_R _26352_ (.A1(_07273_),
    .A2(_07500_),
    .B1(_07905_),
    .B2(_07073_),
    .Y(_07906_));
 XOR2x2_ASAP7_75t_R _26353_ (.A(_01436_),
    .B(_02236_),
    .Y(_07907_));
 NOR2x1_ASAP7_75t_R _26354_ (.A(_07064_),
    .B(_07907_),
    .Y(_07908_));
 AO21x1_ASAP7_75t_R _26355_ (.A1(_00684_),
    .A2(_07064_),
    .B(_07908_),
    .Y(_07909_));
 AND2x2_ASAP7_75t_R _26356_ (.A(_07060_),
    .B(_07909_),
    .Y(_07910_));
 AOI21x1_ASAP7_75t_R _26357_ (.A1(_00684_),
    .A2(_07059_),
    .B(_07910_),
    .Y(_07911_));
 AND3x1_ASAP7_75t_R _26358_ (.A(_00103_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07912_));
 AOI211x1_ASAP7_75t_R _26359_ (.A1(_00102_),
    .A2(_07238_),
    .B(_07912_),
    .C(_07234_),
    .Y(_07913_));
 AO21x1_ASAP7_75t_R _26360_ (.A1(_02371_),
    .A2(_07234_),
    .B(_07913_),
    .Y(_07914_));
 AO221x2_ASAP7_75t_R _26361_ (.A1(net152),
    .A2(_07242_),
    .B1(_07914_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07915_));
 OA21x2_ASAP7_75t_R _26362_ (.A1(net308),
    .A2(_07911_),
    .B(_07915_),
    .Y(_07916_));
 OA211x2_ASAP7_75t_R _26363_ (.A1(_07487_),
    .A2(_07490_),
    .B(_07215_),
    .C(_07310_),
    .Y(_07917_));
 OR3x1_ASAP7_75t_R _26364_ (.A(_07474_),
    .B(_07916_),
    .C(_07917_),
    .Y(_07918_));
 NAND2x1_ASAP7_75t_R _26365_ (.A(_07426_),
    .B(_07571_),
    .Y(_07919_));
 TAPCELL_ASAP7_75t_R PHY_690 ();
 OA22x2_ASAP7_75t_R _26367_ (.A1(_01508_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01477_),
    .Y(_07921_));
 OA22x2_ASAP7_75t_R _26368_ (.A1(_02161_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02055_),
    .Y(_07922_));
 OA22x2_ASAP7_75t_R _26369_ (.A1(_02018_),
    .A2(_07028_),
    .B1(_07745_),
    .B2(net3369),
    .Y(_07923_));
 OA22x2_ASAP7_75t_R _26370_ (.A1(_00657_),
    .A2(_07008_),
    .B1(_07522_),
    .B2(_01948_),
    .Y(_07924_));
 OA211x2_ASAP7_75t_R _26371_ (.A1(_07021_),
    .A2(_07922_),
    .B(_07923_),
    .C(_07924_),
    .Y(_07925_));
 OA22x2_ASAP7_75t_R _26372_ (.A1(_01984_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01570_),
    .Y(_07926_));
 OA222x2_ASAP7_75t_R _26373_ (.A1(_02033_),
    .A2(_07000_),
    .B1(_07367_),
    .B2(_02128_),
    .C1(_07740_),
    .C2(_01456_),
    .Y(_07927_));
 NAND2x1_ASAP7_75t_R _26374_ (.A(_14180_),
    .B(_14238_),
    .Y(_07928_));
 OR4x2_ASAP7_75t_R _26375_ (.A(_13523_),
    .B(_13894_),
    .C(_05563_),
    .D(_07928_),
    .Y(_07929_));
 TAPCELL_ASAP7_75t_R PHY_689 ();
 OR3x1_ASAP7_75t_R _26377_ (.A(_02087_),
    .B(_05589_),
    .C(_07929_),
    .Y(_07931_));
 OA21x2_ASAP7_75t_R _26378_ (.A1(_01934_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_07932_));
 NAND2x2_ASAP7_75t_R _26379_ (.A(net3701),
    .B(_06947_),
    .Y(_07933_));
 AND5x2_ASAP7_75t_R _26380_ (.A(_07926_),
    .B(_07927_),
    .C(_07931_),
    .D(_07932_),
    .E(net3702),
    .Y(_07934_));
 OA211x2_ASAP7_75t_R _26381_ (.A1(_07360_),
    .A2(_07921_),
    .B(_07925_),
    .C(_07934_),
    .Y(_07935_));
 NAND2x1_ASAP7_75t_R _26382_ (.A(_07919_),
    .B(_07935_),
    .Y(_07936_));
 AOI211x1_ASAP7_75t_R _26383_ (.A1(_07215_),
    .A2(_07906_),
    .B(_07918_),
    .C(_07936_),
    .Y(_07937_));
 NOR2x1_ASAP7_75t_R _26384_ (.A(net52),
    .B(net434),
    .Y(_07938_));
 AOI21x1_ASAP7_75t_R _26385_ (.A1(_07548_),
    .A2(net434),
    .B(_07938_),
    .Y(_07939_));
 OR2x2_ASAP7_75t_R _26386_ (.A(net29),
    .B(_07051_),
    .Y(_07940_));
 OA211x2_ASAP7_75t_R _26387_ (.A1(net37),
    .A2(net434),
    .B(_07940_),
    .C(_01642_),
    .Y(_07941_));
 AOI21x1_ASAP7_75t_R _26388_ (.A1(_07039_),
    .A2(_07939_),
    .B(_07941_),
    .Y(_07942_));
 AOI211x1_ASAP7_75t_R _26389_ (.A1(net434),
    .A2(_01852_),
    .B(_07938_),
    .C(_01642_),
    .Y(_07943_));
 TAPCELL_ASAP7_75t_R PHY_688 ();
 OA211x2_ASAP7_75t_R _26391_ (.A1(net434),
    .A2(_07545_),
    .B(_07940_),
    .C(_01642_),
    .Y(_07945_));
 OAI21x1_ASAP7_75t_R _26392_ (.A1(_07943_),
    .A2(_07945_),
    .B(_07036_),
    .Y(_07946_));
 OA211x2_ASAP7_75t_R _26393_ (.A1(_01731_),
    .A2(_07942_),
    .B(_07946_),
    .C(_07823_),
    .Y(_07947_));
 NOR2x2_ASAP7_75t_R _26394_ (.A(_07937_),
    .B(_07947_),
    .Y(_07948_));
 NOR2x1_ASAP7_75t_R _26395_ (.A(_01698_),
    .B(net288),
    .Y(_07949_));
 AO21x1_ASAP7_75t_R _26396_ (.A1(net288),
    .A2(_07948_),
    .B(_07949_),
    .Y(_02667_));
 NOR2x1_ASAP7_75t_R _26397_ (.A(net53),
    .B(net433),
    .Y(_07950_));
 AO21x1_ASAP7_75t_R _26398_ (.A1(net433),
    .A2(_01851_),
    .B(_07950_),
    .Y(_07951_));
 INVx1_ASAP7_75t_R _26399_ (.A(net30),
    .Y(_07952_));
 NAND2x1_ASAP7_75t_R _26400_ (.A(_07952_),
    .B(net433),
    .Y(_07953_));
 OA211x2_ASAP7_75t_R _26401_ (.A1(net433),
    .A2(_07601_),
    .B(_07953_),
    .C(net432),
    .Y(_07954_));
 INVx1_ASAP7_75t_R _26402_ (.A(_07954_),
    .Y(_07955_));
 OA21x2_ASAP7_75t_R _26403_ (.A1(net432),
    .A2(_07951_),
    .B(_07955_),
    .Y(_07956_));
 AOI21x1_ASAP7_75t_R _26404_ (.A1(_07604_),
    .A2(net433),
    .B(_07950_),
    .Y(_07957_));
 OA211x2_ASAP7_75t_R _26405_ (.A1(net39),
    .A2(net433),
    .B(_07953_),
    .C(net432),
    .Y(_07958_));
 AOI21x1_ASAP7_75t_R _26406_ (.A1(_07039_),
    .A2(_07957_),
    .B(_07958_),
    .Y(_07959_));
 OAI22x1_ASAP7_75t_R _26407_ (.A1(_07034_),
    .A2(_07956_),
    .B1(_07959_),
    .B2(_01731_),
    .Y(_07960_));
 OR3x4_ASAP7_75t_R _26408_ (.A(net290),
    .B(_07822_),
    .C(_07960_),
    .Y(_07961_));
 AND3x1_ASAP7_75t_R _26409_ (.A(_07215_),
    .B(_07218_),
    .C(_07125_),
    .Y(_07962_));
 INVx1_ASAP7_75t_R _26410_ (.A(_02239_),
    .Y(_07963_));
 AO32x1_ASAP7_75t_R _26411_ (.A1(_07963_),
    .A2(_07060_),
    .A3(_07062_),
    .B1(_07065_),
    .B2(_00686_),
    .Y(_07964_));
 NAND2x1_ASAP7_75t_R _26412_ (.A(_13817_),
    .B(_07964_),
    .Y(_07965_));
 AND3x1_ASAP7_75t_R _26413_ (.A(_00105_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07966_));
 AOI211x1_ASAP7_75t_R _26414_ (.A1(_00104_),
    .A2(_07238_),
    .B(_07966_),
    .C(_07234_),
    .Y(_07967_));
 AO21x1_ASAP7_75t_R _26415_ (.A1(_02372_),
    .A2(_07234_),
    .B(_07967_),
    .Y(_07968_));
 AO221x2_ASAP7_75t_R _26416_ (.A1(net153),
    .A2(_07242_),
    .B1(_07968_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_07969_));
 AO222x2_ASAP7_75t_R _26417_ (.A1(_07426_),
    .A2(_07493_),
    .B1(_07568_),
    .B2(_07962_),
    .C1(_07965_),
    .C2(_07969_),
    .Y(_07970_));
 AO22x1_ASAP7_75t_R _26418_ (.A1(_07073_),
    .A2(_07513_),
    .B1(_07577_),
    .B2(_07273_),
    .Y(_07971_));
 OAI22x1_ASAP7_75t_R _26419_ (.A1(_01507_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01476_),
    .Y(_07972_));
 OA22x2_ASAP7_75t_R _26420_ (.A1(_02160_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02054_),
    .Y(_07973_));
 OA222x2_ASAP7_75t_R _26421_ (.A1(_00656_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01569_),
    .C1(_02017_),
    .C2(_07028_),
    .Y(_07974_));
 OAI21x1_ASAP7_75t_R _26422_ (.A1(_07021_),
    .A2(_07973_),
    .B(_07974_),
    .Y(_07975_));
 OAI22x1_ASAP7_75t_R _26423_ (.A1(_01933_),
    .A2(_06998_),
    .B1(_07000_),
    .B2(_02032_),
    .Y(_07976_));
 OAI22x1_ASAP7_75t_R _26424_ (.A1(_02127_),
    .A2(_07367_),
    .B1(_07740_),
    .B2(_01455_),
    .Y(_07977_));
 OA22x2_ASAP7_75t_R _26425_ (.A1(_02086_),
    .A2(_06994_),
    .B1(_07023_),
    .B2(_01983_),
    .Y(_07978_));
 NOR2x1_ASAP7_75t_R _26426_ (.A(_05589_),
    .B(_07978_),
    .Y(_07979_));
 AO21x1_ASAP7_75t_R _26427_ (.A1(net3671),
    .A2(_06947_),
    .B(_06958_),
    .Y(_07980_));
 OR5x2_ASAP7_75t_R _26428_ (.A(_07975_),
    .B(_07976_),
    .C(_07977_),
    .D(_07979_),
    .E(net3672),
    .Y(_07981_));
 AO21x2_ASAP7_75t_R _26429_ (.A1(_06950_),
    .A2(_07972_),
    .B(_07981_),
    .Y(_07982_));
 AO21x1_ASAP7_75t_R _26430_ (.A1(_07215_),
    .A2(_07971_),
    .B(_07982_),
    .Y(_07983_));
 OR3x4_ASAP7_75t_R _26431_ (.A(_07474_),
    .B(_07970_),
    .C(_07983_),
    .Y(_07984_));
 AND2x6_ASAP7_75t_R _26432_ (.A(_07961_),
    .B(_07984_),
    .Y(_07985_));
 NOR2x1_ASAP7_75t_R _26433_ (.A(_01697_),
    .B(net288),
    .Y(_07986_));
 AO21x1_ASAP7_75t_R _26434_ (.A1(net288),
    .A2(_07985_),
    .B(_07986_),
    .Y(_02668_));
 OR2x2_ASAP7_75t_R _26435_ (.A(_07626_),
    .B(_07627_),
    .Y(_07987_));
 AO21x1_ASAP7_75t_R _26436_ (.A1(_07620_),
    .A2(_07621_),
    .B(_07152_),
    .Y(_07988_));
 OA211x2_ASAP7_75t_R _26437_ (.A1(_07125_),
    .A2(_07987_),
    .B(_07988_),
    .C(_07218_),
    .Y(_07989_));
 AO21x1_ASAP7_75t_R _26438_ (.A1(_07073_),
    .A2(_07425_),
    .B(_07989_),
    .Y(_07990_));
 NAND2x1_ASAP7_75t_R _26439_ (.A(_07215_),
    .B(_07990_),
    .Y(_07991_));
 AO21x1_ASAP7_75t_R _26440_ (.A1(_07121_),
    .A2(_07401_),
    .B(_07403_),
    .Y(_07992_));
 AND3x1_ASAP7_75t_R _26441_ (.A(_07152_),
    .B(_07389_),
    .C(_07392_),
    .Y(_07993_));
 AO21x1_ASAP7_75t_R _26442_ (.A1(_07125_),
    .A2(_07992_),
    .B(_07993_),
    .Y(_07994_));
 XNOR2x2_ASAP7_75t_R _26443_ (.A(net2146),
    .B(_02238_),
    .Y(_07995_));
 AO32x1_ASAP7_75t_R _26444_ (.A1(_07060_),
    .A2(_07062_),
    .A3(_07995_),
    .B1(_07065_),
    .B2(_00718_),
    .Y(_07996_));
 NAND2x1_ASAP7_75t_R _26445_ (.A(_13817_),
    .B(_07996_),
    .Y(_07997_));
 AND3x1_ASAP7_75t_R _26446_ (.A(_00107_),
    .B(_13618_),
    .C(_06635_),
    .Y(_07998_));
 AOI211x1_ASAP7_75t_R _26447_ (.A1(_00106_),
    .A2(_07238_),
    .B(_07998_),
    .C(_07234_),
    .Y(_07999_));
 AO21x1_ASAP7_75t_R _26448_ (.A1(_02373_),
    .A2(_07234_),
    .B(_07999_),
    .Y(_08000_));
 AO221x2_ASAP7_75t_R _26449_ (.A1(net154),
    .A2(_07242_),
    .B1(_08000_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08001_));
 AO21x1_ASAP7_75t_R _26450_ (.A1(_07997_),
    .A2(_08001_),
    .B(_07474_),
    .Y(_08002_));
 OA22x2_ASAP7_75t_R _26451_ (.A1(_01506_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01475_),
    .Y(_08003_));
 OA33x2_ASAP7_75t_R _26452_ (.A1(_01568_),
    .A2(_05589_),
    .A3(_06938_),
    .B1(_06990_),
    .B2(_07023_),
    .B3(_02016_),
    .Y(_08004_));
 OA22x2_ASAP7_75t_R _26453_ (.A1(_01932_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02126_),
    .Y(_08005_));
 OA21x2_ASAP7_75t_R _26454_ (.A1(_02031_),
    .A2(_07000_),
    .B(_07004_),
    .Y(_08006_));
 NAND2x1_ASAP7_75t_R _26455_ (.A(net3706),
    .B(_06947_),
    .Y(_08007_));
 AND4x2_ASAP7_75t_R _26456_ (.A(_08004_),
    .B(_08005_),
    .C(_08006_),
    .D(_08007_),
    .Y(_08008_));
 OA22x2_ASAP7_75t_R _26457_ (.A1(_02159_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02053_),
    .Y(_08009_));
 OA222x2_ASAP7_75t_R _26458_ (.A1(_01982_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02085_),
    .C1(_07008_),
    .C2(_00108_),
    .Y(_08010_));
 OA21x2_ASAP7_75t_R _26459_ (.A1(_07021_),
    .A2(_08009_),
    .B(_08010_),
    .Y(_08011_));
 OA211x2_ASAP7_75t_R _26460_ (.A1(_07360_),
    .A2(_08003_),
    .B(_08008_),
    .C(_08011_),
    .Y(_08012_));
 INVx1_ASAP7_75t_R _26461_ (.A(_08012_),
    .Y(_08013_));
 AOI211x1_ASAP7_75t_R _26462_ (.A1(_07994_),
    .A2(_07426_),
    .B(_08002_),
    .C(_08013_),
    .Y(_08014_));
 OR2x2_ASAP7_75t_R _26463_ (.A(net31),
    .B(_07051_),
    .Y(_08015_));
 OAI21x1_ASAP7_75t_R _26464_ (.A1(net2482),
    .A2(net433),
    .B(_08015_),
    .Y(_08016_));
 OR2x2_ASAP7_75t_R _26465_ (.A(net54),
    .B(net433),
    .Y(_08017_));
 OA21x2_ASAP7_75t_R _26466_ (.A1(net2476),
    .A2(_07051_),
    .B(_08017_),
    .Y(_08018_));
 NOR2x1_ASAP7_75t_R _26467_ (.A(net432),
    .B(_08018_),
    .Y(_08019_));
 AO21x1_ASAP7_75t_R _26468_ (.A1(net432),
    .A2(_08016_),
    .B(_08019_),
    .Y(_08020_));
 INVx1_ASAP7_75t_R _26469_ (.A(_01850_),
    .Y(_08021_));
 OA211x2_ASAP7_75t_R _26470_ (.A1(_07051_),
    .A2(_08021_),
    .B(_08017_),
    .C(_07039_),
    .Y(_08022_));
 OA211x2_ASAP7_75t_R _26471_ (.A1(net433),
    .A2(_07656_),
    .B(_08015_),
    .C(net432),
    .Y(_08023_));
 OAI21x1_ASAP7_75t_R _26472_ (.A1(_08022_),
    .A2(_08023_),
    .B(_07036_),
    .Y(_08024_));
 OA211x2_ASAP7_75t_R _26473_ (.A1(_01731_),
    .A2(_08020_),
    .B(_08024_),
    .C(_07823_),
    .Y(_08025_));
 AOI21x1_ASAP7_75t_R _26474_ (.A1(_07991_),
    .A2(_08014_),
    .B(_08025_),
    .Y(_08026_));
 NOR2x1_ASAP7_75t_R _26475_ (.A(_01696_),
    .B(_06987_),
    .Y(_08027_));
 AO21x1_ASAP7_75t_R _26476_ (.A1(_06987_),
    .A2(net251),
    .B(_08027_),
    .Y(_02669_));
 NOR2x1_ASAP7_75t_R _26477_ (.A(net55),
    .B(net433),
    .Y(_08028_));
 AOI21x1_ASAP7_75t_R _26478_ (.A1(_07669_),
    .A2(net434),
    .B(_08028_),
    .Y(_08029_));
 INVx1_ASAP7_75t_R _26479_ (.A(net32),
    .Y(_08030_));
 NAND2x1_ASAP7_75t_R _26480_ (.A(_08030_),
    .B(net434),
    .Y(_08031_));
 OA211x2_ASAP7_75t_R _26481_ (.A1(net41),
    .A2(net434),
    .B(_08031_),
    .C(net432),
    .Y(_08032_));
 AOI21x1_ASAP7_75t_R _26482_ (.A1(_07039_),
    .A2(_08029_),
    .B(_08032_),
    .Y(_08033_));
 AOI211x1_ASAP7_75t_R _26483_ (.A1(net434),
    .A2(_01849_),
    .B(_08028_),
    .C(net432),
    .Y(_08034_));
 OA211x2_ASAP7_75t_R _26484_ (.A1(net434),
    .A2(_07666_),
    .B(_08031_),
    .C(net432),
    .Y(_08035_));
 OAI21x1_ASAP7_75t_R _26485_ (.A1(_08034_),
    .A2(_08035_),
    .B(_07036_),
    .Y(_08036_));
 OA211x2_ASAP7_75t_R _26486_ (.A1(_01731_),
    .A2(_08033_),
    .B(_08036_),
    .C(_07823_),
    .Y(_08037_));
 AND2x2_ASAP7_75t_R _26487_ (.A(_07152_),
    .B(_07679_),
    .Y(_08038_));
 OR2x2_ASAP7_75t_R _26488_ (.A(_07152_),
    .B(_07223_),
    .Y(_08039_));
 OA211x2_ASAP7_75t_R _26489_ (.A1(_07125_),
    .A2(_07275_),
    .B(_08039_),
    .C(_07073_),
    .Y(_08040_));
 AO21x1_ASAP7_75t_R _26490_ (.A1(_07218_),
    .A2(_08038_),
    .B(_08040_),
    .Y(_08041_));
 OR3x1_ASAP7_75t_R _26491_ (.A(_07125_),
    .B(_07318_),
    .C(_07325_),
    .Y(_08042_));
 OA211x2_ASAP7_75t_R _26492_ (.A1(_07152_),
    .A2(_07340_),
    .B(_08042_),
    .C(_07426_),
    .Y(_08043_));
 INVx1_ASAP7_75t_R _26493_ (.A(_02241_),
    .Y(_08044_));
 AND3x1_ASAP7_75t_R _26494_ (.A(_00279_),
    .B(_08044_),
    .C(_07062_),
    .Y(_08045_));
 AOI21x1_ASAP7_75t_R _26495_ (.A1(_00750_),
    .A2(_07267_),
    .B(_08045_),
    .Y(_08046_));
 AND3x1_ASAP7_75t_R _26496_ (.A(_00110_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08047_));
 AOI211x1_ASAP7_75t_R _26497_ (.A1(_00109_),
    .A2(_07238_),
    .B(_08047_),
    .C(_07234_),
    .Y(_08048_));
 AO21x1_ASAP7_75t_R _26498_ (.A1(_02374_),
    .A2(_07234_),
    .B(_08048_),
    .Y(_08049_));
 AO221x1_ASAP7_75t_R _26499_ (.A1(net155),
    .A2(_07242_),
    .B1(_08049_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08050_));
 OA21x2_ASAP7_75t_R _26500_ (.A1(net308),
    .A2(_08046_),
    .B(_08050_),
    .Y(_08051_));
 AO21x1_ASAP7_75t_R _26501_ (.A1(_07674_),
    .A2(_07962_),
    .B(_08051_),
    .Y(_08052_));
 OAI22x1_ASAP7_75t_R _26502_ (.A1(_01505_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01474_),
    .Y(_08053_));
 AND2x2_ASAP7_75t_R _26503_ (.A(_06950_),
    .B(_08053_),
    .Y(_08054_));
 OAI22x1_ASAP7_75t_R _26504_ (.A1(_02158_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02052_),
    .Y(_08055_));
 AND2x2_ASAP7_75t_R _26505_ (.A(_06940_),
    .B(_08055_),
    .Y(_08056_));
 AND3x2_ASAP7_75t_R _26506_ (.A(_14358_),
    .B(_05693_),
    .C(_06957_),
    .Y(_08057_));
 OAI22x1_ASAP7_75t_R _26507_ (.A1(_02084_),
    .A2(_07026_),
    .B1(_07028_),
    .B2(_02015_),
    .Y(_08058_));
 NOR2x1_ASAP7_75t_R _26508_ (.A(_02125_),
    .B(_07367_),
    .Y(_08059_));
 NOR2x1_ASAP7_75t_R _26509_ (.A(_01931_),
    .B(_06998_),
    .Y(_08060_));
 OR4x2_ASAP7_75t_R _26510_ (.A(_08057_),
    .B(_08058_),
    .C(_08059_),
    .D(_08060_),
    .Y(_08061_));
 AO21x1_ASAP7_75t_R _26511_ (.A1(net3586),
    .A2(_06947_),
    .B(_08061_),
    .Y(_08062_));
 OA222x2_ASAP7_75t_R _26512_ (.A1(_00111_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01567_),
    .C1(_01981_),
    .C2(_07024_),
    .Y(_08063_));
 INVx1_ASAP7_75t_R _26513_ (.A(_08063_),
    .Y(_08064_));
 OR4x2_ASAP7_75t_R _26514_ (.A(_08054_),
    .B(_08056_),
    .C(_08062_),
    .D(_08064_),
    .Y(_08065_));
 OR4x1_ASAP7_75t_R _26515_ (.A(_07474_),
    .B(_08043_),
    .C(_08052_),
    .D(_08065_),
    .Y(_08066_));
 AOI21x1_ASAP7_75t_R _26516_ (.A1(_07215_),
    .A2(_08041_),
    .B(_08066_),
    .Y(_08067_));
 NOR2x2_ASAP7_75t_R _26517_ (.A(_08037_),
    .B(_08067_),
    .Y(_08068_));
 NOR2x1_ASAP7_75t_R _26518_ (.A(_01695_),
    .B(net288),
    .Y(_08069_));
 AO21x1_ASAP7_75t_R _26519_ (.A1(net288),
    .A2(_08068_),
    .B(_08069_),
    .Y(_02670_));
 NOR2x1_ASAP7_75t_R _26520_ (.A(net56),
    .B(net434),
    .Y(_08070_));
 AO21x1_ASAP7_75t_R _26521_ (.A1(net434),
    .A2(_01733_),
    .B(_08070_),
    .Y(_08071_));
 OR2x2_ASAP7_75t_R _26522_ (.A(net33),
    .B(_07051_),
    .Y(_08072_));
 OA211x2_ASAP7_75t_R _26523_ (.A1(net434),
    .A2(_07753_),
    .B(_08072_),
    .C(_01642_),
    .Y(_08073_));
 INVx1_ASAP7_75t_R _26524_ (.A(_08073_),
    .Y(_08074_));
 OA21x2_ASAP7_75t_R _26525_ (.A1(_01642_),
    .A2(_08071_),
    .B(_08074_),
    .Y(_08075_));
 OA21x2_ASAP7_75t_R _26526_ (.A1(net42),
    .A2(net434),
    .B(_08072_),
    .Y(_08076_));
 AO21x1_ASAP7_75t_R _26527_ (.A1(_07756_),
    .A2(net434),
    .B(_08070_),
    .Y(_08077_));
 NOR2x1_ASAP7_75t_R _26528_ (.A(_01642_),
    .B(_08077_),
    .Y(_08078_));
 AO21x1_ASAP7_75t_R _26529_ (.A1(_01642_),
    .A2(_08076_),
    .B(_08078_),
    .Y(_08079_));
 NAND2x1_ASAP7_75t_R _26530_ (.A(_05750_),
    .B(_08079_),
    .Y(_08080_));
 OA211x2_ASAP7_75t_R _26531_ (.A1(_07034_),
    .A2(_08075_),
    .B(_08080_),
    .C(_07823_),
    .Y(_08081_));
 OA21x2_ASAP7_75t_R _26532_ (.A1(_07125_),
    .A2(_07225_),
    .B(_08039_),
    .Y(_08082_));
 OA222x2_ASAP7_75t_R _26533_ (.A1(_07625_),
    .A2(_07712_),
    .B1(_07716_),
    .B2(_07219_),
    .C1(_07218_),
    .C2(_08082_),
    .Y(_08083_));
 NAND2x1_ASAP7_75t_R _26534_ (.A(_07215_),
    .B(_08083_),
    .Y(_08084_));
 AND3x1_ASAP7_75t_R _26535_ (.A(_00113_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08085_));
 AOI211x1_ASAP7_75t_R _26536_ (.A1(_00112_),
    .A2(_07238_),
    .B(_08085_),
    .C(_07234_),
    .Y(_08086_));
 AO21x1_ASAP7_75t_R _26537_ (.A1(_02375_),
    .A2(_07234_),
    .B(_08086_),
    .Y(_08087_));
 AOI22x1_ASAP7_75t_R _26538_ (.A1(net156),
    .A2(_07242_),
    .B1(_08087_),
    .B2(_07231_),
    .Y(_08088_));
 XOR2x1_ASAP7_75t_R _26539_ (.A(net2237),
    .Y(_08089_),
    .B(_02240_));
 NOR2x1_ASAP7_75t_R _26540_ (.A(_07064_),
    .B(_08089_),
    .Y(_08090_));
 AO21x1_ASAP7_75t_R _26541_ (.A1(_00783_),
    .A2(_07064_),
    .B(_08090_),
    .Y(_08091_));
 AO221x1_ASAP7_75t_R _26542_ (.A1(_00783_),
    .A2(_07059_),
    .B1(_07060_),
    .B2(_08091_),
    .C(net308),
    .Y(_08092_));
 OAI22x1_ASAP7_75t_R _26543_ (.A1(_02157_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02051_),
    .Y(_08093_));
 OAI22x1_ASAP7_75t_R _26544_ (.A1(_01504_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01473_),
    .Y(_08094_));
 OAI22x1_ASAP7_75t_R _26545_ (.A1(_01566_),
    .A2(_05589_),
    .B1(_07447_),
    .B2(_01930_),
    .Y(_08095_));
 AO32x1_ASAP7_75t_R _26546_ (.A1(net302),
    .A2(_05604_),
    .A3(_05693_),
    .B1(_07440_),
    .B2(_08095_),
    .Y(_08096_));
 INVx2_ASAP7_75t_R _26547_ (.A(_00114_),
    .Y(_08097_));
 INVx1_ASAP7_75t_R _26548_ (.A(_07007_),
    .Y(_08098_));
 OAI22x1_ASAP7_75t_R _26549_ (.A1(_02030_),
    .A2(_05589_),
    .B1(_07447_),
    .B2(_02124_),
    .Y(_08099_));
 AO32x1_ASAP7_75t_R _26550_ (.A1(_08097_),
    .A2(_08098_),
    .A3(_07450_),
    .B1(_08099_),
    .B2(_05693_),
    .Y(_08100_));
 AND2x2_ASAP7_75t_R _26551_ (.A(net3746),
    .B(_07443_),
    .Y(_08101_));
 OR2x2_ASAP7_75t_R _26552_ (.A(_07447_),
    .B(_07023_),
    .Y(_08102_));
 OA222x2_ASAP7_75t_R _26553_ (.A1(_01980_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02083_),
    .C1(_08102_),
    .C2(_02014_),
    .Y(_08103_));
 INVx1_ASAP7_75t_R _26554_ (.A(_08103_),
    .Y(_08104_));
 OR4x1_ASAP7_75t_R _26555_ (.A(_08096_),
    .B(_08100_),
    .C(_08101_),
    .D(_08104_),
    .Y(_08105_));
 AOI221x1_ASAP7_75t_R _26556_ (.A1(_07441_),
    .A2(_08093_),
    .B1(_08094_),
    .B2(_07438_),
    .C(_08105_),
    .Y(_08106_));
 OA211x2_ASAP7_75t_R _26557_ (.A1(_13817_),
    .A2(_08088_),
    .B(_08092_),
    .C(_08106_),
    .Y(_08107_));
 OR3x1_ASAP7_75t_R _26558_ (.A(_07073_),
    .B(_07080_),
    .C(_07154_),
    .Y(_08108_));
 AND4x2_ASAP7_75t_R _26559_ (.A(net290),
    .B(_08084_),
    .C(_08107_),
    .D(_08108_),
    .Y(_08109_));
 NOR2x2_ASAP7_75t_R _26560_ (.A(_08081_),
    .B(_08109_),
    .Y(_08110_));
 NOR2x1_ASAP7_75t_R _26561_ (.A(_01694_),
    .B(_06987_),
    .Y(_08111_));
 AO21x1_ASAP7_75t_R _26562_ (.A1(_06987_),
    .A2(_08110_),
    .B(_08111_),
    .Y(_02671_));
 NOR2x1_ASAP7_75t_R _26563_ (.A(_01644_),
    .B(_08080_),
    .Y(_08112_));
 OR3x4_ASAP7_75t_R _26564_ (.A(net290),
    .B(_07822_),
    .C(_08112_),
    .Y(_08113_));
 TAPCELL_ASAP7_75t_R PHY_687 ();
 TAPCELL_ASAP7_75t_R PHY_686 ();
 AO21x1_ASAP7_75t_R _26567_ (.A1(net57),
    .A2(_07051_),
    .B(_07049_),
    .Y(_08116_));
 NAND2x1_ASAP7_75t_R _26568_ (.A(net34),
    .B(net433),
    .Y(_08117_));
 OA211x2_ASAP7_75t_R _26569_ (.A1(net433),
    .A2(_01855_),
    .B(_08117_),
    .C(net432),
    .Y(_08118_));
 INVx1_ASAP7_75t_R _26570_ (.A(_08118_),
    .Y(_08119_));
 TAPCELL_ASAP7_75t_R PHY_685 ();
 OA211x2_ASAP7_75t_R _26572_ (.A1(net432),
    .A2(_08116_),
    .B(_08119_),
    .C(_07036_),
    .Y(_08121_));
 AND3x1_ASAP7_75t_R _26573_ (.A(_00116_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08122_));
 AOI211x1_ASAP7_75t_R _26574_ (.A1(_00115_),
    .A2(_07238_),
    .B(_08122_),
    .C(_07234_),
    .Y(_08123_));
 AO21x1_ASAP7_75t_R _26575_ (.A1(_02376_),
    .A2(_07234_),
    .B(_08123_),
    .Y(_08124_));
 AOI22x1_ASAP7_75t_R _26576_ (.A1(net157),
    .A2(_07242_),
    .B1(_08124_),
    .B2(_07231_),
    .Y(_08125_));
 AND2x2_ASAP7_75t_R _26577_ (.A(_01356_),
    .B(_07064_),
    .Y(_08126_));
 AO21x1_ASAP7_75t_R _26578_ (.A1(_00030_),
    .A2(_07062_),
    .B(_08126_),
    .Y(_08127_));
 AO221x1_ASAP7_75t_R _26579_ (.A1(_00816_),
    .A2(_07059_),
    .B1(_07060_),
    .B2(_08127_),
    .C(net308),
    .Y(_08128_));
 OA21x2_ASAP7_75t_R _26580_ (.A1(_13817_),
    .A2(_08125_),
    .B(_08128_),
    .Y(_08129_));
 OA22x2_ASAP7_75t_R _26581_ (.A1(_01503_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01472_),
    .Y(_08130_));
 OA22x2_ASAP7_75t_R _26582_ (.A1(_02156_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02050_),
    .Y(_08131_));
 OA222x2_ASAP7_75t_R _26583_ (.A1(_00117_),
    .A2(_07008_),
    .B1(_07522_),
    .B2(_01963_),
    .C1(_02013_),
    .C2(_07028_),
    .Y(_08132_));
 OA21x2_ASAP7_75t_R _26584_ (.A1(_07021_),
    .A2(_08131_),
    .B(_08132_),
    .Y(_08133_));
 AND2x4_ASAP7_75t_R _26585_ (.A(_06942_),
    .B(_06965_),
    .Y(_08134_));
 NAND2x1_ASAP7_75t_R _26586_ (.A(net3299),
    .B(_08134_),
    .Y(_08135_));
 OA22x2_ASAP7_75t_R _26587_ (.A1(_01979_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01565_),
    .Y(_08136_));
 OA211x2_ASAP7_75t_R _26588_ (.A1(_02082_),
    .A2(_07026_),
    .B(_08135_),
    .C(_08136_),
    .Y(_08137_));
 NAND2x1_ASAP7_75t_R _26589_ (.A(net3602),
    .B(_06947_),
    .Y(_08138_));
 OA21x2_ASAP7_75t_R _26590_ (.A1(_02123_),
    .A2(_07367_),
    .B(_07004_),
    .Y(_08139_));
 OA21x2_ASAP7_75t_R _26591_ (.A1(_01929_),
    .A2(_06998_),
    .B(_08139_),
    .Y(_08140_));
 AND4x1_ASAP7_75t_R _26592_ (.A(_08133_),
    .B(_08137_),
    .C(net3603),
    .D(_08140_),
    .Y(_08141_));
 OA21x2_ASAP7_75t_R _26593_ (.A1(_07360_),
    .A2(_08130_),
    .B(_08141_),
    .Y(_08142_));
 NAND2x1_ASAP7_75t_R _26594_ (.A(_08129_),
    .B(_08142_),
    .Y(_08143_));
 NOR2x1_ASAP7_75t_R _26595_ (.A(_07216_),
    .B(_07154_),
    .Y(_08144_));
 AND3x1_ASAP7_75t_R _26596_ (.A(_07073_),
    .B(_07077_),
    .C(_08082_),
    .Y(_08145_));
 AO21x1_ASAP7_75t_R _26597_ (.A1(_07218_),
    .A2(_08144_),
    .B(_08145_),
    .Y(_08146_));
 OR2x2_ASAP7_75t_R _26598_ (.A(_07474_),
    .B(_07834_),
    .Y(_08147_));
 OR2x2_ASAP7_75t_R _26599_ (.A(_07152_),
    .B(_07712_),
    .Y(_08148_));
 OA211x2_ASAP7_75t_R _26600_ (.A1(_07125_),
    .A2(_07716_),
    .B(_08148_),
    .C(_07426_),
    .Y(_08149_));
 OR4x1_ASAP7_75t_R _26601_ (.A(_08143_),
    .B(_08146_),
    .C(_08147_),
    .D(_08149_),
    .Y(_08150_));
 OA21x2_ASAP7_75t_R _26602_ (.A1(_08113_),
    .A2(_08121_),
    .B(_08150_),
    .Y(_08151_));
 NOR2x1_ASAP7_75t_R _26603_ (.A(_01693_),
    .B(net288),
    .Y(_08152_));
 AO21x1_ASAP7_75t_R _26604_ (.A1(net288),
    .A2(_08151_),
    .B(_08152_),
    .Y(_02672_));
 AND2x2_ASAP7_75t_R _26605_ (.A(net38),
    .B(net434),
    .Y(_08153_));
 AO21x1_ASAP7_75t_R _26606_ (.A1(net58),
    .A2(_07051_),
    .B(_08153_),
    .Y(_08154_));
 NAND2x1_ASAP7_75t_R _26607_ (.A(net35),
    .B(net434),
    .Y(_08155_));
 OA211x2_ASAP7_75t_R _26608_ (.A1(net434),
    .A2(_01854_),
    .B(_08155_),
    .C(net432),
    .Y(_08156_));
 INVx1_ASAP7_75t_R _26609_ (.A(_08156_),
    .Y(_08157_));
 OA211x2_ASAP7_75t_R _26610_ (.A1(net432),
    .A2(_08154_),
    .B(_08157_),
    .C(_07036_),
    .Y(_08158_));
 AND3x1_ASAP7_75t_R _26611_ (.A(_07218_),
    .B(_07125_),
    .C(_07674_),
    .Y(_08159_));
 OA21x2_ASAP7_75t_R _26612_ (.A1(_08040_),
    .A2(_08159_),
    .B(_07077_),
    .Y(_08160_));
 OAI22x1_ASAP7_75t_R _26613_ (.A1(_01502_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01471_),
    .Y(_08161_));
 NAND2x1_ASAP7_75t_R _26614_ (.A(_06950_),
    .B(_08161_),
    .Y(_08162_));
 OR3x1_ASAP7_75t_R _26615_ (.A(_01978_),
    .B(_05589_),
    .C(_07023_),
    .Y(_08163_));
 OA33x2_ASAP7_75t_R _26616_ (.A1(_01564_),
    .A2(_05589_),
    .A3(_06938_),
    .B1(_06990_),
    .B2(_07023_),
    .B3(_02012_),
    .Y(_08164_));
 OA211x2_ASAP7_75t_R _26617_ (.A1(_01962_),
    .A2(_07522_),
    .B(_08163_),
    .C(_08164_),
    .Y(_08165_));
 OA22x2_ASAP7_75t_R _26618_ (.A1(_02122_),
    .A2(_07367_),
    .B1(_07740_),
    .B2(_01996_),
    .Y(_08166_));
 OA211x2_ASAP7_75t_R _26619_ (.A1(_01928_),
    .A2(_06998_),
    .B(_07004_),
    .C(_08166_),
    .Y(_08167_));
 NAND2x1_ASAP7_75t_R _26620_ (.A(net3658),
    .B(_06947_),
    .Y(_08168_));
 OA22x2_ASAP7_75t_R _26621_ (.A1(_02155_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02049_),
    .Y(_08169_));
 INVx1_ASAP7_75t_R _26622_ (.A(net3665),
    .Y(_08170_));
 OA222x2_ASAP7_75t_R _26623_ (.A1(_02081_),
    .A2(_07026_),
    .B1(_07008_),
    .B2(_00120_),
    .C1(net3666),
    .C2(_07745_),
    .Y(_08171_));
 OA21x2_ASAP7_75t_R _26624_ (.A1(_07021_),
    .A2(_08169_),
    .B(_08171_),
    .Y(_08172_));
 AND5x2_ASAP7_75t_R _26625_ (.A(_08162_),
    .B(_08165_),
    .C(_08167_),
    .D(net3659),
    .E(_08172_),
    .Y(_08173_));
 INVx1_ASAP7_75t_R _26626_ (.A(_08173_),
    .Y(_08174_));
 AND3x1_ASAP7_75t_R _26627_ (.A(_07215_),
    .B(_07218_),
    .C(_07152_),
    .Y(_08175_));
 OR2x2_ASAP7_75t_R _26628_ (.A(_07318_),
    .B(_07325_),
    .Y(_08176_));
 AND3x1_ASAP7_75t_R _26629_ (.A(_00119_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08177_));
 AOI211x1_ASAP7_75t_R _26630_ (.A1(_00118_),
    .A2(_07238_),
    .B(_08177_),
    .C(_07234_),
    .Y(_08178_));
 AO21x1_ASAP7_75t_R _26631_ (.A1(_02377_),
    .A2(_07234_),
    .B(_08178_),
    .Y(_08179_));
 AO221x1_ASAP7_75t_R _26632_ (.A1(net2254),
    .A2(_07242_),
    .B1(_08179_),
    .B2(_07231_),
    .C(_07834_),
    .Y(_08180_));
 XOR2x1_ASAP7_75t_R _26633_ (.A(_00033_),
    .Y(_08181_),
    .B(net2196));
 AND2x2_ASAP7_75t_R _26634_ (.A(_07062_),
    .B(_08181_),
    .Y(_08182_));
 AO21x1_ASAP7_75t_R _26635_ (.A1(_01360_),
    .A2(_07064_),
    .B(_08182_),
    .Y(_08183_));
 AO21x1_ASAP7_75t_R _26636_ (.A1(_07060_),
    .A2(_08183_),
    .B(net308),
    .Y(_08184_));
 AOI21x1_ASAP7_75t_R _26637_ (.A1(_00849_),
    .A2(_07059_),
    .B(_08184_),
    .Y(_08185_));
 AO21x1_ASAP7_75t_R _26638_ (.A1(net308),
    .A2(_08180_),
    .B(_08185_),
    .Y(_08186_));
 AO221x1_ASAP7_75t_R _26639_ (.A1(_07340_),
    .A2(_07962_),
    .B1(_08175_),
    .B2(_08176_),
    .C(_08186_),
    .Y(_08187_));
 AO21x1_ASAP7_75t_R _26640_ (.A1(_07426_),
    .A2(_08038_),
    .B(_08187_),
    .Y(_08188_));
 OR4x2_ASAP7_75t_R _26641_ (.A(_07474_),
    .B(_08160_),
    .C(_08174_),
    .D(_08188_),
    .Y(_08189_));
 OA21x2_ASAP7_75t_R _26642_ (.A1(_08113_),
    .A2(_08158_),
    .B(_08189_),
    .Y(_08190_));
 TAPCELL_ASAP7_75t_R PHY_684 ();
 NOR2x1_ASAP7_75t_R _26644_ (.A(_01692_),
    .B(net288),
    .Y(_08192_));
 AO21x1_ASAP7_75t_R _26645_ (.A1(net288),
    .A2(_08190_),
    .B(_08192_),
    .Y(_02673_));
 AND2x2_ASAP7_75t_R _26646_ (.A(net49),
    .B(net433),
    .Y(_08193_));
 AO21x1_ASAP7_75t_R _26647_ (.A1(net28),
    .A2(_07051_),
    .B(_08193_),
    .Y(_08194_));
 NAND2x1_ASAP7_75t_R _26648_ (.A(net36),
    .B(net433),
    .Y(_08195_));
 OA211x2_ASAP7_75t_R _26649_ (.A1(net433),
    .A2(_01853_),
    .B(_08195_),
    .C(net432),
    .Y(_08196_));
 INVx1_ASAP7_75t_R _26650_ (.A(_08196_),
    .Y(_08197_));
 OA211x2_ASAP7_75t_R _26651_ (.A1(net432),
    .A2(_08194_),
    .B(_08197_),
    .C(_07036_),
    .Y(_08198_));
 AND3x1_ASAP7_75t_R _26652_ (.A(_00122_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08199_));
 AOI211x1_ASAP7_75t_R _26653_ (.A1(_00121_),
    .A2(_07238_),
    .B(_08199_),
    .C(_07234_),
    .Y(_08200_));
 AO21x1_ASAP7_75t_R _26654_ (.A1(_02378_),
    .A2(_07234_),
    .B(_08200_),
    .Y(_08201_));
 AO22x2_ASAP7_75t_R _26655_ (.A1(net159),
    .A2(_07242_),
    .B1(_08201_),
    .B2(_07231_),
    .Y(_08202_));
 OR2x2_ASAP7_75t_R _26656_ (.A(_07073_),
    .B(_08202_),
    .Y(_08203_));
 OA21x2_ASAP7_75t_R _26657_ (.A1(_07218_),
    .A2(_07223_),
    .B(_07215_),
    .Y(_08204_));
 OA21x2_ASAP7_75t_R _26658_ (.A1(_08202_),
    .A2(_08204_),
    .B(net308),
    .Y(_08205_));
 OA21x2_ASAP7_75t_R _26659_ (.A1(_07994_),
    .A2(_08203_),
    .B(_08205_),
    .Y(_08206_));
 NOR2x1_ASAP7_75t_R _26660_ (.A(_02243_),
    .B(_07064_),
    .Y(_08207_));
 AO21x1_ASAP7_75t_R _26661_ (.A1(_01364_),
    .A2(_07064_),
    .B(_08207_),
    .Y(_08208_));
 AO21x1_ASAP7_75t_R _26662_ (.A1(_07060_),
    .A2(_08208_),
    .B(net308),
    .Y(_08209_));
 AOI21x1_ASAP7_75t_R _26663_ (.A1(_00881_),
    .A2(_07059_),
    .B(_08209_),
    .Y(_08210_));
 OAI22x1_ASAP7_75t_R _26664_ (.A1(_01501_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01470_),
    .Y(_08211_));
 AND2x2_ASAP7_75t_R _26665_ (.A(_06950_),
    .B(_08211_),
    .Y(_08212_));
 AND2x2_ASAP7_75t_R _26666_ (.A(_06956_),
    .B(_06960_),
    .Y(_08213_));
 AO32x1_ASAP7_75t_R _26667_ (.A1(_06246_),
    .A2(_06942_),
    .A3(_08213_),
    .B1(_08134_),
    .B2(net3555),
    .Y(_08214_));
 OAI22x1_ASAP7_75t_R _26668_ (.A1(_00123_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01563_),
    .Y(_08215_));
 OA21x2_ASAP7_75t_R _26669_ (.A1(_01927_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_08216_));
 OAI21x1_ASAP7_75t_R _26670_ (.A1(_02121_),
    .A2(_07367_),
    .B(_08216_),
    .Y(_08217_));
 AO21x1_ASAP7_75t_R _26671_ (.A1(net3570),
    .A2(_06947_),
    .B(_08217_),
    .Y(_08218_));
 OA22x2_ASAP7_75t_R _26672_ (.A1(_02154_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02048_),
    .Y(_08219_));
 OA222x2_ASAP7_75t_R _26673_ (.A1(_01977_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02080_),
    .C1(_07028_),
    .C2(_02011_),
    .Y(_08220_));
 OAI21x1_ASAP7_75t_R _26674_ (.A1(_07021_),
    .A2(_08219_),
    .B(_08220_),
    .Y(_08221_));
 OR5x2_ASAP7_75t_R _26675_ (.A(_08212_),
    .B(_08214_),
    .C(_08215_),
    .D(_08218_),
    .E(_08221_),
    .Y(_08222_));
 OR3x1_ASAP7_75t_R _26676_ (.A(_07474_),
    .B(_08210_),
    .C(_08222_),
    .Y(_08223_));
 AO21x1_ASAP7_75t_R _26677_ (.A1(_07077_),
    .A2(_07990_),
    .B(_08223_),
    .Y(_08224_));
 OA22x2_ASAP7_75t_R _26678_ (.A1(_08113_),
    .A2(_08198_),
    .B1(_08206_),
    .B2(_08224_),
    .Y(_08225_));
 NOR2x1_ASAP7_75t_R _26679_ (.A(_01691_),
    .B(_06987_),
    .Y(_08226_));
 AO21x1_ASAP7_75t_R _26680_ (.A1(_06987_),
    .A2(_08225_),
    .B(_08226_),
    .Y(_02674_));
 TAPCELL_ASAP7_75t_R PHY_683 ();
 AND2x2_ASAP7_75t_R _26682_ (.A(net52),
    .B(net434),
    .Y(_08228_));
 AO21x1_ASAP7_75t_R _26683_ (.A1(net29),
    .A2(_07051_),
    .B(_08228_),
    .Y(_08229_));
 NAND2x1_ASAP7_75t_R _26684_ (.A(net37),
    .B(net434),
    .Y(_08230_));
 OA211x2_ASAP7_75t_R _26685_ (.A1(net434),
    .A2(_01852_),
    .B(_08230_),
    .C(_01642_),
    .Y(_08231_));
 INVx1_ASAP7_75t_R _26686_ (.A(_08231_),
    .Y(_08232_));
 OA211x2_ASAP7_75t_R _26687_ (.A1(_01642_),
    .A2(_08229_),
    .B(_08232_),
    .C(_07036_),
    .Y(_08233_));
 AND3x1_ASAP7_75t_R _26688_ (.A(_00125_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08234_));
 AOI211x1_ASAP7_75t_R _26689_ (.A1(_00124_),
    .A2(_07238_),
    .B(_08234_),
    .C(_07234_),
    .Y(_08235_));
 AO21x1_ASAP7_75t_R _26690_ (.A1(_02379_),
    .A2(_07234_),
    .B(_08235_),
    .Y(_08236_));
 AO221x1_ASAP7_75t_R _26691_ (.A1(net160),
    .A2(_07242_),
    .B1(_08236_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08237_));
 OR3x1_ASAP7_75t_R _26692_ (.A(_02231_),
    .B(_05815_),
    .C(_07061_),
    .Y(_08238_));
 XNOR2x1_ASAP7_75t_R _26693_ (.B(_02242_),
    .Y(_08239_),
    .A(net2165));
 NAND2x1_ASAP7_75t_R _26694_ (.A(_07062_),
    .B(_08239_),
    .Y(_08240_));
 AO21x1_ASAP7_75t_R _26695_ (.A1(_08238_),
    .A2(_08240_),
    .B(_05766_),
    .Y(_08241_));
 NAND2x1_ASAP7_75t_R _26696_ (.A(_13570_),
    .B(_00914_),
    .Y(_08242_));
 AO21x1_ASAP7_75t_R _26697_ (.A1(_08241_),
    .A2(_08242_),
    .B(net308),
    .Y(_08243_));
 AO32x1_ASAP7_75t_R _26698_ (.A1(_07215_),
    .A2(_07218_),
    .A3(_07493_),
    .B1(_08237_),
    .B2(_08243_),
    .Y(_08244_));
 OA22x2_ASAP7_75t_R _26699_ (.A1(_01500_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01469_),
    .Y(_08245_));
 OAI22x1_ASAP7_75t_R _26700_ (.A1(_02153_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02047_),
    .Y(_08246_));
 NAND2x1_ASAP7_75t_R _26701_ (.A(_06940_),
    .B(_08246_),
    .Y(_08247_));
 OA22x2_ASAP7_75t_R _26702_ (.A1(_02079_),
    .A2(_07026_),
    .B1(_07008_),
    .B2(_00126_),
    .Y(_08248_));
 NAND2x1_ASAP7_75t_R _26703_ (.A(net3704),
    .B(_08134_),
    .Y(_08249_));
 OA211x2_ASAP7_75t_R _26704_ (.A1(_02010_),
    .A2(_07028_),
    .B(_08248_),
    .C(_08249_),
    .Y(_08250_));
 NAND2x1_ASAP7_75t_R _26705_ (.A(net3710),
    .B(_06947_),
    .Y(_08251_));
 OA21x2_ASAP7_75t_R _26706_ (.A1(_01926_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_08252_));
 OA211x2_ASAP7_75t_R _26707_ (.A1(_02120_),
    .A2(_07367_),
    .B(_08251_),
    .C(_08252_),
    .Y(_08253_));
 OA222x2_ASAP7_75t_R _26708_ (.A1(_01562_),
    .A2(_07369_),
    .B1(_07522_),
    .B2(_01960_),
    .C1(_01976_),
    .C2(_07024_),
    .Y(_08254_));
 AND4x1_ASAP7_75t_R _26709_ (.A(_08247_),
    .B(_08250_),
    .C(_08253_),
    .D(_08254_),
    .Y(_08255_));
 OA21x2_ASAP7_75t_R _26710_ (.A1(_07360_),
    .A2(_08245_),
    .B(_08255_),
    .Y(_08256_));
 INVx1_ASAP7_75t_R _26711_ (.A(_08256_),
    .Y(_08257_));
 AND2x2_ASAP7_75t_R _26712_ (.A(_07125_),
    .B(_07568_),
    .Y(_08258_));
 AO21x1_ASAP7_75t_R _26713_ (.A1(_07152_),
    .A2(_07577_),
    .B(_08258_),
    .Y(_08259_));
 OA21x2_ASAP7_75t_R _26714_ (.A1(_07218_),
    .A2(_07513_),
    .B(_07077_),
    .Y(_08260_));
 OA21x2_ASAP7_75t_R _26715_ (.A1(_07073_),
    .A2(_08259_),
    .B(_08260_),
    .Y(_08261_));
 OR4x2_ASAP7_75t_R _26716_ (.A(_08147_),
    .B(_08244_),
    .C(_08257_),
    .D(_08261_),
    .Y(_08262_));
 OA21x2_ASAP7_75t_R _26717_ (.A1(_08113_),
    .A2(_08233_),
    .B(_08262_),
    .Y(_08263_));
 NOR2x1_ASAP7_75t_R _26718_ (.A(_01690_),
    .B(net288),
    .Y(_08264_));
 AO21x1_ASAP7_75t_R _26719_ (.A1(net288),
    .A2(_08263_),
    .B(_08264_),
    .Y(_02675_));
 AND3x1_ASAP7_75t_R _26720_ (.A(_00128_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08265_));
 AOI211x1_ASAP7_75t_R _26721_ (.A1(_00127_),
    .A2(_07238_),
    .B(_08265_),
    .C(_07234_),
    .Y(_08266_));
 AO21x1_ASAP7_75t_R _26722_ (.A1(_02380_),
    .A2(_07234_),
    .B(_08266_),
    .Y(_08267_));
 AO22x2_ASAP7_75t_R _26723_ (.A1(net161),
    .A2(_07242_),
    .B1(_08267_),
    .B2(_07231_),
    .Y(_08268_));
 NOR2x1_ASAP7_75t_R _26724_ (.A(_01376_),
    .B(_07062_),
    .Y(_08269_));
 AO21x1_ASAP7_75t_R _26725_ (.A1(_02245_),
    .A2(_07062_),
    .B(_08269_),
    .Y(_08270_));
 OA21x2_ASAP7_75t_R _26726_ (.A1(_05766_),
    .A2(_08270_),
    .B(_13817_),
    .Y(_08271_));
 NAND2x1_ASAP7_75t_R _26727_ (.A(_00946_),
    .B(_07059_),
    .Y(_08272_));
 AO22x1_ASAP7_75t_R _26728_ (.A1(net308),
    .A2(_08268_),
    .B1(_08271_),
    .B2(_08272_),
    .Y(_08273_));
 OA211x2_ASAP7_75t_R _26729_ (.A1(_07487_),
    .A2(_07490_),
    .B(_07077_),
    .C(_07310_),
    .Y(_08274_));
 AOI211x1_ASAP7_75t_R _26730_ (.A1(_07571_),
    .A2(_08204_),
    .B(_08273_),
    .C(_08274_),
    .Y(_08275_));
 OA22x2_ASAP7_75t_R _26731_ (.A1(_01499_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01468_),
    .Y(_08276_));
 OA22x2_ASAP7_75t_R _26732_ (.A1(_02152_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02046_),
    .Y(_08277_));
 OA22x2_ASAP7_75t_R _26733_ (.A1(_01975_),
    .A2(_07024_),
    .B1(_07008_),
    .B2(_00129_),
    .Y(_08278_));
 OA22x2_ASAP7_75t_R _26734_ (.A1(_01959_),
    .A2(_07522_),
    .B1(_07745_),
    .B2(_06283_),
    .Y(_08279_));
 OA211x2_ASAP7_75t_R _26735_ (.A1(_07021_),
    .A2(_08277_),
    .B(_08278_),
    .C(_08279_),
    .Y(_08280_));
 OA222x2_ASAP7_75t_R _26736_ (.A1(_01925_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02119_),
    .C1(_07369_),
    .C2(_01561_),
    .Y(_08281_));
 OA33x2_ASAP7_75t_R _26737_ (.A1(_02078_),
    .A2(_05589_),
    .A3(_06994_),
    .B1(_07023_),
    .B2(_06990_),
    .B3(_02009_),
    .Y(_08282_));
 NAND2x1_ASAP7_75t_R _26738_ (.A(net3680),
    .B(_06947_),
    .Y(_08283_));
 AND4x1_ASAP7_75t_R _26739_ (.A(_07791_),
    .B(_08281_),
    .C(_08282_),
    .D(_08283_),
    .Y(_08284_));
 OA211x2_ASAP7_75t_R _26740_ (.A1(_07360_),
    .A2(_08276_),
    .B(_08280_),
    .C(_08284_),
    .Y(_08285_));
 NAND2x1_ASAP7_75t_R _26741_ (.A(_08275_),
    .B(_08285_),
    .Y(_08286_));
 AO21x1_ASAP7_75t_R _26742_ (.A1(_07077_),
    .A2(_07906_),
    .B(_08147_),
    .Y(_08287_));
 NAND2x1_ASAP7_75t_R _26743_ (.A(net53),
    .B(net433),
    .Y(_08288_));
 OA211x2_ASAP7_75t_R _26744_ (.A1(_07952_),
    .A2(net433),
    .B(_08288_),
    .C(_07039_),
    .Y(_08289_));
 NAND2x1_ASAP7_75t_R _26745_ (.A(net39),
    .B(net433),
    .Y(_08290_));
 OA211x2_ASAP7_75t_R _26746_ (.A1(net433),
    .A2(_01851_),
    .B(_08290_),
    .C(net432),
    .Y(_08291_));
 NOR2x1_ASAP7_75t_R _26747_ (.A(_08289_),
    .B(_08291_),
    .Y(_08292_));
 AO21x2_ASAP7_75t_R _26748_ (.A1(_07036_),
    .A2(_08292_),
    .B(_08113_),
    .Y(_08293_));
 OA21x2_ASAP7_75t_R _26749_ (.A1(_08286_),
    .A2(_08287_),
    .B(_08293_),
    .Y(_08294_));
 NOR2x1_ASAP7_75t_R _26750_ (.A(_01689_),
    .B(_06987_),
    .Y(_08295_));
 AO21x1_ASAP7_75t_R _26751_ (.A1(_06987_),
    .A2(_08294_),
    .B(_08295_),
    .Y(_02676_));
 OA211x2_ASAP7_75t_R _26752_ (.A1(_07218_),
    .A2(_07617_),
    .B(_07888_),
    .C(_07077_),
    .Y(_08296_));
 OAI21x1_ASAP7_75t_R _26753_ (.A1(_07073_),
    .A2(_07886_),
    .B(_08204_),
    .Y(_08297_));
 AND3x1_ASAP7_75t_R _26754_ (.A(_00131_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08298_));
 AOI211x1_ASAP7_75t_R _26755_ (.A1(_00130_),
    .A2(_07238_),
    .B(_08298_),
    .C(_07234_),
    .Y(_08299_));
 AO21x1_ASAP7_75t_R _26756_ (.A1(_02381_),
    .A2(_07234_),
    .B(_08299_),
    .Y(_08300_));
 AO22x1_ASAP7_75t_R _26757_ (.A1(net162),
    .A2(_07242_),
    .B1(_08300_),
    .B2(_07231_),
    .Y(_08301_));
 XNOR2x2_ASAP7_75t_R _26758_ (.A(_00044_),
    .B(_02244_),
    .Y(_08302_));
 NAND2x1_ASAP7_75t_R _26759_ (.A(_07062_),
    .B(_08302_),
    .Y(_08303_));
 OA21x2_ASAP7_75t_R _26760_ (.A1(_07062_),
    .A2(_07639_),
    .B(_08303_),
    .Y(_08304_));
 OA21x2_ASAP7_75t_R _26761_ (.A1(_05766_),
    .A2(_08304_),
    .B(_13817_),
    .Y(_08305_));
 NAND2x1_ASAP7_75t_R _26762_ (.A(_00979_),
    .B(_07059_),
    .Y(_08306_));
 AOI22x1_ASAP7_75t_R _26763_ (.A1(net308),
    .A2(_08301_),
    .B1(_08305_),
    .B2(_08306_),
    .Y(_08307_));
 OA22x2_ASAP7_75t_R _26764_ (.A1(_01498_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01467_),
    .Y(_08308_));
 OA22x2_ASAP7_75t_R _26765_ (.A1(_02151_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02045_),
    .Y(_08309_));
 INVx1_ASAP7_75t_R _26766_ (.A(net3533),
    .Y(_08310_));
 OA222x2_ASAP7_75t_R _26767_ (.A1(_02077_),
    .A2(_07026_),
    .B1(_07522_),
    .B2(_01958_),
    .C1(_08310_),
    .C2(_07745_),
    .Y(_08311_));
 OA21x2_ASAP7_75t_R _26768_ (.A1(_07021_),
    .A2(_08309_),
    .B(_08311_),
    .Y(_08312_));
 OA22x2_ASAP7_75t_R _26769_ (.A1(_02008_),
    .A2(_07028_),
    .B1(_07008_),
    .B2(_00132_),
    .Y(_08313_));
 OA22x2_ASAP7_75t_R _26770_ (.A1(_01974_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01560_),
    .Y(_08314_));
 OA22x2_ASAP7_75t_R _26771_ (.A1(_02118_),
    .A2(_07367_),
    .B1(_07740_),
    .B2(_01997_),
    .Y(_08315_));
 OA211x2_ASAP7_75t_R _26772_ (.A1(_01924_),
    .A2(_06998_),
    .B(_07004_),
    .C(_08315_),
    .Y(_08316_));
 NAND2x1_ASAP7_75t_R _26773_ (.A(net3675),
    .B(_06947_),
    .Y(_08317_));
 AND5x1_ASAP7_75t_R _26774_ (.A(_08312_),
    .B(_08313_),
    .C(_08314_),
    .D(_08316_),
    .E(net3676),
    .Y(_08318_));
 OA21x2_ASAP7_75t_R _26775_ (.A1(_07360_),
    .A2(_08308_),
    .B(_08318_),
    .Y(_08319_));
 AND3x2_ASAP7_75t_R _26776_ (.A(_06981_),
    .B(_08307_),
    .C(_08319_),
    .Y(_08320_));
 NAND2x1_ASAP7_75t_R _26777_ (.A(_08297_),
    .B(_08320_),
    .Y(_08321_));
 AND2x2_ASAP7_75t_R _26778_ (.A(net54),
    .B(net433),
    .Y(_08322_));
 AO21x1_ASAP7_75t_R _26779_ (.A1(net31),
    .A2(_07051_),
    .B(_08322_),
    .Y(_08323_));
 NAND2x1_ASAP7_75t_R _26780_ (.A(net40),
    .B(net433),
    .Y(_08324_));
 OA211x2_ASAP7_75t_R _26781_ (.A1(net433),
    .A2(_01850_),
    .B(_08324_),
    .C(net432),
    .Y(_08325_));
 INVx1_ASAP7_75t_R _26782_ (.A(_08325_),
    .Y(_08326_));
 OA211x2_ASAP7_75t_R _26783_ (.A1(net432),
    .A2(_08323_),
    .B(_08326_),
    .C(_07036_),
    .Y(_08327_));
 OA22x2_ASAP7_75t_R _26784_ (.A1(_08296_),
    .A2(_08321_),
    .B1(_08327_),
    .B2(_08113_),
    .Y(_08328_));
 NOR2x1_ASAP7_75t_R _26785_ (.A(_01688_),
    .B(net288),
    .Y(_08329_));
 AO21x1_ASAP7_75t_R _26786_ (.A1(net288),
    .A2(_08328_),
    .B(_08329_),
    .Y(_02677_));
 NAND2x1_ASAP7_75t_R _26787_ (.A(net55),
    .B(net434),
    .Y(_08330_));
 OA211x2_ASAP7_75t_R _26788_ (.A1(_08030_),
    .A2(net434),
    .B(_08330_),
    .C(_07039_),
    .Y(_08331_));
 NAND2x1_ASAP7_75t_R _26789_ (.A(net41),
    .B(net434),
    .Y(_08332_));
 OA211x2_ASAP7_75t_R _26790_ (.A1(net434),
    .A2(_01849_),
    .B(_08332_),
    .C(net432),
    .Y(_08333_));
 NOR2x1_ASAP7_75t_R _26791_ (.A(_08331_),
    .B(_08333_),
    .Y(_08334_));
 AOI21x1_ASAP7_75t_R _26792_ (.A1(_07036_),
    .A2(_08334_),
    .B(_08113_),
    .Y(_08335_));
 NAND2x1_ASAP7_75t_R _26793_ (.A(_07215_),
    .B(_07835_),
    .Y(_08336_));
 AND2x2_ASAP7_75t_R _26794_ (.A(_07073_),
    .B(_07077_),
    .Y(_08337_));
 OA211x2_ASAP7_75t_R _26795_ (.A1(_07125_),
    .A2(_07829_),
    .B(_07426_),
    .C(_07830_),
    .Y(_08338_));
 AOI21x1_ASAP7_75t_R _26796_ (.A1(_07828_),
    .A2(_08337_),
    .B(_08338_),
    .Y(_08339_));
 AND3x1_ASAP7_75t_R _26797_ (.A(_00134_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08340_));
 AOI211x1_ASAP7_75t_R _26798_ (.A1(_00133_),
    .A2(_07238_),
    .B(_08340_),
    .C(_07234_),
    .Y(_08341_));
 AO21x1_ASAP7_75t_R _26799_ (.A1(_02382_),
    .A2(_07234_),
    .B(_08341_),
    .Y(_08342_));
 AOI22x1_ASAP7_75t_R _26800_ (.A1(net163),
    .A2(_07242_),
    .B1(_08342_),
    .B2(_07231_),
    .Y(_08343_));
 NOR2x1_ASAP7_75t_R _26801_ (.A(_02247_),
    .B(_07064_),
    .Y(_08344_));
 AO21x1_ASAP7_75t_R _26802_ (.A1(_07684_),
    .A2(_07064_),
    .B(_08344_),
    .Y(_08345_));
 AO221x1_ASAP7_75t_R _26803_ (.A1(_01011_),
    .A2(_07059_),
    .B1(_07060_),
    .B2(_08345_),
    .C(net308),
    .Y(_08346_));
 OA211x2_ASAP7_75t_R _26804_ (.A1(_13817_),
    .A2(_08343_),
    .B(_08346_),
    .C(_06981_),
    .Y(_08347_));
 OA22x2_ASAP7_75t_R _26805_ (.A1(_01497_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01466_),
    .Y(_08348_));
 OA22x2_ASAP7_75t_R _26806_ (.A1(_02150_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02044_),
    .Y(_08349_));
 INVx1_ASAP7_75t_R _26807_ (.A(net3566),
    .Y(_08350_));
 OA222x2_ASAP7_75t_R _26808_ (.A1(_02076_),
    .A2(_07026_),
    .B1(_07008_),
    .B2(_00135_),
    .C1(_08350_),
    .C2(_07745_),
    .Y(_08351_));
 OA21x2_ASAP7_75t_R _26809_ (.A1(_07021_),
    .A2(_08349_),
    .B(_08351_),
    .Y(_08352_));
 OA22x2_ASAP7_75t_R _26810_ (.A1(_02007_),
    .A2(_07028_),
    .B1(_07522_),
    .B2(_01957_),
    .Y(_08353_));
 OA22x2_ASAP7_75t_R _26811_ (.A1(_01973_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01559_),
    .Y(_08354_));
 OA22x2_ASAP7_75t_R _26812_ (.A1(_01923_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02117_),
    .Y(_08355_));
 NAND2x1_ASAP7_75t_R _26813_ (.A(net3688),
    .B(_07700_),
    .Y(_08356_));
 AND5x2_ASAP7_75t_R _26814_ (.A(_07004_),
    .B(_08353_),
    .C(_08354_),
    .D(_08355_),
    .E(net3689),
    .Y(_08357_));
 OA211x2_ASAP7_75t_R _26815_ (.A1(_07360_),
    .A2(_08348_),
    .B(_08352_),
    .C(_08357_),
    .Y(_08358_));
 AND4x2_ASAP7_75t_R _26816_ (.A(_08336_),
    .B(_08339_),
    .C(_08347_),
    .D(_08358_),
    .Y(_08359_));
 NOR2x2_ASAP7_75t_R _26817_ (.A(_08335_),
    .B(_08359_),
    .Y(_08360_));
 NOR2x1_ASAP7_75t_R _26818_ (.A(_01687_),
    .B(_06987_),
    .Y(_08361_));
 AO21x1_ASAP7_75t_R _26819_ (.A1(_06987_),
    .A2(_08360_),
    .B(_08361_),
    .Y(_02678_));
 AND2x2_ASAP7_75t_R _26820_ (.A(_07077_),
    .B(_07774_),
    .Y(_08362_));
 OA21x2_ASAP7_75t_R _26821_ (.A1(_07073_),
    .A2(_07714_),
    .B(_08204_),
    .Y(_08363_));
 AND3x1_ASAP7_75t_R _26822_ (.A(_00137_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08364_));
 AOI211x1_ASAP7_75t_R _26823_ (.A1(_00136_),
    .A2(_07238_),
    .B(_08364_),
    .C(_07234_),
    .Y(_08365_));
 AO21x1_ASAP7_75t_R _26824_ (.A1(_02383_),
    .A2(_07234_),
    .B(_08365_),
    .Y(_08366_));
 AO22x1_ASAP7_75t_R _26825_ (.A1(net164),
    .A2(_07242_),
    .B1(_08366_),
    .B2(_07231_),
    .Y(_08367_));
 XNOR2x1_ASAP7_75t_R _26826_ (.B(_02246_),
    .Y(_08368_),
    .A(net2135));
 AND2x2_ASAP7_75t_R _26827_ (.A(_07062_),
    .B(_08368_),
    .Y(_08369_));
 AO21x1_ASAP7_75t_R _26828_ (.A1(_07064_),
    .A2(_07727_),
    .B(_08369_),
    .Y(_08370_));
 NAND2x2_ASAP7_75t_R _26829_ (.A(_07060_),
    .B(_08370_),
    .Y(_08371_));
 NAND2x1_ASAP7_75t_R _26830_ (.A(_01045_),
    .B(_07059_),
    .Y(_08372_));
 AND3x1_ASAP7_75t_R _26831_ (.A(_13817_),
    .B(_08371_),
    .C(_08372_),
    .Y(_08373_));
 AO21x1_ASAP7_75t_R _26832_ (.A1(net308),
    .A2(_08367_),
    .B(_08373_),
    .Y(_08374_));
 NAND2x1_ASAP7_75t_R _26833_ (.A(_14180_),
    .B(_14239_),
    .Y(_08375_));
 AO21x1_ASAP7_75t_R _26834_ (.A1(_14239_),
    .A2(_05662_),
    .B(_14180_),
    .Y(_08376_));
 AND2x2_ASAP7_75t_R _26835_ (.A(_13894_),
    .B(_14239_),
    .Y(_08377_));
 AO221x1_ASAP7_75t_R _26836_ (.A1(_05707_),
    .A2(_08375_),
    .B1(_08376_),
    .B2(_13525_),
    .C(_08377_),
    .Y(_08378_));
 AND3x1_ASAP7_75t_R _26837_ (.A(_14179_),
    .B(_14238_),
    .C(_05662_),
    .Y(_08379_));
 AO21x1_ASAP7_75t_R _26838_ (.A1(_14297_),
    .A2(_05610_),
    .B(_08379_),
    .Y(_08380_));
 AO221x1_ASAP7_75t_R _26839_ (.A1(_14239_),
    .A2(_05610_),
    .B1(_08378_),
    .B2(net302),
    .C(_08380_),
    .Y(_08381_));
 INVx1_ASAP7_75t_R _26840_ (.A(_05711_),
    .Y(_08382_));
 AND2x2_ASAP7_75t_R _26841_ (.A(_14297_),
    .B(_14359_),
    .Y(_08383_));
 OA211x2_ASAP7_75t_R _26842_ (.A1(_08382_),
    .A2(_05707_),
    .B(_05652_),
    .C(_08383_),
    .Y(_08384_));
 AOI211x1_ASAP7_75t_R _26843_ (.A1(_14359_),
    .A2(_08381_),
    .B(_08384_),
    .C(_05563_),
    .Y(_08385_));
 AO22x1_ASAP7_75t_R _26844_ (.A1(_05594_),
    .A2(_14424_),
    .B1(_05595_),
    .B2(_13474_),
    .Y(_08386_));
 OA22x2_ASAP7_75t_R _26845_ (.A1(_01496_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01465_),
    .Y(_08387_));
 AO21x1_ASAP7_75t_R _26846_ (.A1(net310),
    .A2(_08386_),
    .B(_08387_),
    .Y(_08388_));
 OR3x1_ASAP7_75t_R _26847_ (.A(_05623_),
    .B(_08385_),
    .C(_08388_),
    .Y(_08389_));
 OAI22x1_ASAP7_75t_R _26848_ (.A1(_00138_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01558_),
    .Y(_08390_));
 AO32x1_ASAP7_75t_R _26849_ (.A1(_06239_),
    .A2(_06942_),
    .A3(_08213_),
    .B1(_08134_),
    .B2(net3492),
    .Y(_08391_));
 NOR2x1_ASAP7_75t_R _26850_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 NAND2x1_ASAP7_75t_R _26851_ (.A(net3579),
    .B(_06947_),
    .Y(_08393_));
 OR3x1_ASAP7_75t_R _26852_ (.A(_01922_),
    .B(_06938_),
    .C(_06990_),
    .Y(_08394_));
 OA211x2_ASAP7_75t_R _26853_ (.A1(_02116_),
    .A2(_07367_),
    .B(_08394_),
    .C(_07004_),
    .Y(_08395_));
 OA22x2_ASAP7_75t_R _26854_ (.A1(_02149_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02043_),
    .Y(_08396_));
 OA222x2_ASAP7_75t_R _26855_ (.A1(_01972_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02075_),
    .C1(_07028_),
    .C2(_02006_),
    .Y(_08397_));
 OA21x2_ASAP7_75t_R _26856_ (.A1(_07021_),
    .A2(_08396_),
    .B(_08397_),
    .Y(_08398_));
 AND5x2_ASAP7_75t_R _26857_ (.A(_08389_),
    .B(_08392_),
    .C(_08393_),
    .D(_08395_),
    .E(_08398_),
    .Y(_08399_));
 INVx1_ASAP7_75t_R _26858_ (.A(_08399_),
    .Y(_08400_));
 OR4x1_ASAP7_75t_R _26859_ (.A(_07474_),
    .B(_08363_),
    .C(_08374_),
    .D(_08400_),
    .Y(_08401_));
 INVx1_ASAP7_75t_R _26860_ (.A(_01733_),
    .Y(_08402_));
 OA211x2_ASAP7_75t_R _26861_ (.A1(net434),
    .A2(_08402_),
    .B(_07819_),
    .C(net432),
    .Y(_08403_));
 AO21x1_ASAP7_75t_R _26862_ (.A1(_07039_),
    .A2(_07818_),
    .B(_08403_),
    .Y(_08404_));
 AO21x2_ASAP7_75t_R _26863_ (.A1(_07036_),
    .A2(_08404_),
    .B(_08113_),
    .Y(_08405_));
 OA21x2_ASAP7_75t_R _26864_ (.A1(_08362_),
    .A2(_08401_),
    .B(_08405_),
    .Y(_08406_));
 NOR2x1_ASAP7_75t_R _26865_ (.A(_01686_),
    .B(_06987_),
    .Y(_08407_));
 AO21x1_ASAP7_75t_R _26866_ (.A1(_06987_),
    .A2(_08406_),
    .B(_08407_),
    .Y(_02679_));
 AND3x1_ASAP7_75t_R _26867_ (.A(_00140_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08408_));
 AOI211x1_ASAP7_75t_R _26868_ (.A1(_00139_),
    .A2(_07238_),
    .B(_08408_),
    .C(_07234_),
    .Y(_08409_));
 AO21x1_ASAP7_75t_R _26869_ (.A1(_02384_),
    .A2(_07234_),
    .B(_08409_),
    .Y(_08410_));
 AO221x2_ASAP7_75t_R _26870_ (.A1(net165),
    .A2(_07242_),
    .B1(_08410_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08411_));
 OA211x2_ASAP7_75t_R _26871_ (.A1(_07733_),
    .A2(_07125_),
    .B(_07227_),
    .C(_07215_),
    .Y(_08412_));
 TAPCELL_ASAP7_75t_R PHY_682 ();
 AND2x2_ASAP7_75t_R _26873_ (.A(_02249_),
    .B(_07062_),
    .Y(_08414_));
 AO221x1_ASAP7_75t_R _26874_ (.A1(_13537_),
    .A2(_07059_),
    .B1(_07064_),
    .B2(_02235_),
    .C(_08414_),
    .Y(_08415_));
 INVx1_ASAP7_75t_R _26875_ (.A(_08415_),
    .Y(_08416_));
 AOI21x1_ASAP7_75t_R _26876_ (.A1(_01077_),
    .A2(_07059_),
    .B(_08416_),
    .Y(_08417_));
 OA33x2_ASAP7_75t_R _26877_ (.A1(_07834_),
    .A2(_08411_),
    .A3(_08412_),
    .B1(_08417_),
    .B2(_05545_),
    .B3(_13612_),
    .Y(_08418_));
 OR2x2_ASAP7_75t_R _26878_ (.A(_07125_),
    .B(_07718_),
    .Y(_08419_));
 OA211x2_ASAP7_75t_R _26879_ (.A1(_07152_),
    .A2(_07716_),
    .B(_08419_),
    .C(_07426_),
    .Y(_08420_));
 AO21x1_ASAP7_75t_R _26880_ (.A1(_07714_),
    .A2(_08337_),
    .B(_07474_),
    .Y(_08421_));
 OAI22x1_ASAP7_75t_R _26881_ (.A1(_01495_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01464_),
    .Y(_08422_));
 OR3x1_ASAP7_75t_R _26882_ (.A(_13525_),
    .B(net305),
    .C(_05563_),
    .Y(_08423_));
 AO21x1_ASAP7_75t_R _26883_ (.A1(_14239_),
    .A2(_05645_),
    .B(_14179_),
    .Y(_08424_));
 AND3x1_ASAP7_75t_R _26884_ (.A(_13525_),
    .B(_13894_),
    .C(_06954_),
    .Y(_08425_));
 AND2x2_ASAP7_75t_R _26885_ (.A(_05568_),
    .B(_05616_),
    .Y(_08426_));
 OA211x2_ASAP7_75t_R _26886_ (.A1(_05693_),
    .A2(_08425_),
    .B(_08426_),
    .C(_08383_),
    .Y(_08427_));
 OA21x2_ASAP7_75t_R _26887_ (.A1(_08424_),
    .A2(_08427_),
    .B(net310),
    .Y(_08428_));
 AO21x1_ASAP7_75t_R _26888_ (.A1(_06968_),
    .A2(_08423_),
    .B(_08428_),
    .Y(_08429_));
 OR3x1_ASAP7_75t_R _26889_ (.A(_07440_),
    .B(_07530_),
    .C(_08428_),
    .Y(_08430_));
 AND3x1_ASAP7_75t_R _26890_ (.A(_14297_),
    .B(_14359_),
    .C(net310),
    .Y(_08431_));
 OA211x2_ASAP7_75t_R _26891_ (.A1(_05707_),
    .A2(_05667_),
    .B(_05682_),
    .C(_14359_),
    .Y(_08432_));
 AO221x1_ASAP7_75t_R _26892_ (.A1(_05627_),
    .A2(_08429_),
    .B1(_08430_),
    .B2(_08431_),
    .C(_08432_),
    .Y(_08433_));
 OAI22x1_ASAP7_75t_R _26893_ (.A1(_02148_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02042_),
    .Y(_08434_));
 AND2x2_ASAP7_75t_R _26894_ (.A(_08426_),
    .B(_08434_),
    .Y(_08435_));
 OAI22x1_ASAP7_75t_R _26895_ (.A1(_01921_),
    .A2(_06938_),
    .B1(_07023_),
    .B2(_02005_),
    .Y(_08436_));
 INVx1_ASAP7_75t_R _26896_ (.A(_02115_),
    .Y(_08437_));
 AO32x1_ASAP7_75t_R _26897_ (.A1(net3521),
    .A2(_05647_),
    .A3(_05707_),
    .B1(_05693_),
    .B2(_08437_),
    .Y(_08438_));
 OA21x2_ASAP7_75t_R _26898_ (.A1(_08436_),
    .A2(_08438_),
    .B(_06965_),
    .Y(_08439_));
 OAI22x1_ASAP7_75t_R _26899_ (.A1(_00141_),
    .A2(_07008_),
    .B1(_07522_),
    .B2(_01955_),
    .Y(_08440_));
 OAI22x1_ASAP7_75t_R _26900_ (.A1(_01971_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02074_),
    .Y(_08441_));
 OAI21x1_ASAP7_75t_R _26901_ (.A1(_01557_),
    .A2(_07369_),
    .B(_07004_),
    .Y(_08442_));
 AO21x1_ASAP7_75t_R _26902_ (.A1(net3590),
    .A2(_06947_),
    .B(_08442_),
    .Y(_08443_));
 OR4x1_ASAP7_75t_R _26903_ (.A(_08439_),
    .B(_08440_),
    .C(_08441_),
    .D(_08443_),
    .Y(_08444_));
 AO221x2_ASAP7_75t_R _26904_ (.A1(_06950_),
    .A2(_08422_),
    .B1(_08433_),
    .B2(_08435_),
    .C(_08444_),
    .Y(_08445_));
 OR3x1_ASAP7_75t_R _26905_ (.A(_08420_),
    .B(_08421_),
    .C(_08445_),
    .Y(_08446_));
 OA211x2_ASAP7_75t_R _26906_ (.A1(net34),
    .A2(net433),
    .B(_07807_),
    .C(_07039_),
    .Y(_08447_));
 AO21x1_ASAP7_75t_R _26907_ (.A1(net432),
    .A2(_07804_),
    .B(_08447_),
    .Y(_08448_));
 AO21x2_ASAP7_75t_R _26908_ (.A1(_07036_),
    .A2(_08448_),
    .B(_08113_),
    .Y(_08449_));
 OA21x2_ASAP7_75t_R _26909_ (.A1(_08418_),
    .A2(_08446_),
    .B(_08449_),
    .Y(_08450_));
 NOR2x1_ASAP7_75t_R _26910_ (.A(_01685_),
    .B(_06987_),
    .Y(_08451_));
 AO21x1_ASAP7_75t_R _26911_ (.A1(_06987_),
    .A2(_08450_),
    .B(_08451_),
    .Y(_02680_));
 NAND2x1_ASAP7_75t_R _26912_ (.A(net432),
    .B(_07856_),
    .Y(_08452_));
 OA211x2_ASAP7_75t_R _26913_ (.A1(net432),
    .A2(_07858_),
    .B(_08452_),
    .C(_07036_),
    .Y(_08453_));
 OA211x2_ASAP7_75t_R _26914_ (.A1(_07218_),
    .A2(_07676_),
    .B(_07682_),
    .C(_07077_),
    .Y(_08454_));
 AO21x1_ASAP7_75t_R _26915_ (.A1(_07273_),
    .A2(_07340_),
    .B(_07276_),
    .Y(_08455_));
 AND2x2_ASAP7_75t_R _26916_ (.A(_07215_),
    .B(_08455_),
    .Y(_08456_));
 AND3x1_ASAP7_75t_R _26917_ (.A(_00143_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08457_));
 AOI211x1_ASAP7_75t_R _26918_ (.A1(_00142_),
    .A2(_07238_),
    .B(_08457_),
    .C(_07234_),
    .Y(_08458_));
 AO21x1_ASAP7_75t_R _26919_ (.A1(_02385_),
    .A2(_07234_),
    .B(_08458_),
    .Y(_08459_));
 AO22x2_ASAP7_75t_R _26920_ (.A1(net166),
    .A2(_07242_),
    .B1(_08459_),
    .B2(_07231_),
    .Y(_08460_));
 XNOR2x2_ASAP7_75t_R _26921_ (.A(_00055_),
    .B(_02248_),
    .Y(_08461_));
 NAND2x1_ASAP7_75t_R _26922_ (.A(_07062_),
    .B(_08461_),
    .Y(_08462_));
 OA21x2_ASAP7_75t_R _26923_ (.A1(_07062_),
    .A2(_07837_),
    .B(_08462_),
    .Y(_08463_));
 OA21x2_ASAP7_75t_R _26924_ (.A1(_05766_),
    .A2(_08463_),
    .B(_13817_),
    .Y(_08464_));
 NAND2x1_ASAP7_75t_R _26925_ (.A(_01110_),
    .B(_07059_),
    .Y(_08465_));
 AO22x1_ASAP7_75t_R _26926_ (.A1(net308),
    .A2(_08460_),
    .B1(_08464_),
    .B2(_08465_),
    .Y(_08466_));
 OAI22x1_ASAP7_75t_R _26927_ (.A1(_01494_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01463_),
    .Y(_08467_));
 INVx2_ASAP7_75t_R _26928_ (.A(_00144_),
    .Y(_08468_));
 AO32x1_ASAP7_75t_R _26929_ (.A1(_08468_),
    .A2(_05612_),
    .A3(_05647_),
    .B1(_06942_),
    .B2(_06255_),
    .Y(_08469_));
 OAI22x1_ASAP7_75t_R _26930_ (.A1(_07457_),
    .A2(_06992_),
    .B1(_07024_),
    .B2(_01970_),
    .Y(_08470_));
 AO221x1_ASAP7_75t_R _26931_ (.A1(net3637),
    .A2(_07443_),
    .B1(_07450_),
    .B2(_08469_),
    .C(_08470_),
    .Y(_08471_));
 OAI22x1_ASAP7_75t_R _26932_ (.A1(_02114_),
    .A2(_06992_),
    .B1(_06938_),
    .B2(_01920_),
    .Y(_08472_));
 AO21x1_ASAP7_75t_R _26933_ (.A1(net3477),
    .A2(_06942_),
    .B(_08472_),
    .Y(_08473_));
 OAI22x1_ASAP7_75t_R _26934_ (.A1(_02147_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02041_),
    .Y(_08474_));
 OA222x2_ASAP7_75t_R _26935_ (.A1(_01556_),
    .A2(_07369_),
    .B1(_08102_),
    .B2(_02004_),
    .C1(_02073_),
    .C2(_07026_),
    .Y(_08475_));
 INVx1_ASAP7_75t_R _26936_ (.A(_08475_),
    .Y(_08476_));
 AO221x1_ASAP7_75t_R _26937_ (.A1(_05632_),
    .A2(_08473_),
    .B1(_08474_),
    .B2(_07441_),
    .C(_08476_),
    .Y(_08477_));
 AOI211x1_ASAP7_75t_R _26938_ (.A1(_07438_),
    .A2(_08467_),
    .B(net3638),
    .C(_08477_),
    .Y(_08478_));
 INVx1_ASAP7_75t_R _26939_ (.A(_08478_),
    .Y(_08479_));
 OR5x2_ASAP7_75t_R _26940_ (.A(_07474_),
    .B(_08454_),
    .C(_08456_),
    .D(_08466_),
    .E(_08479_),
    .Y(_08480_));
 OA21x2_ASAP7_75t_R _26941_ (.A1(_08113_),
    .A2(_08453_),
    .B(_08480_),
    .Y(_08481_));
 NOR2x1_ASAP7_75t_R _26942_ (.A(_01684_),
    .B(net288),
    .Y(_08482_));
 AO21x1_ASAP7_75t_R _26943_ (.A1(net288),
    .A2(_08481_),
    .B(_08482_),
    .Y(_02681_));
 OA21x2_ASAP7_75t_R _26944_ (.A1(_07073_),
    .A2(_07617_),
    .B(_08204_),
    .Y(_08483_));
 AND3x1_ASAP7_75t_R _26945_ (.A(_00146_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08484_));
 AOI211x1_ASAP7_75t_R _26946_ (.A1(_00145_),
    .A2(_07238_),
    .B(_08484_),
    .C(_07234_),
    .Y(_08485_));
 AO21x1_ASAP7_75t_R _26947_ (.A1(_02386_),
    .A2(_07234_),
    .B(_08485_),
    .Y(_08486_));
 AOI22x1_ASAP7_75t_R _26948_ (.A1(net167),
    .A2(_07242_),
    .B1(_08486_),
    .B2(_07231_),
    .Y(_08487_));
 NOR2x1_ASAP7_75t_R _26949_ (.A(_02251_),
    .B(_07064_),
    .Y(_08488_));
 AO21x1_ASAP7_75t_R _26950_ (.A1(_07868_),
    .A2(_07064_),
    .B(_08488_),
    .Y(_08489_));
 AO21x1_ASAP7_75t_R _26951_ (.A1(_07060_),
    .A2(_08489_),
    .B(net308),
    .Y(_08490_));
 AO21x1_ASAP7_75t_R _26952_ (.A1(_01142_),
    .A2(_07059_),
    .B(_08490_),
    .Y(_08491_));
 OA211x2_ASAP7_75t_R _26953_ (.A1(_13817_),
    .A2(_08487_),
    .B(_08491_),
    .C(net290),
    .Y(_08492_));
 OA22x2_ASAP7_75t_R _26954_ (.A1(_01493_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01462_),
    .Y(_08493_));
 OA22x2_ASAP7_75t_R _26955_ (.A1(_01969_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01555_),
    .Y(_08494_));
 OA22x2_ASAP7_75t_R _26956_ (.A1(_00147_),
    .A2(_07008_),
    .B1(_07745_),
    .B2(net3408),
    .Y(_08495_));
 OR2x2_ASAP7_75t_R _26957_ (.A(_01919_),
    .B(_06998_),
    .Y(_08496_));
 NAND2x1_ASAP7_75t_R _26958_ (.A(net3750),
    .B(_06947_),
    .Y(_08497_));
 OA21x2_ASAP7_75t_R _26959_ (.A1(_02113_),
    .A2(_07367_),
    .B(_07004_),
    .Y(_08498_));
 AND5x2_ASAP7_75t_R _26960_ (.A(_08494_),
    .B(_08495_),
    .C(_08496_),
    .D(net3751),
    .E(_08498_),
    .Y(_08499_));
 OA22x2_ASAP7_75t_R _26961_ (.A1(_02146_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02040_),
    .Y(_08500_));
 OA222x2_ASAP7_75t_R _26962_ (.A1(_02072_),
    .A2(_07026_),
    .B1(_07028_),
    .B2(_02003_),
    .C1(_01953_),
    .C2(_07522_),
    .Y(_08501_));
 OA21x2_ASAP7_75t_R _26963_ (.A1(_07021_),
    .A2(_08500_),
    .B(_08501_),
    .Y(_08502_));
 OA211x2_ASAP7_75t_R _26964_ (.A1(_07360_),
    .A2(_08493_),
    .B(_08499_),
    .C(_08502_),
    .Y(_08503_));
 NAND2x1_ASAP7_75t_R _26965_ (.A(_08492_),
    .B(_08503_),
    .Y(_08504_));
 AO21x1_ASAP7_75t_R _26966_ (.A1(_07077_),
    .A2(_07631_),
    .B(_08504_),
    .Y(_08505_));
 NOR2x1_ASAP7_75t_R _26967_ (.A(_07039_),
    .B(_07897_),
    .Y(_08506_));
 OA211x2_ASAP7_75t_R _26968_ (.A1(net36),
    .A2(net433),
    .B(_07893_),
    .C(_07039_),
    .Y(_08507_));
 OA21x2_ASAP7_75t_R _26969_ (.A1(_08506_),
    .A2(_08507_),
    .B(_07036_),
    .Y(_08508_));
 OA22x2_ASAP7_75t_R _26970_ (.A1(_08483_),
    .A2(_08505_),
    .B1(_08508_),
    .B2(_08113_),
    .Y(_08509_));
 NOR2x1_ASAP7_75t_R _26971_ (.A(_01683_),
    .B(net288),
    .Y(_08510_));
 AO21x1_ASAP7_75t_R _26972_ (.A1(net288),
    .A2(_08509_),
    .B(_08510_),
    .Y(_02682_));
 OA211x2_ASAP7_75t_R _26973_ (.A1(net37),
    .A2(net434),
    .B(_07940_),
    .C(_07039_),
    .Y(_08511_));
 AO21x1_ASAP7_75t_R _26974_ (.A1(_01642_),
    .A2(_07939_),
    .B(_08511_),
    .Y(_08512_));
 AOI21x1_ASAP7_75t_R _26975_ (.A1(_07036_),
    .A2(_08512_),
    .B(_08113_),
    .Y(_08513_));
 XNOR2x2_ASAP7_75t_R _26976_ (.A(_00058_),
    .B(_02250_),
    .Y(_08514_));
 NOR2x1_ASAP7_75t_R _26977_ (.A(_07062_),
    .B(_07907_),
    .Y(_08515_));
 AO21x1_ASAP7_75t_R _26978_ (.A1(_07062_),
    .A2(_08514_),
    .B(_08515_),
    .Y(_08516_));
 AO221x1_ASAP7_75t_R _26979_ (.A1(_01176_),
    .A2(_07059_),
    .B1(_07060_),
    .B2(_08516_),
    .C(net308),
    .Y(_08517_));
 AND3x1_ASAP7_75t_R _26980_ (.A(_00149_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08518_));
 AOI211x1_ASAP7_75t_R _26981_ (.A1(_00148_),
    .A2(_07238_),
    .B(_08518_),
    .C(_07234_),
    .Y(_08519_));
 AO21x1_ASAP7_75t_R _26982_ (.A1(_02387_),
    .A2(_07234_),
    .B(_08519_),
    .Y(_08520_));
 AO222x2_ASAP7_75t_R _26983_ (.A1(net2157),
    .A2(_07242_),
    .B1(_07561_),
    .B2(_07215_),
    .C1(_08520_),
    .C2(_07231_),
    .Y(_08521_));
 NAND2x1_ASAP7_75t_R _26984_ (.A(net308),
    .B(_08521_),
    .Y(_08522_));
 NAND2x1_ASAP7_75t_R _26985_ (.A(_07077_),
    .B(_07582_),
    .Y(_08523_));
 OA22x2_ASAP7_75t_R _26986_ (.A1(_01492_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01461_),
    .Y(_08524_));
 OA22x2_ASAP7_75t_R _26987_ (.A1(_02145_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02039_),
    .Y(_08525_));
 OA222x2_ASAP7_75t_R _26988_ (.A1(_00150_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01554_),
    .C1(_02002_),
    .C2(_07028_),
    .Y(_08526_));
 OA21x2_ASAP7_75t_R _26989_ (.A1(_07021_),
    .A2(_08525_),
    .B(_08526_),
    .Y(_08527_));
 AO32x1_ASAP7_75t_R _26990_ (.A1(_06280_),
    .A2(_06942_),
    .A3(_08213_),
    .B1(_08134_),
    .B2(net3505),
    .Y(_08528_));
 OAI22x1_ASAP7_75t_R _26991_ (.A1(_01968_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02071_),
    .Y(_08529_));
 NOR2x1_ASAP7_75t_R _26992_ (.A(_08528_),
    .B(_08529_),
    .Y(_08530_));
 NAND2x1_ASAP7_75t_R _26993_ (.A(net3592),
    .B(_06947_),
    .Y(_08531_));
 OA21x2_ASAP7_75t_R _26994_ (.A1(_01918_),
    .A2(_06998_),
    .B(_07004_),
    .Y(_08532_));
 OA21x2_ASAP7_75t_R _26995_ (.A1(_02112_),
    .A2(_07367_),
    .B(_08532_),
    .Y(_08533_));
 AND4x1_ASAP7_75t_R _26996_ (.A(_08527_),
    .B(_08530_),
    .C(net3593),
    .D(_08533_),
    .Y(_08534_));
 OA21x2_ASAP7_75t_R _26997_ (.A1(_07360_),
    .A2(_08524_),
    .B(_08534_),
    .Y(_08535_));
 AND5x2_ASAP7_75t_R _26998_ (.A(net290),
    .B(_08517_),
    .C(_08522_),
    .D(_08523_),
    .E(_08535_),
    .Y(_08536_));
 NOR2x2_ASAP7_75t_R _26999_ (.A(_08513_),
    .B(_08536_),
    .Y(_08537_));
 NOR2x1_ASAP7_75t_R _27000_ (.A(_01682_),
    .B(net288),
    .Y(_08538_));
 AO21x1_ASAP7_75t_R _27001_ (.A1(net288),
    .A2(_08537_),
    .B(_08538_),
    .Y(_02683_));
 NAND2x1_ASAP7_75t_R _27002_ (.A(_02253_),
    .B(_07062_),
    .Y(_08539_));
 OA211x2_ASAP7_75t_R _27003_ (.A1(_07963_),
    .A2(_07062_),
    .B(_08539_),
    .C(_07060_),
    .Y(_08540_));
 AO21x1_ASAP7_75t_R _27004_ (.A1(_01208_),
    .A2(_07059_),
    .B(_08540_),
    .Y(_08541_));
 NAND2x1_ASAP7_75t_R _27005_ (.A(_13817_),
    .B(_08541_),
    .Y(_08542_));
 AND3x1_ASAP7_75t_R _27006_ (.A(_00152_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08543_));
 AOI211x1_ASAP7_75t_R _27007_ (.A1(_00151_),
    .A2(_07238_),
    .B(_08543_),
    .C(_07234_),
    .Y(_08544_));
 AO21x1_ASAP7_75t_R _27008_ (.A1(_02388_),
    .A2(_07234_),
    .B(_08544_),
    .Y(_08545_));
 AO221x1_ASAP7_75t_R _27009_ (.A1(net169),
    .A2(_07242_),
    .B1(_08545_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08546_));
 OA21x2_ASAP7_75t_R _27010_ (.A1(_07073_),
    .A2(_07513_),
    .B(_08204_),
    .Y(_08547_));
 AO221x1_ASAP7_75t_R _27011_ (.A1(_07077_),
    .A2(_07508_),
    .B1(_08542_),
    .B2(_08546_),
    .C(_08547_),
    .Y(_08548_));
 OAI22x1_ASAP7_75t_R _27012_ (.A1(_01491_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01460_),
    .Y(_08549_));
 OA22x2_ASAP7_75t_R _27013_ (.A1(_02144_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02038_),
    .Y(_08550_));
 OA222x2_ASAP7_75t_R _27014_ (.A1(_01967_),
    .A2(_07024_),
    .B1(_07026_),
    .B2(_02070_),
    .C1(_07028_),
    .C2(_02001_),
    .Y(_08551_));
 OAI21x1_ASAP7_75t_R _27015_ (.A1(_07021_),
    .A2(_08550_),
    .B(_08551_),
    .Y(_08552_));
 AO32x1_ASAP7_75t_R _27016_ (.A1(_06261_),
    .A2(_06942_),
    .A3(_08213_),
    .B1(_08134_),
    .B2(net3372),
    .Y(_08553_));
 OAI22x1_ASAP7_75t_R _27017_ (.A1(_00153_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01553_),
    .Y(_08554_));
 OAI22x1_ASAP7_75t_R _27018_ (.A1(_01917_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02111_),
    .Y(_08555_));
 AND2x2_ASAP7_75t_R _27019_ (.A(net3740),
    .B(_07700_),
    .Y(_08556_));
 OR5x2_ASAP7_75t_R _27020_ (.A(_08057_),
    .B(_08553_),
    .C(_08554_),
    .D(_08555_),
    .E(net3741),
    .Y(_08557_));
 AOI211x1_ASAP7_75t_R _27021_ (.A1(_06950_),
    .A2(_08549_),
    .B(_08552_),
    .C(_08557_),
    .Y(_08558_));
 NAND2x1_ASAP7_75t_R _27022_ (.A(net290),
    .B(_08558_),
    .Y(_08559_));
 OA211x2_ASAP7_75t_R _27023_ (.A1(net39),
    .A2(net433),
    .B(_07953_),
    .C(_07039_),
    .Y(_08560_));
 AO21x1_ASAP7_75t_R _27024_ (.A1(net432),
    .A2(_07957_),
    .B(_08560_),
    .Y(_08561_));
 AO21x2_ASAP7_75t_R _27025_ (.A1(_07036_),
    .A2(_08561_),
    .B(_08113_),
    .Y(_08562_));
 OA21x2_ASAP7_75t_R _27026_ (.A1(_08548_),
    .A2(_08559_),
    .B(_08562_),
    .Y(_08563_));
 NOR2x1_ASAP7_75t_R _27027_ (.A(_01681_),
    .B(_06987_),
    .Y(_08564_));
 AO21x1_ASAP7_75t_R _27028_ (.A1(_06987_),
    .A2(_08563_),
    .B(_08564_),
    .Y(_02684_));
 OR3x1_ASAP7_75t_R _27029_ (.A(_07080_),
    .B(_07406_),
    .C(_07418_),
    .Y(_08565_));
 AND3x1_ASAP7_75t_R _27030_ (.A(_00155_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08566_));
 AOI211x1_ASAP7_75t_R _27031_ (.A1(_00154_),
    .A2(_07238_),
    .B(_08566_),
    .C(_07234_),
    .Y(_08567_));
 AO21x1_ASAP7_75t_R _27032_ (.A1(_02389_),
    .A2(_07234_),
    .B(_08567_),
    .Y(_08568_));
 OA21x2_ASAP7_75t_R _27033_ (.A1(_07073_),
    .A2(_07425_),
    .B(_08204_),
    .Y(_08569_));
 AO221x2_ASAP7_75t_R _27034_ (.A1(net2136),
    .A2(_07242_),
    .B1(_08568_),
    .B2(_07231_),
    .C(_08569_),
    .Y(_08570_));
 NAND2x1_ASAP7_75t_R _27035_ (.A(net308),
    .B(_08570_),
    .Y(_08571_));
 XNOR2x1_ASAP7_75t_R _27036_ (.B(_02252_),
    .Y(_08572_),
    .A(_00061_));
 AND2x2_ASAP7_75t_R _27037_ (.A(_07062_),
    .B(_08572_),
    .Y(_08573_));
 AO21x1_ASAP7_75t_R _27038_ (.A1(_07064_),
    .A2(_07995_),
    .B(_08573_),
    .Y(_08574_));
 AO221x1_ASAP7_75t_R _27039_ (.A1(_01242_),
    .A2(_07059_),
    .B1(_07060_),
    .B2(_08574_),
    .C(net308),
    .Y(_08575_));
 OA22x2_ASAP7_75t_R _27040_ (.A1(_01490_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01459_),
    .Y(_08576_));
 OA22x2_ASAP7_75t_R _27041_ (.A1(_02143_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02037_),
    .Y(_08577_));
 NAND2x1_ASAP7_75t_R _27042_ (.A(net3387),
    .B(_08134_),
    .Y(_08578_));
 OA22x2_ASAP7_75t_R _27043_ (.A1(_01966_),
    .A2(_07024_),
    .B1(_07369_),
    .B2(_01552_),
    .Y(_08579_));
 OA211x2_ASAP7_75t_R _27044_ (.A1(_02069_),
    .A2(_07026_),
    .B(_08578_),
    .C(_08579_),
    .Y(_08580_));
 OA21x2_ASAP7_75t_R _27045_ (.A1(_07021_),
    .A2(_08577_),
    .B(_08580_),
    .Y(_08581_));
 OA22x2_ASAP7_75t_R _27046_ (.A1(_02110_),
    .A2(_06992_),
    .B1(_06938_),
    .B2(_01916_),
    .Y(_08582_));
 OA21x2_ASAP7_75t_R _27047_ (.A1(_02000_),
    .A2(_07028_),
    .B(_07004_),
    .Y(_08583_));
 INVx1_ASAP7_75t_R _27048_ (.A(_00156_),
    .Y(_08584_));
 AO32x1_ASAP7_75t_R _27049_ (.A1(_08584_),
    .A2(_05612_),
    .A3(_05647_),
    .B1(_06942_),
    .B2(_06260_),
    .Y(_08585_));
 AOI22x1_ASAP7_75t_R _27050_ (.A1(net3607),
    .A2(_06947_),
    .B1(_08585_),
    .B2(_08213_),
    .Y(_08586_));
 OA211x2_ASAP7_75t_R _27051_ (.A1(_06990_),
    .A2(_08582_),
    .B(_08583_),
    .C(net3608),
    .Y(_08587_));
 OA211x2_ASAP7_75t_R _27052_ (.A1(_07360_),
    .A2(_08576_),
    .B(_08581_),
    .C(net3609),
    .Y(_08588_));
 AND4x1_ASAP7_75t_R _27053_ (.A(net290),
    .B(_08571_),
    .C(_08575_),
    .D(_08588_),
    .Y(_08589_));
 NOR2x1_ASAP7_75t_R _27054_ (.A(net432),
    .B(_08016_),
    .Y(_08590_));
 AO21x1_ASAP7_75t_R _27055_ (.A1(net432),
    .A2(_08018_),
    .B(_08590_),
    .Y(_08591_));
 AOI21x1_ASAP7_75t_R _27056_ (.A1(_07036_),
    .A2(_08591_),
    .B(_08113_),
    .Y(_08592_));
 AOI21x1_ASAP7_75t_R _27057_ (.A1(_08565_),
    .A2(_08589_),
    .B(_08592_),
    .Y(_08593_));
 NOR2x1_ASAP7_75t_R _27058_ (.A(_01680_),
    .B(net288),
    .Y(_08594_));
 AO21x1_ASAP7_75t_R _27059_ (.A1(net288),
    .A2(net250),
    .B(_08594_),
    .Y(_02685_));
 AND2x2_ASAP7_75t_R _27060_ (.A(_07077_),
    .B(_07342_),
    .Y(_08595_));
 OA22x2_ASAP7_75t_R _27061_ (.A1(_01489_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01458_),
    .Y(_08596_));
 OA22x2_ASAP7_75t_R _27062_ (.A1(_02142_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02036_),
    .Y(_08597_));
 OA22x2_ASAP7_75t_R _27063_ (.A1(_01915_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02109_),
    .Y(_08598_));
 NAND2x1_ASAP7_75t_R _27064_ (.A(net3695),
    .B(_07700_),
    .Y(_08599_));
 AND4x1_ASAP7_75t_R _27065_ (.A(_07791_),
    .B(_07000_),
    .C(_08598_),
    .D(net3696),
    .Y(_08600_));
 INVx1_ASAP7_75t_R _27066_ (.A(net3354),
    .Y(_08601_));
 OA222x2_ASAP7_75t_R _27067_ (.A1(_01999_),
    .A2(_07028_),
    .B1(_07369_),
    .B2(_01551_),
    .C1(_08601_),
    .C2(_07745_),
    .Y(_08602_));
 OA22x2_ASAP7_75t_R _27068_ (.A1(_02068_),
    .A2(_07026_),
    .B1(_07008_),
    .B2(_00159_),
    .Y(_08603_));
 OA22x2_ASAP7_75t_R _27069_ (.A1(_01965_),
    .A2(_07024_),
    .B1(_07522_),
    .B2(_01949_),
    .Y(_08604_));
 AND3x1_ASAP7_75t_R _27070_ (.A(_08602_),
    .B(_08603_),
    .C(_08604_),
    .Y(_08605_));
 OA211x2_ASAP7_75t_R _27071_ (.A1(_07021_),
    .A2(_08597_),
    .B(_08600_),
    .C(_08605_),
    .Y(_08606_));
 OAI21x1_ASAP7_75t_R _27072_ (.A1(_07360_),
    .A2(_08596_),
    .B(_08606_),
    .Y(_08607_));
 AND3x1_ASAP7_75t_R _27073_ (.A(_00158_),
    .B(_13618_),
    .C(_06635_),
    .Y(_08608_));
 AOI211x1_ASAP7_75t_R _27074_ (.A1(_00157_),
    .A2(_07238_),
    .B(_08608_),
    .C(_07234_),
    .Y(_08609_));
 AO21x1_ASAP7_75t_R _27075_ (.A1(_02390_),
    .A2(_07234_),
    .B(_08609_),
    .Y(_08610_));
 AO222x2_ASAP7_75t_R _27076_ (.A1(net172),
    .A2(_07242_),
    .B1(_07277_),
    .B2(_07215_),
    .C1(_08610_),
    .C2(_07231_),
    .Y(_08611_));
 NAND2x1_ASAP7_75t_R _27077_ (.A(_02255_),
    .B(_07062_),
    .Y(_08612_));
 OA211x2_ASAP7_75t_R _27078_ (.A1(_08044_),
    .A2(_07062_),
    .B(_08612_),
    .C(_07060_),
    .Y(_08613_));
 AO21x1_ASAP7_75t_R _27079_ (.A1(_01274_),
    .A2(_07059_),
    .B(_08613_),
    .Y(_08614_));
 NAND2x1_ASAP7_75t_R _27080_ (.A(_13817_),
    .B(_08614_),
    .Y(_08615_));
 OA21x2_ASAP7_75t_R _27081_ (.A1(_13817_),
    .A2(_08611_),
    .B(_08615_),
    .Y(_08616_));
 OR3x1_ASAP7_75t_R _27082_ (.A(_07474_),
    .B(_08607_),
    .C(_08616_),
    .Y(_08617_));
 OA211x2_ASAP7_75t_R _27083_ (.A1(net41),
    .A2(net434),
    .B(_08031_),
    .C(_07039_),
    .Y(_08618_));
 AO21x1_ASAP7_75t_R _27084_ (.A1(net432),
    .A2(_08029_),
    .B(_08618_),
    .Y(_08619_));
 AO21x2_ASAP7_75t_R _27085_ (.A1(_07036_),
    .A2(_08619_),
    .B(_08113_),
    .Y(_08620_));
 OA21x2_ASAP7_75t_R _27086_ (.A1(_08595_),
    .A2(_08617_),
    .B(_08620_),
    .Y(_08621_));
 NOR2x1_ASAP7_75t_R _27087_ (.A(_01679_),
    .B(_06987_),
    .Y(_08622_));
 AO21x1_ASAP7_75t_R _27088_ (.A1(_06987_),
    .A2(net2197),
    .B(_08622_),
    .Y(_02686_));
 AO221x1_ASAP7_75t_R _27089_ (.A1(_07073_),
    .A2(_07154_),
    .B1(_07196_),
    .B2(_07213_),
    .C(_07080_),
    .Y(_08623_));
 OAI22x1_ASAP7_75t_R _27090_ (.A1(_01488_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_01457_),
    .Y(_08624_));
 OAI22x1_ASAP7_75t_R _27091_ (.A1(_02141_),
    .A2(_07014_),
    .B1(_07016_),
    .B2(_02035_),
    .Y(_08625_));
 OAI22x1_ASAP7_75t_R _27092_ (.A1(_00161_),
    .A2(_07008_),
    .B1(_07369_),
    .B2(_01550_),
    .Y(_08626_));
 OAI22x1_ASAP7_75t_R _27093_ (.A1(_01964_),
    .A2(_07024_),
    .B1(_07028_),
    .B2(_01998_),
    .Y(_08627_));
 OAI22x1_ASAP7_75t_R _27094_ (.A1(_02067_),
    .A2(_05589_),
    .B1(_06990_),
    .B2(_01908_),
    .Y(_08628_));
 AO21x1_ASAP7_75t_R _27095_ (.A1(_07530_),
    .A2(_08628_),
    .B(_08057_),
    .Y(_08629_));
 OAI22x1_ASAP7_75t_R _27096_ (.A1(_01914_),
    .A2(_06998_),
    .B1(_07367_),
    .B2(_02108_),
    .Y(_08630_));
 AND2x2_ASAP7_75t_R _27097_ (.A(net3575),
    .B(_06947_),
    .Y(_08631_));
 OR5x2_ASAP7_75t_R _27098_ (.A(_08626_),
    .B(_08627_),
    .C(_08629_),
    .D(_08630_),
    .E(_08631_),
    .Y(_08632_));
 AOI221x1_ASAP7_75t_R _27099_ (.A1(_06950_),
    .A2(_08624_),
    .B1(_08625_),
    .B2(_06940_),
    .C(_08632_),
    .Y(_08633_));
 XNOR2x2_ASAP7_75t_R _27100_ (.A(_00064_),
    .B(_02254_),
    .Y(_08634_));
 NAND2x1_ASAP7_75t_R _27101_ (.A(_07062_),
    .B(_08634_),
    .Y(_08635_));
 OA211x2_ASAP7_75t_R _27102_ (.A1(_07062_),
    .A2(_08089_),
    .B(_08635_),
    .C(_07060_),
    .Y(_08636_));
 AO21x1_ASAP7_75t_R _27103_ (.A1(_05536_),
    .A2(_05766_),
    .B(net308),
    .Y(_08637_));
 OA211x2_ASAP7_75t_R _27104_ (.A1(_07219_),
    .A2(_07225_),
    .B(_07227_),
    .C(_07215_),
    .Y(_08638_));
 AND2x2_ASAP7_75t_R _27105_ (.A(_01310_),
    .B(_07238_),
    .Y(_08639_));
 AOI211x1_ASAP7_75t_R _27106_ (.A1(_00160_),
    .A2(_07237_),
    .B(_08639_),
    .C(_07234_),
    .Y(_08640_));
 AO21x1_ASAP7_75t_R _27107_ (.A1(_02282_),
    .A2(_07234_),
    .B(_08640_),
    .Y(_08641_));
 AO221x2_ASAP7_75t_R _27108_ (.A1(net173),
    .A2(_07242_),
    .B1(_08641_),
    .B2(_07231_),
    .C(_13817_),
    .Y(_08642_));
 OAI22x1_ASAP7_75t_R _27109_ (.A1(_08636_),
    .A2(_08637_),
    .B1(_08638_),
    .B2(_08642_),
    .Y(_08643_));
 AND3x1_ASAP7_75t_R _27110_ (.A(_06981_),
    .B(_08633_),
    .C(_08643_),
    .Y(_08644_));
 NAND2x1_ASAP7_75t_R _27111_ (.A(_01642_),
    .B(_08077_),
    .Y(_08645_));
 OA211x2_ASAP7_75t_R _27112_ (.A1(_01642_),
    .A2(_08076_),
    .B(_08645_),
    .C(_07036_),
    .Y(_08646_));
 NOR2x2_ASAP7_75t_R _27113_ (.A(_08113_),
    .B(_08646_),
    .Y(_08647_));
 AO21x2_ASAP7_75t_R _27114_ (.A1(_08623_),
    .A2(_08644_),
    .B(_08647_),
    .Y(_08648_));
 TAPCELL_ASAP7_75t_R PHY_681 ();
 NAND2x1_ASAP7_75t_R _27116_ (.A(_06987_),
    .B(_08648_),
    .Y(_08650_));
 OA21x2_ASAP7_75t_R _27117_ (.A1(_05481_),
    .A2(_06987_),
    .B(_08650_),
    .Y(_02687_));
 NAND2x2_ASAP7_75t_R _27118_ (.A(_01873_),
    .B(_13771_),
    .Y(_08651_));
 AND2x2_ASAP7_75t_R _27119_ (.A(_05513_),
    .B(_05950_),
    .Y(_08652_));
 NAND2x2_ASAP7_75t_R _27120_ (.A(_13604_),
    .B(_07059_),
    .Y(_08653_));
 OR2x2_ASAP7_75t_R _27121_ (.A(_01519_),
    .B(_05547_),
    .Y(_08654_));
 NAND2x2_ASAP7_75t_R _27122_ (.A(_05513_),
    .B(_05950_),
    .Y(_08655_));
 AND4x1_ASAP7_75t_R _27123_ (.A(_13604_),
    .B(_07059_),
    .C(_05944_),
    .D(_08655_),
    .Y(_08656_));
 AO21x1_ASAP7_75t_R _27124_ (.A1(_06752_),
    .A2(_08652_),
    .B(_08656_),
    .Y(_08657_));
 AO221x1_ASAP7_75t_R _27125_ (.A1(_08652_),
    .A2(_08653_),
    .B1(_08654_),
    .B2(_08657_),
    .C(_00285_),
    .Y(_08658_));
 OA21x2_ASAP7_75t_R _27126_ (.A1(_05782_),
    .A2(_08651_),
    .B(_08658_),
    .Y(_08659_));
 OA21x2_ASAP7_75t_R _27127_ (.A1(_07060_),
    .A2(_08659_),
    .B(_14843_),
    .Y(_08660_));
 TAPCELL_ASAP7_75t_R PHY_680 ();
 TAPCELL_ASAP7_75t_R PHY_679 ();
 TAPCELL_ASAP7_75t_R PHY_678 ();
 NOR2x2_ASAP7_75t_R _27131_ (.A(_05547_),
    .B(_08653_),
    .Y(_08664_));
 OR3x4_ASAP7_75t_R _27132_ (.A(_07060_),
    .B(_08651_),
    .C(_08664_),
    .Y(_08665_));
 TAPCELL_ASAP7_75t_R PHY_677 ();
 TAPCELL_ASAP7_75t_R PHY_676 ();
 AND2x6_ASAP7_75t_R _27135_ (.A(_01873_),
    .B(_13771_),
    .Y(_08668_));
 NOR2x1_ASAP7_75t_R _27136_ (.A(_02291_),
    .B(_05771_),
    .Y(_08669_));
 XNOR2x2_ASAP7_75t_R _27137_ (.A(_01318_),
    .B(_08669_),
    .Y(_08670_));
 XNOR2x2_ASAP7_75t_R _27138_ (.A(_01322_),
    .B(_02292_),
    .Y(_08671_));
 INVx2_ASAP7_75t_R _27139_ (.A(_08671_),
    .Y(_08672_));
 TAPCELL_ASAP7_75t_R PHY_675 ();
 TAPCELL_ASAP7_75t_R PHY_674 ();
 INVx1_ASAP7_75t_R _27142_ (.A(_01673_),
    .Y(_08675_));
 TAPCELL_ASAP7_75t_R PHY_673 ();
 NOR2x1_ASAP7_75t_R _27144_ (.A(net314),
    .B(_01675_),
    .Y(_08677_));
 AO21x1_ASAP7_75t_R _27145_ (.A1(net314),
    .A2(_08675_),
    .B(_08677_),
    .Y(_08678_));
 INVx1_ASAP7_75t_R _27146_ (.A(_01676_),
    .Y(_08679_));
 TAPCELL_ASAP7_75t_R PHY_672 ();
 NAND2x1_ASAP7_75t_R _27148_ (.A(net314),
    .B(_01674_),
    .Y(_08681_));
 OA211x2_ASAP7_75t_R _27149_ (.A1(net314),
    .A2(_08679_),
    .B(_08681_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08682_));
 AO21x1_ASAP7_75t_R _27150_ (.A1(_17818_),
    .A2(_08678_),
    .B(_08682_),
    .Y(_08683_));
 INVx1_ASAP7_75t_R _27151_ (.A(_01668_),
    .Y(_08684_));
 NAND2x1_ASAP7_75t_R _27152_ (.A(net313),
    .B(_01666_),
    .Y(_08685_));
 OA211x2_ASAP7_75t_R _27153_ (.A1(net313),
    .A2(_08684_),
    .B(_08685_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08686_));
 INVx1_ASAP7_75t_R _27154_ (.A(_01667_),
    .Y(_08687_));
 NAND2x1_ASAP7_75t_R _27155_ (.A(net314),
    .B(_01665_),
    .Y(_08688_));
 OA211x2_ASAP7_75t_R _27156_ (.A1(net314),
    .A2(_08687_),
    .B(_08688_),
    .C(_17818_),
    .Y(_08689_));
 OR3x1_ASAP7_75t_R _27157_ (.A(_08671_),
    .B(_08686_),
    .C(_08689_),
    .Y(_08690_));
 INVx1_ASAP7_75t_R _27158_ (.A(_02293_),
    .Y(_08691_));
 OA211x2_ASAP7_75t_R _27159_ (.A1(_08672_),
    .A2(_08683_),
    .B(_08690_),
    .C(_08691_),
    .Y(_08692_));
 INVx1_ASAP7_75t_R _27160_ (.A(_01672_),
    .Y(_08693_));
 NAND2x1_ASAP7_75t_R _27161_ (.A(net313),
    .B(_01670_),
    .Y(_08694_));
 OA211x2_ASAP7_75t_R _27162_ (.A1(net313),
    .A2(_08693_),
    .B(_08694_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08695_));
 INVx1_ASAP7_75t_R _27163_ (.A(_01671_),
    .Y(_08696_));
 NAND2x1_ASAP7_75t_R _27164_ (.A(net314),
    .B(_01669_),
    .Y(_08697_));
 OA211x2_ASAP7_75t_R _27165_ (.A1(net314),
    .A2(_08696_),
    .B(_08697_),
    .C(_17818_),
    .Y(_08698_));
 OR3x1_ASAP7_75t_R _27166_ (.A(_08672_),
    .B(_08695_),
    .C(_08698_),
    .Y(_08699_));
 INVx1_ASAP7_75t_R _27167_ (.A(_01664_),
    .Y(_08700_));
 NAND2x1_ASAP7_75t_R _27168_ (.A(net313),
    .B(_01662_),
    .Y(_08701_));
 OA211x2_ASAP7_75t_R _27169_ (.A1(net313),
    .A2(_08700_),
    .B(_08701_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08702_));
 INVx1_ASAP7_75t_R _27170_ (.A(_01663_),
    .Y(_08703_));
 NAND2x1_ASAP7_75t_R _27171_ (.A(net314),
    .B(_01661_),
    .Y(_08704_));
 OA211x2_ASAP7_75t_R _27172_ (.A1(net314),
    .A2(_08703_),
    .B(_08704_),
    .C(_17818_),
    .Y(_08705_));
 OR3x1_ASAP7_75t_R _27173_ (.A(_08671_),
    .B(_08702_),
    .C(_08705_),
    .Y(_08706_));
 AND3x1_ASAP7_75t_R _27174_ (.A(_02293_),
    .B(_08699_),
    .C(_08706_),
    .Y(_08707_));
 NOR2x1_ASAP7_75t_R _27175_ (.A(_08692_),
    .B(_08707_),
    .Y(_08708_));
 INVx1_ASAP7_75t_R _27176_ (.A(_01660_),
    .Y(_08709_));
 NAND2x1_ASAP7_75t_R _27177_ (.A(net313),
    .B(_01658_),
    .Y(_08710_));
 OA211x2_ASAP7_75t_R _27178_ (.A1(net313),
    .A2(_08709_),
    .B(_08710_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08711_));
 INVx1_ASAP7_75t_R _27179_ (.A(_01659_),
    .Y(_08712_));
 NAND2x1_ASAP7_75t_R _27180_ (.A(net313),
    .B(_01657_),
    .Y(_08713_));
 OA211x2_ASAP7_75t_R _27181_ (.A1(net313),
    .A2(_08712_),
    .B(_08713_),
    .C(_17818_),
    .Y(_08714_));
 OR3x1_ASAP7_75t_R _27182_ (.A(_08672_),
    .B(_08711_),
    .C(_08714_),
    .Y(_08715_));
 INVx1_ASAP7_75t_R _27183_ (.A(_01652_),
    .Y(_08716_));
 NAND2x1_ASAP7_75t_R _27184_ (.A(net313),
    .B(_01650_),
    .Y(_08717_));
 OA211x2_ASAP7_75t_R _27185_ (.A1(net313),
    .A2(_08716_),
    .B(_08717_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08718_));
 INVx1_ASAP7_75t_R _27186_ (.A(_01651_),
    .Y(_08719_));
 NAND2x1_ASAP7_75t_R _27187_ (.A(net313),
    .B(_01649_),
    .Y(_08720_));
 OA211x2_ASAP7_75t_R _27188_ (.A1(net313),
    .A2(_08719_),
    .B(_08720_),
    .C(_17818_),
    .Y(_08721_));
 OR3x1_ASAP7_75t_R _27189_ (.A(_08671_),
    .B(_08718_),
    .C(_08721_),
    .Y(_08722_));
 AND3x1_ASAP7_75t_R _27190_ (.A(_08691_),
    .B(_08715_),
    .C(_08722_),
    .Y(_08723_));
 INVx1_ASAP7_75t_R _27191_ (.A(_01648_),
    .Y(_08724_));
 NAND2x1_ASAP7_75t_R _27192_ (.A(net314),
    .B(_01646_),
    .Y(_08725_));
 OA211x2_ASAP7_75t_R _27193_ (.A1(net314),
    .A2(_08724_),
    .B(_08725_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08726_));
 INVx1_ASAP7_75t_R _27194_ (.A(_01647_),
    .Y(_08727_));
 NAND2x1_ASAP7_75t_R _27195_ (.A(net313),
    .B(_01645_),
    .Y(_08728_));
 OA211x2_ASAP7_75t_R _27196_ (.A1(net313),
    .A2(_08727_),
    .B(_08728_),
    .C(_17818_),
    .Y(_08729_));
 OR3x1_ASAP7_75t_R _27197_ (.A(_08671_),
    .B(_08726_),
    .C(_08729_),
    .Y(_08730_));
 INVx1_ASAP7_75t_R _27198_ (.A(_01656_),
    .Y(_08731_));
 NAND2x1_ASAP7_75t_R _27199_ (.A(net314),
    .B(_01654_),
    .Y(_08732_));
 OA211x2_ASAP7_75t_R _27200_ (.A1(net314),
    .A2(_08731_),
    .B(_08732_),
    .C(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .Y(_08733_));
 INVx1_ASAP7_75t_R _27201_ (.A(_01655_),
    .Y(_08734_));
 NAND2x1_ASAP7_75t_R _27202_ (.A(net314),
    .B(_01653_),
    .Y(_08735_));
 OA211x2_ASAP7_75t_R _27203_ (.A1(net314),
    .A2(_08734_),
    .B(_08735_),
    .C(_17818_),
    .Y(_08736_));
 OR3x1_ASAP7_75t_R _27204_ (.A(_08672_),
    .B(_08733_),
    .C(_08736_),
    .Y(_08737_));
 AND3x1_ASAP7_75t_R _27205_ (.A(_02293_),
    .B(_08730_),
    .C(_08737_),
    .Y(_08738_));
 OAI21x1_ASAP7_75t_R _27206_ (.A1(_08723_),
    .A2(_08738_),
    .B(_08670_),
    .Y(_08739_));
 OA21x2_ASAP7_75t_R _27207_ (.A1(_08670_),
    .A2(_08708_),
    .B(_08739_),
    .Y(_08740_));
 NOR2x1_ASAP7_75t_R _27208_ (.A(_01357_),
    .B(_08740_),
    .Y(_08741_));
 INVx1_ASAP7_75t_R _27209_ (.A(_01645_),
    .Y(_08742_));
 AO22x1_ASAP7_75t_R _27210_ (.A1(_13775_),
    .A2(\ex_block_i.alu_adder_result_ex_o[0] ),
    .B1(_08742_),
    .B2(_05776_),
    .Y(_08743_));
 OR3x4_ASAP7_75t_R _27211_ (.A(_00279_),
    .B(_13559_),
    .C(_13538_),
    .Y(_08744_));
 INVx1_ASAP7_75t_R _27212_ (.A(_02202_),
    .Y(_08745_));
 MAJx3_ASAP7_75t_R _27213_ (.A(_01308_),
    .B(_08745_),
    .C(net173),
    .Y(_08746_));
 TAPCELL_ASAP7_75t_R PHY_671 ();
 MAJx3_ASAP7_75t_R _27215_ (.A(_05536_),
    .B(_02202_),
    .C(_05542_),
    .Y(_08748_));
 AND2x2_ASAP7_75t_R _27216_ (.A(_16721_),
    .B(_08748_),
    .Y(_08749_));
 AO21x1_ASAP7_75t_R _27217_ (.A1(_00324_),
    .A2(_08746_),
    .B(_08749_),
    .Y(_08750_));
 TAPCELL_ASAP7_75t_R PHY_670 ();
 OR3x4_ASAP7_75t_R _27219_ (.A(_05773_),
    .B(_05771_),
    .C(_08746_),
    .Y(_08752_));
 OA211x2_ASAP7_75t_R _27220_ (.A1(_01321_),
    .A2(_08752_),
    .B(_08664_),
    .C(_01323_),
    .Y(_08753_));
 AOI211x1_ASAP7_75t_R _27221_ (.A1(_08744_),
    .A2(_08750_),
    .B(_01727_),
    .C(_08753_),
    .Y(_08754_));
 OR5x2_ASAP7_75t_R _27222_ (.A(_07060_),
    .B(_08668_),
    .C(_08741_),
    .D(_08743_),
    .E(_08754_),
    .Y(_08755_));
 NAND2x1_ASAP7_75t_R _27223_ (.A(_00324_),
    .B(_07064_),
    .Y(_08756_));
 TAPCELL_ASAP7_75t_R PHY_669 ();
 NAND2x1_ASAP7_75t_R _27225_ (.A(_01356_),
    .B(_07062_),
    .Y(_08758_));
 AO21x1_ASAP7_75t_R _27226_ (.A1(_08756_),
    .A2(_08758_),
    .B(_05766_),
    .Y(_08759_));
 OA211x2_ASAP7_75t_R _27227_ (.A1(_13981_),
    .A2(_08665_),
    .B(_08755_),
    .C(_08759_),
    .Y(_08760_));
 TAPCELL_ASAP7_75t_R PHY_668 ();
 NOR2x1_ASAP7_75t_R _27229_ (.A(_00324_),
    .B(_08660_),
    .Y(_08762_));
 AO21x1_ASAP7_75t_R _27230_ (.A1(_08660_),
    .A2(_08760_),
    .B(_08762_),
    .Y(_02688_));
 NAND2x1_ASAP7_75t_R _27231_ (.A(_00291_),
    .B(_07064_),
    .Y(_08763_));
 NAND2x1_ASAP7_75t_R _27232_ (.A(_01360_),
    .B(_07062_),
    .Y(_08764_));
 AO21x1_ASAP7_75t_R _27233_ (.A1(_08763_),
    .A2(_08764_),
    .B(_05766_),
    .Y(_08765_));
 TAPCELL_ASAP7_75t_R PHY_667 ();
 TAPCELL_ASAP7_75t_R PHY_666 ();
 OR3x1_ASAP7_75t_R _27236_ (.A(_05771_),
    .B(_05774_),
    .C(_08746_),
    .Y(_08768_));
 TAPCELL_ASAP7_75t_R PHY_665 ();
 TAPCELL_ASAP7_75t_R PHY_664 ();
 AND2x2_ASAP7_75t_R _27239_ (.A(_16717_),
    .B(_08748_),
    .Y(_08771_));
 AO21x1_ASAP7_75t_R _27240_ (.A1(_00291_),
    .A2(_08746_),
    .B(_08771_),
    .Y(_08772_));
 TAPCELL_ASAP7_75t_R PHY_663 ();
 AO32x1_ASAP7_75t_R _27242_ (.A1(_01324_),
    .A2(_08664_),
    .A3(_08768_),
    .B1(_08772_),
    .B2(_08744_),
    .Y(_08774_));
 TAPCELL_ASAP7_75t_R PHY_662 ();
 TAPCELL_ASAP7_75t_R PHY_661 ();
 AND2x6_ASAP7_75t_R _27245_ (.A(_05766_),
    .B(_08651_),
    .Y(_08777_));
 OA21x2_ASAP7_75t_R _27246_ (.A1(_00285_),
    .A2(_16717_),
    .B(_08777_),
    .Y(_08778_));
 OA21x2_ASAP7_75t_R _27247_ (.A1(_01357_),
    .A2(_08750_),
    .B(_08778_),
    .Y(_08779_));
 OAI21x1_ASAP7_75t_R _27248_ (.A1(_01727_),
    .A2(_08774_),
    .B(_08779_),
    .Y(_08780_));
 OA211x2_ASAP7_75t_R _27249_ (.A1(_13767_),
    .A2(_08665_),
    .B(_08765_),
    .C(_08780_),
    .Y(_08781_));
 NOR2x1_ASAP7_75t_R _27250_ (.A(_00291_),
    .B(_08660_),
    .Y(_08782_));
 AO21x1_ASAP7_75t_R _27251_ (.A1(_08660_),
    .A2(_08781_),
    .B(_08782_),
    .Y(_02689_));
 NAND2x1_ASAP7_75t_R _27252_ (.A(_00663_),
    .B(_07064_),
    .Y(_08783_));
 NAND2x1_ASAP7_75t_R _27253_ (.A(_01364_),
    .B(_07062_),
    .Y(_08784_));
 AO21x1_ASAP7_75t_R _27254_ (.A1(_08783_),
    .A2(_08784_),
    .B(_05766_),
    .Y(_08785_));
 OA211x2_ASAP7_75t_R _27255_ (.A1(_01326_),
    .A2(_08752_),
    .B(_08664_),
    .C(_01325_),
    .Y(_08786_));
 TAPCELL_ASAP7_75t_R PHY_660 ();
 AND2x2_ASAP7_75t_R _27257_ (.A(_05792_),
    .B(_08748_),
    .Y(_08788_));
 AO21x1_ASAP7_75t_R _27258_ (.A1(_00663_),
    .A2(_08746_),
    .B(_08788_),
    .Y(_08789_));
 TAPCELL_ASAP7_75t_R PHY_659 ();
 AO21x1_ASAP7_75t_R _27260_ (.A1(_08744_),
    .A2(_08789_),
    .B(_01727_),
    .Y(_08791_));
 OA21x2_ASAP7_75t_R _27261_ (.A1(_00285_),
    .A2(_05792_),
    .B(_08777_),
    .Y(_08792_));
 OA21x2_ASAP7_75t_R _27262_ (.A1(_01357_),
    .A2(_08772_),
    .B(_08792_),
    .Y(_08793_));
 OAI21x1_ASAP7_75t_R _27263_ (.A1(_08786_),
    .A2(_08791_),
    .B(_08793_),
    .Y(_08794_));
 OA211x2_ASAP7_75t_R _27264_ (.A1(_14921_),
    .A2(_08665_),
    .B(_08785_),
    .C(_08794_),
    .Y(_08795_));
 NOR2x1_ASAP7_75t_R _27265_ (.A(_00663_),
    .B(_08660_),
    .Y(_08796_));
 AO21x1_ASAP7_75t_R _27266_ (.A1(_08660_),
    .A2(_08795_),
    .B(_08796_),
    .Y(_02690_));
 TAPCELL_ASAP7_75t_R PHY_658 ();
 CKINVDCx10_ASAP7_75t_R _27268_ (.A(_08660_),
    .Y(_08798_));
 TAPCELL_ASAP7_75t_R PHY_657 ();
 NAND2x1_ASAP7_75t_R _27270_ (.A(_02231_),
    .B(_07062_),
    .Y(_08800_));
 TAPCELL_ASAP7_75t_R PHY_656 ();
 OA211x2_ASAP7_75t_R _27272_ (.A1(_00665_),
    .A2(_07062_),
    .B(_08800_),
    .C(_07060_),
    .Y(_08802_));
 NOR2x1_ASAP7_75t_R _27273_ (.A(_14980_),
    .B(_08665_),
    .Y(_08803_));
 AND2x2_ASAP7_75t_R _27274_ (.A(_06317_),
    .B(_08748_),
    .Y(_08804_));
 AO21x1_ASAP7_75t_R _27275_ (.A1(_00665_),
    .A2(_08746_),
    .B(_08804_),
    .Y(_08805_));
 AND3x4_ASAP7_75t_R _27276_ (.A(_13570_),
    .B(_00282_),
    .C(_13817_),
    .Y(_08806_));
 OA211x2_ASAP7_75t_R _27277_ (.A1(_01320_),
    .A2(_08752_),
    .B(_08806_),
    .C(_01327_),
    .Y(_08807_));
 AO21x1_ASAP7_75t_R _27278_ (.A1(_08744_),
    .A2(_08805_),
    .B(_08807_),
    .Y(_08808_));
 OA21x2_ASAP7_75t_R _27279_ (.A1(_00285_),
    .A2(_06317_),
    .B(_08777_),
    .Y(_08809_));
 OA21x2_ASAP7_75t_R _27280_ (.A1(_01357_),
    .A2(_08789_),
    .B(_08809_),
    .Y(_08810_));
 OA21x2_ASAP7_75t_R _27281_ (.A1(_01727_),
    .A2(_08808_),
    .B(_08810_),
    .Y(_08811_));
 OR4x1_ASAP7_75t_R _27282_ (.A(_08798_),
    .B(_08802_),
    .C(_08803_),
    .D(_08811_),
    .Y(_08812_));
 OAI21x1_ASAP7_75t_R _27283_ (.A1(_00665_),
    .A2(_08660_),
    .B(_08812_),
    .Y(_02691_));
 TAPCELL_ASAP7_75t_R PHY_655 ();
 TAPCELL_ASAP7_75t_R PHY_654 ();
 TAPCELL_ASAP7_75t_R PHY_653 ();
 TAPCELL_ASAP7_75t_R PHY_652 ();
 AND2x2_ASAP7_75t_R _27288_ (.A(_05791_),
    .B(_08748_),
    .Y(_08817_));
 AO21x1_ASAP7_75t_R _27289_ (.A1(_00668_),
    .A2(_08746_),
    .B(_08817_),
    .Y(_08818_));
 INVx2_ASAP7_75t_R _27290_ (.A(_01322_),
    .Y(_08819_));
 TAPCELL_ASAP7_75t_R PHY_651 ();
 OR3x2_ASAP7_75t_R _27292_ (.A(_08819_),
    .B(_17825_),
    .C(_08746_),
    .Y(_08821_));
 OR2x4_ASAP7_75t_R _27293_ (.A(_05773_),
    .B(_08821_),
    .Y(_08822_));
 OA211x2_ASAP7_75t_R _27294_ (.A1(_01321_),
    .A2(_08822_),
    .B(_08664_),
    .C(_01328_),
    .Y(_08823_));
 AOI211x1_ASAP7_75t_R _27295_ (.A1(_08744_),
    .A2(_08818_),
    .B(_08823_),
    .C(_01727_),
    .Y(_08824_));
 TAPCELL_ASAP7_75t_R PHY_650 ();
 TAPCELL_ASAP7_75t_R PHY_649 ();
 OA21x2_ASAP7_75t_R _27298_ (.A1(_00285_),
    .A2(_05791_),
    .B(_08777_),
    .Y(_08827_));
 OAI21x1_ASAP7_75t_R _27299_ (.A1(_01357_),
    .A2(_08805_),
    .B(_08827_),
    .Y(_08828_));
 NAND2x1_ASAP7_75t_R _27300_ (.A(_01376_),
    .B(_07062_),
    .Y(_08829_));
 OA21x2_ASAP7_75t_R _27301_ (.A1(_06760_),
    .A2(_07062_),
    .B(_08829_),
    .Y(_08830_));
 OA22x2_ASAP7_75t_R _27302_ (.A1(net2322),
    .A2(_08665_),
    .B1(_08830_),
    .B2(_05766_),
    .Y(_08831_));
 OA211x2_ASAP7_75t_R _27303_ (.A1(_08824_),
    .A2(_08828_),
    .B(_08660_),
    .C(_08831_),
    .Y(_08832_));
 AO21x1_ASAP7_75t_R _27304_ (.A1(_06760_),
    .A2(_08798_),
    .B(_08832_),
    .Y(_02692_));
 OA21x2_ASAP7_75t_R _27305_ (.A1(_00285_),
    .A2(_06345_),
    .B(_08777_),
    .Y(_08833_));
 OAI21x1_ASAP7_75t_R _27306_ (.A1(_01357_),
    .A2(_08818_),
    .B(_08833_),
    .Y(_08834_));
 AND2x2_ASAP7_75t_R _27307_ (.A(_06345_),
    .B(_08748_),
    .Y(_08835_));
 AO21x1_ASAP7_75t_R _27308_ (.A1(_00670_),
    .A2(_08746_),
    .B(_08835_),
    .Y(_08836_));
 OA211x2_ASAP7_75t_R _27309_ (.A1(_05774_),
    .A2(_08821_),
    .B(_08664_),
    .C(_01329_),
    .Y(_08837_));
 AOI211x1_ASAP7_75t_R _27310_ (.A1(_08744_),
    .A2(_08836_),
    .B(_08837_),
    .C(_01727_),
    .Y(_08838_));
 AND2x2_ASAP7_75t_R _27311_ (.A(_07062_),
    .B(_07639_),
    .Y(_08839_));
 AO21x1_ASAP7_75t_R _27312_ (.A1(_15105_),
    .A2(_07064_),
    .B(_08839_),
    .Y(_08840_));
 OA222x2_ASAP7_75t_R _27313_ (.A1(_15103_),
    .A2(_08665_),
    .B1(_08834_),
    .B2(_08838_),
    .C1(_08840_),
    .C2(_05766_),
    .Y(_08841_));
 NOR2x1_ASAP7_75t_R _27314_ (.A(_00670_),
    .B(_08660_),
    .Y(_08842_));
 AO21x1_ASAP7_75t_R _27315_ (.A1(_08660_),
    .A2(_08841_),
    .B(_08842_),
    .Y(_02693_));
 TAPCELL_ASAP7_75t_R PHY_648 ();
 TAPCELL_ASAP7_75t_R PHY_647 ();
 AND2x2_ASAP7_75t_R _27318_ (.A(_05793_),
    .B(_08748_),
    .Y(_08845_));
 AO21x1_ASAP7_75t_R _27319_ (.A1(_00672_),
    .A2(_08746_),
    .B(_08845_),
    .Y(_08846_));
 TAPCELL_ASAP7_75t_R PHY_646 ();
 OA211x2_ASAP7_75t_R _27321_ (.A1(_01326_),
    .A2(_08822_),
    .B(_08806_),
    .C(_01330_),
    .Y(_08848_));
 AO21x1_ASAP7_75t_R _27322_ (.A1(_08744_),
    .A2(_08846_),
    .B(_08848_),
    .Y(_08849_));
 AND3x4_ASAP7_75t_R _27323_ (.A(_14843_),
    .B(_05766_),
    .C(_08659_),
    .Y(_08850_));
 OR2x6_ASAP7_75t_R _27324_ (.A(_08651_),
    .B(_08664_),
    .Y(_08851_));
 TAPCELL_ASAP7_75t_R PHY_645 ();
 TAPCELL_ASAP7_75t_R PHY_644 ();
 OA21x2_ASAP7_75t_R _27327_ (.A1(_00285_),
    .A2(_05793_),
    .B(_08651_),
    .Y(_08854_));
 OAI21x1_ASAP7_75t_R _27328_ (.A1(_01357_),
    .A2(_08836_),
    .B(_08854_),
    .Y(_08855_));
 OAI21x1_ASAP7_75t_R _27329_ (.A1(_15167_),
    .A2(_08851_),
    .B(_08855_),
    .Y(_08856_));
 OA211x2_ASAP7_75t_R _27330_ (.A1(_01727_),
    .A2(_08849_),
    .B(_08850_),
    .C(_08856_),
    .Y(_08857_));
 NAND2x1_ASAP7_75t_R _27331_ (.A(_07062_),
    .B(_08660_),
    .Y(_08858_));
 AO32x1_ASAP7_75t_R _27332_ (.A1(_07684_),
    .A2(_14843_),
    .A3(_07519_),
    .B1(_08858_),
    .B2(_00672_),
    .Y(_08859_));
 NOR2x1_ASAP7_75t_R _27333_ (.A(_08857_),
    .B(_08859_),
    .Y(_02694_));
 OA211x2_ASAP7_75t_R _27334_ (.A1(_01320_),
    .A2(_08822_),
    .B(_08664_),
    .C(_01331_),
    .Y(_08860_));
 AND2x2_ASAP7_75t_R _27335_ (.A(_00676_),
    .B(_08748_),
    .Y(_08861_));
 AO21x1_ASAP7_75t_R _27336_ (.A1(_00674_),
    .A2(_08746_),
    .B(_08861_),
    .Y(_08862_));
 AO21x1_ASAP7_75t_R _27337_ (.A1(_08744_),
    .A2(_08862_),
    .B(_01727_),
    .Y(_08863_));
 OA21x2_ASAP7_75t_R _27338_ (.A1(_00285_),
    .A2(_00676_),
    .B(_08777_),
    .Y(_08864_));
 OA21x2_ASAP7_75t_R _27339_ (.A1(_01357_),
    .A2(_08846_),
    .B(_08864_),
    .Y(_08865_));
 OA21x2_ASAP7_75t_R _27340_ (.A1(_08860_),
    .A2(_08863_),
    .B(_08865_),
    .Y(_08866_));
 NOR2x1_ASAP7_75t_R _27341_ (.A(_07060_),
    .B(_08851_),
    .Y(_08867_));
 AO21x1_ASAP7_75t_R _27342_ (.A1(_05885_),
    .A2(_08867_),
    .B(_07730_),
    .Y(_08868_));
 OR3x1_ASAP7_75t_R _27343_ (.A(_08798_),
    .B(_08866_),
    .C(_08868_),
    .Y(_08869_));
 OAI21x1_ASAP7_75t_R _27344_ (.A1(_00674_),
    .A2(_08660_),
    .B(_08869_),
    .Y(_02695_));
 AND2x2_ASAP7_75t_R _27345_ (.A(_05798_),
    .B(_08748_),
    .Y(_08870_));
 AO21x1_ASAP7_75t_R _27346_ (.A1(_00677_),
    .A2(_08746_),
    .B(_08870_),
    .Y(_08871_));
 INVx1_ASAP7_75t_R _27347_ (.A(_17825_),
    .Y(_08872_));
 NAND2x2_ASAP7_75t_R _27348_ (.A(_01318_),
    .B(_08819_),
    .Y(_08873_));
 OR3x4_ASAP7_75t_R _27349_ (.A(_08872_),
    .B(_08746_),
    .C(_08873_),
    .Y(_08874_));
 OA211x2_ASAP7_75t_R _27350_ (.A1(_01321_),
    .A2(_08874_),
    .B(_08664_),
    .C(_01332_),
    .Y(_08875_));
 AO21x1_ASAP7_75t_R _27351_ (.A1(_08744_),
    .A2(_08871_),
    .B(_08875_),
    .Y(_08876_));
 OA211x2_ASAP7_75t_R _27352_ (.A1(_00285_),
    .A2(_05798_),
    .B(_08651_),
    .C(_08850_),
    .Y(_08877_));
 OA21x2_ASAP7_75t_R _27353_ (.A1(_01357_),
    .A2(_08862_),
    .B(_08877_),
    .Y(_08878_));
 OA21x2_ASAP7_75t_R _27354_ (.A1(_01727_),
    .A2(_08876_),
    .B(_08878_),
    .Y(_08879_));
 NOR2x1_ASAP7_75t_R _27355_ (.A(_15279_),
    .B(_08851_),
    .Y(_08880_));
 AO32x1_ASAP7_75t_R _27356_ (.A1(_07763_),
    .A2(_14843_),
    .A3(_07519_),
    .B1(_08850_),
    .B2(_08880_),
    .Y(_08881_));
 AOI211x1_ASAP7_75t_R _27357_ (.A1(_00677_),
    .A2(_08858_),
    .B(_08879_),
    .C(_08881_),
    .Y(_02696_));
 AND2x2_ASAP7_75t_R _27358_ (.A(_06391_),
    .B(_08748_),
    .Y(_08882_));
 AO21x1_ASAP7_75t_R _27359_ (.A1(_00680_),
    .A2(_08746_),
    .B(_08882_),
    .Y(_08883_));
 NAND2x2_ASAP7_75t_R _27360_ (.A(_17825_),
    .B(_08748_),
    .Y(_08884_));
 OR3x1_ASAP7_75t_R _27361_ (.A(_01322_),
    .B(_05774_),
    .C(_08884_),
    .Y(_08885_));
 AND3x1_ASAP7_75t_R _27362_ (.A(_01333_),
    .B(_08806_),
    .C(_08885_),
    .Y(_08886_));
 AOI211x1_ASAP7_75t_R _27363_ (.A1(_08744_),
    .A2(_08883_),
    .B(_08886_),
    .C(_01727_),
    .Y(_08887_));
 OA21x2_ASAP7_75t_R _27364_ (.A1(_00285_),
    .A2(_06391_),
    .B(_08777_),
    .Y(_08888_));
 OAI21x1_ASAP7_75t_R _27365_ (.A1(_01357_),
    .A2(_08871_),
    .B(_08888_),
    .Y(_08889_));
 OR3x1_ASAP7_75t_R _27366_ (.A(_15282_),
    .B(_05815_),
    .C(_07061_),
    .Y(_08890_));
 OA21x2_ASAP7_75t_R _27367_ (.A1(_07064_),
    .A2(_07837_),
    .B(_08890_),
    .Y(_08891_));
 OA222x2_ASAP7_75t_R _27368_ (.A1(_15331_),
    .A2(_08665_),
    .B1(_08887_),
    .B2(_08889_),
    .C1(_08891_),
    .C2(_05766_),
    .Y(_08892_));
 NOR2x1_ASAP7_75t_R _27369_ (.A(_00680_),
    .B(_08660_),
    .Y(_08893_));
 AO21x1_ASAP7_75t_R _27370_ (.A1(_08660_),
    .A2(_08892_),
    .B(_08893_),
    .Y(_02697_));
 OR2x2_ASAP7_75t_R _27371_ (.A(_00682_),
    .B(_08748_),
    .Y(_08894_));
 NAND2x1_ASAP7_75t_R _27372_ (.A(net151),
    .B(_08748_),
    .Y(_08895_));
 AND3x1_ASAP7_75t_R _27373_ (.A(_08744_),
    .B(_08894_),
    .C(_08895_),
    .Y(_08896_));
 OA211x2_ASAP7_75t_R _27374_ (.A1(_01326_),
    .A2(_08874_),
    .B(_08806_),
    .C(_01334_),
    .Y(_08897_));
 OR3x1_ASAP7_75t_R _27375_ (.A(_01727_),
    .B(_08896_),
    .C(_08897_),
    .Y(_08898_));
 OA21x2_ASAP7_75t_R _27376_ (.A1(_00285_),
    .A2(_05797_),
    .B(_08777_),
    .Y(_08899_));
 OA211x2_ASAP7_75t_R _27377_ (.A1(_01357_),
    .A2(_08883_),
    .B(_08898_),
    .C(_08899_),
    .Y(_08900_));
 OR3x1_ASAP7_75t_R _27378_ (.A(_00682_),
    .B(_05815_),
    .C(_07061_),
    .Y(_08901_));
 OA211x2_ASAP7_75t_R _27379_ (.A1(_07868_),
    .A2(_07064_),
    .B(_08901_),
    .C(_07060_),
    .Y(_08902_));
 NOR2x1_ASAP7_75t_R _27380_ (.A(net2311),
    .B(_08665_),
    .Y(_08903_));
 OR5x1_ASAP7_75t_R _27381_ (.A(net308),
    .B(_08798_),
    .C(_08900_),
    .D(_08902_),
    .E(_08903_),
    .Y(_08904_));
 OAI21x1_ASAP7_75t_R _27382_ (.A1(_00682_),
    .A2(_08660_),
    .B(_08904_),
    .Y(_02698_));
 INVx1_ASAP7_75t_R _27383_ (.A(net152),
    .Y(_08905_));
 AND2x2_ASAP7_75t_R _27384_ (.A(_08905_),
    .B(_08748_),
    .Y(_08906_));
 AO21x1_ASAP7_75t_R _27385_ (.A1(_00684_),
    .A2(_08746_),
    .B(_08906_),
    .Y(_08907_));
 OA211x2_ASAP7_75t_R _27386_ (.A1(_01320_),
    .A2(_08874_),
    .B(_08806_),
    .C(_01335_),
    .Y(_08908_));
 AO21x1_ASAP7_75t_R _27387_ (.A1(_08744_),
    .A2(_08907_),
    .B(_08908_),
    .Y(_08909_));
 AO21x1_ASAP7_75t_R _27388_ (.A1(_08894_),
    .A2(_08895_),
    .B(_01357_),
    .Y(_08910_));
 OA211x2_ASAP7_75t_R _27389_ (.A1(_00285_),
    .A2(_08905_),
    .B(_08777_),
    .C(_08910_),
    .Y(_08911_));
 OA21x2_ASAP7_75t_R _27390_ (.A1(_01727_),
    .A2(_08909_),
    .B(_08911_),
    .Y(_08912_));
 NOR2x1_ASAP7_75t_R _27391_ (.A(_14783_),
    .B(_08665_),
    .Y(_08913_));
 OR4x1_ASAP7_75t_R _27392_ (.A(_07910_),
    .B(_08798_),
    .C(_08912_),
    .D(_08913_),
    .Y(_08914_));
 OAI21x1_ASAP7_75t_R _27393_ (.A1(_00684_),
    .A2(_08660_),
    .B(_08914_),
    .Y(_02699_));
 AO32x1_ASAP7_75t_R _27394_ (.A1(_07963_),
    .A2(_14843_),
    .A3(_07519_),
    .B1(_08858_),
    .B2(_00686_),
    .Y(_08915_));
 OA21x2_ASAP7_75t_R _27395_ (.A1(_00285_),
    .A2(_05796_),
    .B(_08651_),
    .Y(_08916_));
 OA21x2_ASAP7_75t_R _27396_ (.A1(_01357_),
    .A2(_08907_),
    .B(_08916_),
    .Y(_08917_));
 NOR2x1_ASAP7_75t_R _27397_ (.A(_14099_),
    .B(_08851_),
    .Y(_08918_));
 OR2x2_ASAP7_75t_R _27398_ (.A(_00686_),
    .B(_08748_),
    .Y(_08919_));
 NAND2x1_ASAP7_75t_R _27399_ (.A(net153),
    .B(_08748_),
    .Y(_08920_));
 AO21x1_ASAP7_75t_R _27400_ (.A1(_08919_),
    .A2(_08920_),
    .B(_08806_),
    .Y(_08921_));
 OR4x1_ASAP7_75t_R _27401_ (.A(_01321_),
    .B(_17825_),
    .C(_08746_),
    .D(_08873_),
    .Y(_08922_));
 AO21x1_ASAP7_75t_R _27402_ (.A1(_01336_),
    .A2(_08922_),
    .B(_08744_),
    .Y(_08923_));
 AO21x1_ASAP7_75t_R _27403_ (.A1(_08921_),
    .A2(_08923_),
    .B(_01727_),
    .Y(_08924_));
 OA211x2_ASAP7_75t_R _27404_ (.A1(_08917_),
    .A2(_08918_),
    .B(_08850_),
    .C(_08924_),
    .Y(_08925_));
 NOR2x1_ASAP7_75t_R _27405_ (.A(_08915_),
    .B(_08925_),
    .Y(_02700_));
 OR4x1_ASAP7_75t_R _27406_ (.A(_01322_),
    .B(_17825_),
    .C(_05774_),
    .D(_08746_),
    .Y(_08926_));
 AND2x4_ASAP7_75t_R _27407_ (.A(_13604_),
    .B(_05766_),
    .Y(_08927_));
 AND2x2_ASAP7_75t_R _27408_ (.A(_06428_),
    .B(_08748_),
    .Y(_08928_));
 AO21x1_ASAP7_75t_R _27409_ (.A1(_00718_),
    .A2(_08746_),
    .B(_08928_),
    .Y(_08929_));
 AO32x1_ASAP7_75t_R _27410_ (.A1(_01337_),
    .A2(_08926_),
    .A3(_08927_),
    .B1(_08744_),
    .B2(_08929_),
    .Y(_08930_));
 OA21x2_ASAP7_75t_R _27411_ (.A1(_00285_),
    .A2(_06428_),
    .B(_08777_),
    .Y(_08931_));
 AO21x1_ASAP7_75t_R _27412_ (.A1(_08919_),
    .A2(_08920_),
    .B(_01357_),
    .Y(_08932_));
 OA211x2_ASAP7_75t_R _27413_ (.A1(_01727_),
    .A2(_08930_),
    .B(_08931_),
    .C(_08932_),
    .Y(_08933_));
 NOR2x1_ASAP7_75t_R _27414_ (.A(_15643_),
    .B(_08665_),
    .Y(_08934_));
 AND2x2_ASAP7_75t_R _27415_ (.A(_07062_),
    .B(_07995_),
    .Y(_08935_));
 AO21x1_ASAP7_75t_R _27416_ (.A1(_00718_),
    .A2(_07064_),
    .B(_08935_),
    .Y(_08936_));
 AO21x1_ASAP7_75t_R _27417_ (.A1(_07060_),
    .A2(_08936_),
    .B(net308),
    .Y(_08937_));
 OR4x1_ASAP7_75t_R _27418_ (.A(_08798_),
    .B(_08933_),
    .C(_08934_),
    .D(_08937_),
    .Y(_08938_));
 OAI21x1_ASAP7_75t_R _27419_ (.A1(_00718_),
    .A2(_08660_),
    .B(_08938_),
    .Y(_02701_));
 OR3x1_ASAP7_75t_R _27420_ (.A(_00750_),
    .B(_05815_),
    .C(_07061_),
    .Y(_08939_));
 OA211x2_ASAP7_75t_R _27421_ (.A1(_08044_),
    .A2(_07064_),
    .B(_08939_),
    .C(_07060_),
    .Y(_08940_));
 NOR2x1_ASAP7_75t_R _27422_ (.A(_15773_),
    .B(_08665_),
    .Y(_08941_));
 OR3x4_ASAP7_75t_R _27423_ (.A(_17825_),
    .B(_08746_),
    .C(_08873_),
    .Y(_08942_));
 OA211x2_ASAP7_75t_R _27424_ (.A1(_01326_),
    .A2(_08942_),
    .B(_08927_),
    .C(_01338_),
    .Y(_08943_));
 AND2x2_ASAP7_75t_R _27425_ (.A(_15778_),
    .B(_08748_),
    .Y(_08944_));
 AO21x1_ASAP7_75t_R _27426_ (.A1(_00750_),
    .A2(_08746_),
    .B(_08944_),
    .Y(_08945_));
 AO21x1_ASAP7_75t_R _27427_ (.A1(_08744_),
    .A2(_08945_),
    .B(_01727_),
    .Y(_08946_));
 OA21x2_ASAP7_75t_R _27428_ (.A1(_00285_),
    .A2(_15778_),
    .B(_08777_),
    .Y(_08947_));
 OA21x2_ASAP7_75t_R _27429_ (.A1(_01357_),
    .A2(_08929_),
    .B(_08947_),
    .Y(_08948_));
 OA21x2_ASAP7_75t_R _27430_ (.A1(_08943_),
    .A2(_08946_),
    .B(_08948_),
    .Y(_08949_));
 OR4x1_ASAP7_75t_R _27431_ (.A(_08798_),
    .B(_08940_),
    .C(_08941_),
    .D(_08949_),
    .Y(_08950_));
 OAI21x1_ASAP7_75t_R _27432_ (.A1(_00750_),
    .A2(_08660_),
    .B(_08950_),
    .Y(_02702_));
 OA211x2_ASAP7_75t_R _27433_ (.A1(_01320_),
    .A2(_08942_),
    .B(_08806_),
    .C(_01339_),
    .Y(_08951_));
 AND2x2_ASAP7_75t_R _27434_ (.A(_00785_),
    .B(_08748_),
    .Y(_08952_));
 AO21x1_ASAP7_75t_R _27435_ (.A1(_00783_),
    .A2(_08746_),
    .B(_08952_),
    .Y(_08953_));
 AO21x1_ASAP7_75t_R _27436_ (.A1(_08744_),
    .A2(_08953_),
    .B(_01727_),
    .Y(_08954_));
 OA21x2_ASAP7_75t_R _27437_ (.A1(_00285_),
    .A2(_00785_),
    .B(_08777_),
    .Y(_08955_));
 OA21x2_ASAP7_75t_R _27438_ (.A1(_01357_),
    .A2(_08945_),
    .B(_08955_),
    .Y(_08956_));
 OAI21x1_ASAP7_75t_R _27439_ (.A1(_08951_),
    .A2(_08954_),
    .B(_08956_),
    .Y(_08957_));
 NAND2x1_ASAP7_75t_R _27440_ (.A(_07060_),
    .B(_08091_),
    .Y(_08958_));
 OA211x2_ASAP7_75t_R _27441_ (.A1(_05957_),
    .A2(_08665_),
    .B(_08958_),
    .C(_13817_),
    .Y(_08959_));
 AND3x1_ASAP7_75t_R _27442_ (.A(_08660_),
    .B(_08957_),
    .C(_08959_),
    .Y(_08960_));
 AO21x1_ASAP7_75t_R _27443_ (.A1(_06853_),
    .A2(_08798_),
    .B(_08960_),
    .Y(_02703_));
 OA21x2_ASAP7_75t_R _27444_ (.A1(_00285_),
    .A2(_05795_),
    .B(_08651_),
    .Y(_08961_));
 OAI21x1_ASAP7_75t_R _27445_ (.A1(_01357_),
    .A2(_08953_),
    .B(_08961_),
    .Y(_08962_));
 OAI21x1_ASAP7_75t_R _27446_ (.A1(_05823_),
    .A2(_08851_),
    .B(_08962_),
    .Y(_08963_));
 OR3x4_ASAP7_75t_R _27447_ (.A(_01318_),
    .B(_05771_),
    .C(_08746_),
    .Y(_08964_));
 OA211x2_ASAP7_75t_R _27448_ (.A1(_01321_),
    .A2(_08964_),
    .B(_08927_),
    .C(_01340_),
    .Y(_08965_));
 AND2x2_ASAP7_75t_R _27449_ (.A(_05795_),
    .B(_08748_),
    .Y(_08966_));
 AO21x1_ASAP7_75t_R _27450_ (.A1(_00816_),
    .A2(_08746_),
    .B(_08966_),
    .Y(_08967_));
 AO21x1_ASAP7_75t_R _27451_ (.A1(_08744_),
    .A2(_08967_),
    .B(_01727_),
    .Y(_08968_));
 OA21x2_ASAP7_75t_R _27452_ (.A1(_08965_),
    .A2(_08968_),
    .B(_05766_),
    .Y(_08969_));
 AOI221x1_ASAP7_75t_R _27453_ (.A1(_07060_),
    .A2(_08127_),
    .B1(_08963_),
    .B2(_08969_),
    .C(net308),
    .Y(_08970_));
 NOR2x1_ASAP7_75t_R _27454_ (.A(_00816_),
    .B(_08660_),
    .Y(_08971_));
 AO21x1_ASAP7_75t_R _27455_ (.A1(_08660_),
    .A2(_08970_),
    .B(_08971_),
    .Y(_02704_));
 OR4x2_ASAP7_75t_R _27456_ (.A(_01319_),
    .B(_01318_),
    .C(_05771_),
    .D(_08746_),
    .Y(_08972_));
 NOR2x1_ASAP7_75t_R _27457_ (.A(net2255),
    .B(_08746_),
    .Y(_08973_));
 AO21x1_ASAP7_75t_R _27458_ (.A1(_00849_),
    .A2(_08746_),
    .B(_08973_),
    .Y(_08974_));
 AO32x1_ASAP7_75t_R _27459_ (.A1(_01341_),
    .A2(_08664_),
    .A3(_08972_),
    .B1(_08974_),
    .B2(_08744_),
    .Y(_08975_));
 NAND2x1_ASAP7_75t_R _27460_ (.A(_13775_),
    .B(net2256),
    .Y(_08976_));
 OA211x2_ASAP7_75t_R _27461_ (.A1(_01357_),
    .A2(_08967_),
    .B(_08976_),
    .C(_08777_),
    .Y(_08977_));
 OA21x2_ASAP7_75t_R _27462_ (.A1(_01727_),
    .A2(_08975_),
    .B(_08977_),
    .Y(_08978_));
 NOR2x1_ASAP7_75t_R _27463_ (.A(_16138_),
    .B(_08665_),
    .Y(_08979_));
 OR4x1_ASAP7_75t_R _27464_ (.A(_08184_),
    .B(_08798_),
    .C(_08978_),
    .D(_08979_),
    .Y(_08980_));
 OAI21x1_ASAP7_75t_R _27465_ (.A1(_00849_),
    .A2(_08660_),
    .B(_08980_),
    .Y(_02705_));
 OA21x2_ASAP7_75t_R _27466_ (.A1(_01326_),
    .A2(_08964_),
    .B(_01342_),
    .Y(_08981_));
 AND2x2_ASAP7_75t_R _27467_ (.A(_16263_),
    .B(_08748_),
    .Y(_08982_));
 AO21x1_ASAP7_75t_R _27468_ (.A1(_00881_),
    .A2(_08746_),
    .B(_08982_),
    .Y(_08983_));
 AO21x1_ASAP7_75t_R _27469_ (.A1(_08744_),
    .A2(_08983_),
    .B(_01727_),
    .Y(_08984_));
 AO21x1_ASAP7_75t_R _27470_ (.A1(_08806_),
    .A2(_08981_),
    .B(_08984_),
    .Y(_08985_));
 OA21x2_ASAP7_75t_R _27471_ (.A1(_00285_),
    .A2(_16263_),
    .B(_08777_),
    .Y(_08986_));
 OA21x2_ASAP7_75t_R _27472_ (.A1(_01357_),
    .A2(_08974_),
    .B(_08986_),
    .Y(_08987_));
 AO221x1_ASAP7_75t_R _27473_ (.A1(_16261_),
    .A2(_08867_),
    .B1(_08985_),
    .B2(_08987_),
    .C(_08209_),
    .Y(_08988_));
 AND2x2_ASAP7_75t_R _27474_ (.A(_00881_),
    .B(_08798_),
    .Y(_08989_));
 AOI21x1_ASAP7_75t_R _27475_ (.A1(_08660_),
    .A2(_08988_),
    .B(_08989_),
    .Y(_02706_));
 INVx1_ASAP7_75t_R _27476_ (.A(_00914_),
    .Y(_08990_));
 OA211x2_ASAP7_75t_R _27477_ (.A1(_01320_),
    .A2(_08964_),
    .B(_08664_),
    .C(_01343_),
    .Y(_08991_));
 AND2x2_ASAP7_75t_R _27478_ (.A(_06472_),
    .B(_08748_),
    .Y(_08992_));
 AO21x1_ASAP7_75t_R _27479_ (.A1(_00914_),
    .A2(_08746_),
    .B(_08992_),
    .Y(_08993_));
 AO21x1_ASAP7_75t_R _27480_ (.A1(_08744_),
    .A2(_08993_),
    .B(_01727_),
    .Y(_08994_));
 OA21x2_ASAP7_75t_R _27481_ (.A1(_00285_),
    .A2(_06472_),
    .B(_08777_),
    .Y(_08995_));
 OA21x2_ASAP7_75t_R _27482_ (.A1(_01357_),
    .A2(_08983_),
    .B(_08995_),
    .Y(_08996_));
 OAI21x1_ASAP7_75t_R _27483_ (.A1(_08991_),
    .A2(_08994_),
    .B(_08996_),
    .Y(_08997_));
 OA211x2_ASAP7_75t_R _27484_ (.A1(_16378_),
    .A2(_08665_),
    .B(_08660_),
    .C(_08241_),
    .Y(_08998_));
 AO22x1_ASAP7_75t_R _27485_ (.A1(_08990_),
    .A2(_08798_),
    .B1(_08997_),
    .B2(_08998_),
    .Y(_02707_));
 OAI22x1_ASAP7_75t_R _27486_ (.A1(_00285_),
    .A2(_16509_),
    .B1(_08993_),
    .B2(_01357_),
    .Y(_08999_));
 OA22x2_ASAP7_75t_R _27487_ (.A1(_05861_),
    .A2(_08851_),
    .B1(_08999_),
    .B2(_08668_),
    .Y(_09000_));
 NAND2x2_ASAP7_75t_R _27488_ (.A(_05773_),
    .B(_01322_),
    .Y(_09001_));
 OR4x1_ASAP7_75t_R _27489_ (.A(_01321_),
    .B(_17825_),
    .C(_08746_),
    .D(_09001_),
    .Y(_09002_));
 AND3x1_ASAP7_75t_R _27490_ (.A(_01344_),
    .B(_08806_),
    .C(_09002_),
    .Y(_09003_));
 NAND2x1_ASAP7_75t_R _27491_ (.A(_16509_),
    .B(_08748_),
    .Y(_09004_));
 NAND2x1_ASAP7_75t_R _27492_ (.A(_00946_),
    .B(_08746_),
    .Y(_09005_));
 AOI21x1_ASAP7_75t_R _27493_ (.A1(_09004_),
    .A2(_09005_),
    .B(_08806_),
    .Y(_09006_));
 OR3x1_ASAP7_75t_R _27494_ (.A(_01727_),
    .B(_09003_),
    .C(_09006_),
    .Y(_09007_));
 NAND2x1_ASAP7_75t_R _27495_ (.A(_08850_),
    .B(_09007_),
    .Y(_09008_));
 NOR2x1_ASAP7_75t_R _27496_ (.A(_00946_),
    .B(_08660_),
    .Y(_09009_));
 AO21x1_ASAP7_75t_R _27497_ (.A1(_08271_),
    .A2(_08660_),
    .B(_09009_),
    .Y(_09010_));
 OA21x2_ASAP7_75t_R _27498_ (.A1(_09000_),
    .A2(_09008_),
    .B(_09010_),
    .Y(_02708_));
 NAND2x1_ASAP7_75t_R _27499_ (.A(_08305_),
    .B(_08660_),
    .Y(_09011_));
 OA21x2_ASAP7_75t_R _27500_ (.A1(_00979_),
    .A2(_08660_),
    .B(_09011_),
    .Y(_09012_));
 OR3x2_ASAP7_75t_R _27501_ (.A(_01319_),
    .B(_01318_),
    .C(_08821_),
    .Y(_09013_));
 AND3x1_ASAP7_75t_R _27502_ (.A(_01345_),
    .B(_08664_),
    .C(_09013_),
    .Y(_09014_));
 NOR2x1_ASAP7_75t_R _27503_ (.A(net162),
    .B(_08746_),
    .Y(_09015_));
 AO21x1_ASAP7_75t_R _27504_ (.A1(_00979_),
    .A2(_08746_),
    .B(_09015_),
    .Y(_09016_));
 AO21x1_ASAP7_75t_R _27505_ (.A1(_08744_),
    .A2(_09016_),
    .B(_01727_),
    .Y(_09017_));
 AND3x1_ASAP7_75t_R _27506_ (.A(_05765_),
    .B(_09004_),
    .C(_09005_),
    .Y(_09018_));
 AO21x1_ASAP7_75t_R _27507_ (.A1(_13775_),
    .A2(net162),
    .B(_08668_),
    .Y(_09019_));
 OAI22x1_ASAP7_75t_R _27508_ (.A1(_16617_),
    .A2(_08851_),
    .B1(_09018_),
    .B2(_09019_),
    .Y(_09020_));
 OA211x2_ASAP7_75t_R _27509_ (.A1(_09014_),
    .A2(_09017_),
    .B(_09020_),
    .C(_08850_),
    .Y(_09021_));
 NOR2x1_ASAP7_75t_R _27510_ (.A(_09012_),
    .B(_09021_),
    .Y(_02709_));
 OR3x4_ASAP7_75t_R _27511_ (.A(_17825_),
    .B(_08746_),
    .C(_09001_),
    .Y(_09022_));
 OA211x2_ASAP7_75t_R _27512_ (.A1(_01326_),
    .A2(_09022_),
    .B(_08927_),
    .C(_01346_),
    .Y(_09023_));
 AND2x2_ASAP7_75t_R _27513_ (.A(_04517_),
    .B(_08748_),
    .Y(_09024_));
 AO21x1_ASAP7_75t_R _27514_ (.A1(_01011_),
    .A2(_08746_),
    .B(_09024_),
    .Y(_09025_));
 AO21x1_ASAP7_75t_R _27515_ (.A1(_08744_),
    .A2(_09025_),
    .B(_01727_),
    .Y(_09026_));
 OAI22x1_ASAP7_75t_R _27516_ (.A1(_00285_),
    .A2(_04517_),
    .B1(_09016_),
    .B2(_01357_),
    .Y(_09027_));
 OAI22x1_ASAP7_75t_R _27517_ (.A1(_05877_),
    .A2(_08851_),
    .B1(_09027_),
    .B2(_08668_),
    .Y(_09028_));
 OA211x2_ASAP7_75t_R _27518_ (.A1(_09023_),
    .A2(_09026_),
    .B(_09028_),
    .C(_05766_),
    .Y(_09029_));
 AOI211x1_ASAP7_75t_R _27519_ (.A1(_07060_),
    .A2(_08345_),
    .B(_08798_),
    .C(net308),
    .Y(_09030_));
 INVx1_ASAP7_75t_R _27520_ (.A(_09030_),
    .Y(_09031_));
 OAI22x1_ASAP7_75t_R _27521_ (.A1(_01011_),
    .A2(_08660_),
    .B1(_09029_),
    .B2(_09031_),
    .Y(_02710_));
 INVx1_ASAP7_75t_R _27522_ (.A(_01045_),
    .Y(_09032_));
 OA211x2_ASAP7_75t_R _27523_ (.A1(_01320_),
    .A2(_09022_),
    .B(_08927_),
    .C(_01347_),
    .Y(_09033_));
 AND2x2_ASAP7_75t_R _27524_ (.A(_06498_),
    .B(_08748_),
    .Y(_09034_));
 AO21x1_ASAP7_75t_R _27525_ (.A1(_01045_),
    .A2(_08746_),
    .B(_09034_),
    .Y(_09035_));
 AO21x1_ASAP7_75t_R _27526_ (.A1(_08744_),
    .A2(_09035_),
    .B(_01727_),
    .Y(_09036_));
 OA21x2_ASAP7_75t_R _27527_ (.A1(_00285_),
    .A2(_06498_),
    .B(_08777_),
    .Y(_09037_));
 OA21x2_ASAP7_75t_R _27528_ (.A1(_01357_),
    .A2(_09025_),
    .B(_09037_),
    .Y(_09038_));
 OAI21x1_ASAP7_75t_R _27529_ (.A1(_09033_),
    .A2(_09036_),
    .B(_09038_),
    .Y(_09039_));
 OA211x2_ASAP7_75t_R _27530_ (.A1(_04624_),
    .A2(_08665_),
    .B(_08371_),
    .C(_13817_),
    .Y(_09040_));
 AND3x1_ASAP7_75t_R _27531_ (.A(_08660_),
    .B(_09039_),
    .C(_09040_),
    .Y(_09041_));
 AO21x1_ASAP7_75t_R _27532_ (.A1(_09032_),
    .A2(_08798_),
    .B(_09041_),
    .Y(_02711_));
 OAI21x1_ASAP7_75t_R _27533_ (.A1(_05892_),
    .A2(_08665_),
    .B(_08660_),
    .Y(_09042_));
 OA21x2_ASAP7_75t_R _27534_ (.A1(_01077_),
    .A2(_08660_),
    .B(_09042_),
    .Y(_09043_));
 OA211x2_ASAP7_75t_R _27535_ (.A1(_00285_),
    .A2(_04747_),
    .B(_08651_),
    .C(_08850_),
    .Y(_09044_));
 OR3x4_ASAP7_75t_R _27536_ (.A(_01318_),
    .B(_01322_),
    .C(_08884_),
    .Y(_09045_));
 OA211x2_ASAP7_75t_R _27537_ (.A1(_01321_),
    .A2(_09045_),
    .B(_08664_),
    .C(_01348_),
    .Y(_09046_));
 OR2x2_ASAP7_75t_R _27538_ (.A(_01077_),
    .B(_08748_),
    .Y(_09047_));
 NAND2x1_ASAP7_75t_R _27539_ (.A(net165),
    .B(_08748_),
    .Y(_09048_));
 AND3x1_ASAP7_75t_R _27540_ (.A(_08744_),
    .B(_09047_),
    .C(_09048_),
    .Y(_09049_));
 OR3x1_ASAP7_75t_R _27541_ (.A(_01727_),
    .B(_09046_),
    .C(_09049_),
    .Y(_09050_));
 OA211x2_ASAP7_75t_R _27542_ (.A1(_01357_),
    .A2(_09035_),
    .B(_09044_),
    .C(_09050_),
    .Y(_09051_));
 AOI211x1_ASAP7_75t_R _27543_ (.A1(_14843_),
    .A2(_08416_),
    .B(_09043_),
    .C(_09051_),
    .Y(_02712_));
 AND2x2_ASAP7_75t_R _27544_ (.A(_06511_),
    .B(_08748_),
    .Y(_09052_));
 AO21x1_ASAP7_75t_R _27545_ (.A1(_01110_),
    .A2(_08746_),
    .B(_09052_),
    .Y(_09053_));
 OR3x2_ASAP7_75t_R _27546_ (.A(_01319_),
    .B(_01318_),
    .C(_01322_),
    .Y(_09054_));
 OA211x2_ASAP7_75t_R _27547_ (.A1(_08884_),
    .A2(_09054_),
    .B(_01349_),
    .C(_08806_),
    .Y(_09055_));
 AO21x1_ASAP7_75t_R _27548_ (.A1(_08744_),
    .A2(_09053_),
    .B(_09055_),
    .Y(_09056_));
 AO21x1_ASAP7_75t_R _27549_ (.A1(_09047_),
    .A2(_09048_),
    .B(_01357_),
    .Y(_09057_));
 OA211x2_ASAP7_75t_R _27550_ (.A1(_00285_),
    .A2(_06511_),
    .B(_08777_),
    .C(_09057_),
    .Y(_09058_));
 OAI21x1_ASAP7_75t_R _27551_ (.A1(_01727_),
    .A2(_09056_),
    .B(_09058_),
    .Y(_09059_));
 OA211x2_ASAP7_75t_R _27552_ (.A1(_04854_),
    .A2(_08665_),
    .B(_09059_),
    .C(_08464_),
    .Y(_09060_));
 NOR2x1_ASAP7_75t_R _27553_ (.A(_01110_),
    .B(_08660_),
    .Y(_09061_));
 AO21x1_ASAP7_75t_R _27554_ (.A1(_08660_),
    .A2(_09060_),
    .B(_09061_),
    .Y(_02713_));
 OA211x2_ASAP7_75t_R _27555_ (.A1(_01326_),
    .A2(_09045_),
    .B(_08806_),
    .C(_01350_),
    .Y(_09062_));
 AND2x2_ASAP7_75t_R _27556_ (.A(_04968_),
    .B(_08748_),
    .Y(_09063_));
 AO21x1_ASAP7_75t_R _27557_ (.A1(_01142_),
    .A2(_08746_),
    .B(_09063_),
    .Y(_09064_));
 AO21x1_ASAP7_75t_R _27558_ (.A1(_08744_),
    .A2(_09064_),
    .B(_01727_),
    .Y(_09065_));
 OA21x2_ASAP7_75t_R _27559_ (.A1(_00285_),
    .A2(_04968_),
    .B(_08777_),
    .Y(_09066_));
 OA21x2_ASAP7_75t_R _27560_ (.A1(_01357_),
    .A2(_09053_),
    .B(_09066_),
    .Y(_09067_));
 OA21x2_ASAP7_75t_R _27561_ (.A1(_09062_),
    .A2(_09065_),
    .B(_09067_),
    .Y(_09068_));
 NOR2x1_ASAP7_75t_R _27562_ (.A(_04965_),
    .B(_08665_),
    .Y(_09069_));
 OR4x1_ASAP7_75t_R _27563_ (.A(_08490_),
    .B(_08798_),
    .C(_09068_),
    .D(_09069_),
    .Y(_09070_));
 OAI21x1_ASAP7_75t_R _27564_ (.A1(_01142_),
    .A2(_08660_),
    .B(_09070_),
    .Y(_02714_));
 OA211x2_ASAP7_75t_R _27565_ (.A1(_01320_),
    .A2(_09045_),
    .B(_08664_),
    .C(_01351_),
    .Y(_09071_));
 AND2x2_ASAP7_75t_R _27566_ (.A(_06526_),
    .B(_08748_),
    .Y(_09072_));
 AO21x1_ASAP7_75t_R _27567_ (.A1(_01176_),
    .A2(_08746_),
    .B(_09072_),
    .Y(_09073_));
 AO21x1_ASAP7_75t_R _27568_ (.A1(_08744_),
    .A2(_09073_),
    .B(_01727_),
    .Y(_09074_));
 OA21x2_ASAP7_75t_R _27569_ (.A1(_00285_),
    .A2(_06526_),
    .B(_08777_),
    .Y(_09075_));
 OA21x2_ASAP7_75t_R _27570_ (.A1(_01357_),
    .A2(_09064_),
    .B(_09075_),
    .Y(_09076_));
 OA21x2_ASAP7_75t_R _27571_ (.A1(_09071_),
    .A2(_09074_),
    .B(_09076_),
    .Y(_09077_));
 NOR2x1_ASAP7_75t_R _27572_ (.A(_05075_),
    .B(_08665_),
    .Y(_09078_));
 AO21x1_ASAP7_75t_R _27573_ (.A1(_07060_),
    .A2(_08516_),
    .B(_09078_),
    .Y(_09079_));
 OR3x1_ASAP7_75t_R _27574_ (.A(_08798_),
    .B(_09077_),
    .C(_09079_),
    .Y(_09080_));
 OAI21x1_ASAP7_75t_R _27575_ (.A1(_01176_),
    .A2(_08660_),
    .B(_09080_),
    .Y(_02715_));
 AND2x2_ASAP7_75t_R _27576_ (.A(_05185_),
    .B(_08748_),
    .Y(_09081_));
 AO21x1_ASAP7_75t_R _27577_ (.A1(_01208_),
    .A2(_08746_),
    .B(_09081_),
    .Y(_09082_));
 OR4x2_ASAP7_75t_R _27578_ (.A(_01318_),
    .B(_01322_),
    .C(_17825_),
    .D(_08746_),
    .Y(_09083_));
 OA211x2_ASAP7_75t_R _27579_ (.A1(_01321_),
    .A2(_09083_),
    .B(_08806_),
    .C(_01352_),
    .Y(_09084_));
 AO21x1_ASAP7_75t_R _27580_ (.A1(_08744_),
    .A2(_09082_),
    .B(_09084_),
    .Y(_09085_));
 OA21x2_ASAP7_75t_R _27581_ (.A1(_00285_),
    .A2(_05185_),
    .B(_08651_),
    .Y(_09086_));
 OAI21x1_ASAP7_75t_R _27582_ (.A1(_01357_),
    .A2(_09073_),
    .B(_09086_),
    .Y(_09087_));
 OAI21x1_ASAP7_75t_R _27583_ (.A1(_05924_),
    .A2(_08851_),
    .B(_09087_),
    .Y(_09088_));
 OA211x2_ASAP7_75t_R _27584_ (.A1(_01727_),
    .A2(_09085_),
    .B(_09088_),
    .C(_08850_),
    .Y(_09089_));
 AOI221x1_ASAP7_75t_R _27585_ (.A1(_14843_),
    .A2(_08540_),
    .B1(_08798_),
    .B2(_01208_),
    .C(_09089_),
    .Y(_02716_));
 NOR2x1_ASAP7_75t_R _27586_ (.A(_01357_),
    .B(_09082_),
    .Y(_09090_));
 AO21x1_ASAP7_75t_R _27587_ (.A1(_13775_),
    .A2(net2137),
    .B(_08668_),
    .Y(_09091_));
 OAI22x1_ASAP7_75t_R _27588_ (.A1(_05936_),
    .A2(_08851_),
    .B1(_09090_),
    .B2(_09091_),
    .Y(_09092_));
 OR3x1_ASAP7_75t_R _27589_ (.A(_17825_),
    .B(_08746_),
    .C(_09054_),
    .Y(_09093_));
 AND2x2_ASAP7_75t_R _27590_ (.A(_06541_),
    .B(_08748_),
    .Y(_09094_));
 AO21x1_ASAP7_75t_R _27591_ (.A1(_01242_),
    .A2(_08746_),
    .B(_09094_),
    .Y(_09095_));
 AO32x1_ASAP7_75t_R _27592_ (.A1(_01353_),
    .A2(_08664_),
    .A3(_09093_),
    .B1(_09095_),
    .B2(_08744_),
    .Y(_09096_));
 OA21x2_ASAP7_75t_R _27593_ (.A1(_01727_),
    .A2(_09096_),
    .B(_05766_),
    .Y(_09097_));
 AOI221x1_ASAP7_75t_R _27594_ (.A1(_07060_),
    .A2(_08574_),
    .B1(_09092_),
    .B2(_09097_),
    .C(net308),
    .Y(_09098_));
 NOR2x1_ASAP7_75t_R _27595_ (.A(_01242_),
    .B(_08660_),
    .Y(_09099_));
 AO21x1_ASAP7_75t_R _27596_ (.A1(_08660_),
    .A2(_09098_),
    .B(_09099_),
    .Y(_02717_));
 OA211x2_ASAP7_75t_R _27597_ (.A1(_01326_),
    .A2(_09083_),
    .B(_08927_),
    .C(_01354_),
    .Y(_09100_));
 AND2x2_ASAP7_75t_R _27598_ (.A(_05404_),
    .B(_08748_),
    .Y(_09101_));
 AO21x1_ASAP7_75t_R _27599_ (.A1(_01274_),
    .A2(_08746_),
    .B(_09101_),
    .Y(_09102_));
 AO21x1_ASAP7_75t_R _27600_ (.A1(_08744_),
    .A2(_09102_),
    .B(_01727_),
    .Y(_09103_));
 OAI22x1_ASAP7_75t_R _27601_ (.A1(_00285_),
    .A2(_05404_),
    .B1(_09095_),
    .B2(_01357_),
    .Y(_09104_));
 OAI22x1_ASAP7_75t_R _27602_ (.A1(_05400_),
    .A2(_08851_),
    .B1(_09104_),
    .B2(_08668_),
    .Y(_09105_));
 OA211x2_ASAP7_75t_R _27603_ (.A1(_09100_),
    .A2(_09103_),
    .B(_09105_),
    .C(_08850_),
    .Y(_09106_));
 AOI221x1_ASAP7_75t_R _27604_ (.A1(_14843_),
    .A2(_08613_),
    .B1(_08798_),
    .B2(_01274_),
    .C(_09106_),
    .Y(_02718_));
 OA211x2_ASAP7_75t_R _27605_ (.A1(_01320_),
    .A2(_09083_),
    .B(_08664_),
    .C(_01355_),
    .Y(_09107_));
 OR3x1_ASAP7_75t_R _27606_ (.A(_01308_),
    .B(_05540_),
    .C(_05541_),
    .Y(_09108_));
 AO21x1_ASAP7_75t_R _27607_ (.A1(_08744_),
    .A2(_09108_),
    .B(_01727_),
    .Y(_09109_));
 OA21x2_ASAP7_75t_R _27608_ (.A1(_00285_),
    .A2(_05542_),
    .B(_08651_),
    .Y(_09110_));
 OA21x2_ASAP7_75t_R _27609_ (.A1(_01357_),
    .A2(_09102_),
    .B(_09110_),
    .Y(_09111_));
 OAI21x1_ASAP7_75t_R _27610_ (.A1(_09107_),
    .A2(_09109_),
    .B(_09111_),
    .Y(_09112_));
 TAPCELL_ASAP7_75t_R PHY_643 ();
 OA21x2_ASAP7_75t_R _27612_ (.A1(_05513_),
    .A2(_08851_),
    .B(_08850_),
    .Y(_09114_));
 AND2x2_ASAP7_75t_R _27613_ (.A(_08636_),
    .B(_08660_),
    .Y(_09115_));
 AO221x1_ASAP7_75t_R _27614_ (.A1(_05536_),
    .A2(_08798_),
    .B1(_09112_),
    .B2(_09114_),
    .C(_09115_),
    .Y(_02719_));
 OA33x2_ASAP7_75t_R _27615_ (.A1(_01308_),
    .A2(_01357_),
    .A3(_05542_),
    .B1(_05547_),
    .B2(_08651_),
    .B3(_08653_),
    .Y(_09116_));
 AND3x1_ASAP7_75t_R _27616_ (.A(_02261_),
    .B(_07060_),
    .C(_07062_),
    .Y(_09117_));
 INVx1_ASAP7_75t_R _27617_ (.A(_09117_),
    .Y(_09118_));
 OA211x2_ASAP7_75t_R _27618_ (.A1(_07060_),
    .A2(_09116_),
    .B(_09118_),
    .C(_08660_),
    .Y(_09119_));
 AOI21x1_ASAP7_75t_R _27619_ (.A1(_01677_),
    .A2(_08798_),
    .B(_09119_),
    .Y(_02720_));
 INVx1_ASAP7_75t_R _27620_ (.A(_00034_),
    .Y(_09120_));
 XNOR2x1_ASAP7_75t_R _27621_ (.B(_02256_),
    .Y(_09121_),
    .A(_00070_));
 XNOR2x1_ASAP7_75t_R _27622_ (.B(_17744_),
    .Y(_09122_),
    .A(_00069_));
 XNOR2x1_ASAP7_75t_R _27623_ (.B(_09122_),
    .Y(_09123_),
    .A(_09121_));
 XNOR2x1_ASAP7_75t_R _27624_ (.B(_17720_),
    .Y(_09124_),
    .A(_00068_));
 XNOR2x1_ASAP7_75t_R _27625_ (.B(_09124_),
    .Y(_09125_),
    .A(_09123_));
 XOR2x1_ASAP7_75t_R _27626_ (.A(net2125),
    .Y(_09126_),
    .B(net2159));
 XNOR2x1_ASAP7_75t_R _27627_ (.B(_00071_),
    .Y(_09127_),
    .A(_17689_));
 XNOR2x1_ASAP7_75t_R _27628_ (.B(_09127_),
    .Y(_09128_),
    .A(_09126_));
 XNOR2x1_ASAP7_75t_R _27629_ (.B(_02260_),
    .Y(_09129_),
    .A(_02259_));
 XNOR2x1_ASAP7_75t_R _27630_ (.B(_02258_),
    .Y(_09130_),
    .A(_02257_));
 XNOR2x1_ASAP7_75t_R _27631_ (.B(_09130_),
    .Y(_09131_),
    .A(_09129_));
 XNOR2x1_ASAP7_75t_R _27632_ (.B(_09131_),
    .Y(_09132_),
    .A(_09128_));
 XNOR2x1_ASAP7_75t_R _27633_ (.B(_09132_),
    .Y(_09133_),
    .A(_09125_));
 OA21x2_ASAP7_75t_R _27634_ (.A1(_00034_),
    .A2(_05548_),
    .B(_05967_),
    .Y(_09134_));
 XNOR2x1_ASAP7_75t_R _27635_ (.B(_09134_),
    .Y(_09135_),
    .A(_09133_));
 NAND2x1_ASAP7_75t_R _27636_ (.A(_17712_),
    .B(_17736_),
    .Y(_09136_));
 XNOR2x1_ASAP7_75t_R _27637_ (.B(_09136_),
    .Y(_09137_),
    .A(_09135_));
 AO221x1_ASAP7_75t_R _27638_ (.A1(_08668_),
    .A2(_08664_),
    .B1(_09137_),
    .B2(_07519_),
    .C(_08798_),
    .Y(_09138_));
 OA21x2_ASAP7_75t_R _27639_ (.A1(_09120_),
    .A2(_08660_),
    .B(_09138_),
    .Y(_02721_));
 NAND2x2_ASAP7_75t_R _27640_ (.A(_05781_),
    .B(_05777_),
    .Y(_09139_));
 TAPCELL_ASAP7_75t_R PHY_642 ();
 TAPCELL_ASAP7_75t_R PHY_641 ();
 AND2x6_ASAP7_75t_R _27643_ (.A(_05781_),
    .B(_05777_),
    .Y(_09142_));
 TAPCELL_ASAP7_75t_R PHY_640 ();
 TAPCELL_ASAP7_75t_R PHY_639 ();
 NAND2x1_ASAP7_75t_R _27646_ (.A(_13981_),
    .B(_08655_),
    .Y(_09145_));
 OA211x2_ASAP7_75t_R _27647_ (.A1(_16721_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09145_),
    .Y(_09146_));
 AOI21x1_ASAP7_75t_R _27648_ (.A1(_01676_),
    .A2(_09139_),
    .B(_09146_),
    .Y(_02722_));
 TAPCELL_ASAP7_75t_R PHY_638 ();
 NAND2x1_ASAP7_75t_R _27650_ (.A(_13767_),
    .B(_08655_),
    .Y(_09148_));
 OA211x2_ASAP7_75t_R _27651_ (.A1(_16717_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09148_),
    .Y(_09149_));
 AOI21x1_ASAP7_75t_R _27652_ (.A1(_01675_),
    .A2(_09139_),
    .B(_09149_),
    .Y(_02723_));
 NAND2x1_ASAP7_75t_R _27653_ (.A(_14921_),
    .B(_08655_),
    .Y(_09150_));
 OA211x2_ASAP7_75t_R _27654_ (.A1(_05792_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09150_),
    .Y(_09151_));
 AOI21x1_ASAP7_75t_R _27655_ (.A1(_01674_),
    .A2(_09139_),
    .B(_09151_),
    .Y(_02724_));
 TAPCELL_ASAP7_75t_R PHY_637 ();
 TAPCELL_ASAP7_75t_R PHY_636 ();
 TAPCELL_ASAP7_75t_R PHY_635 ();
 TAPCELL_ASAP7_75t_R PHY_634 ();
 AO21x1_ASAP7_75t_R _27660_ (.A1(_05513_),
    .A2(_05950_),
    .B(_14980_),
    .Y(_09156_));
 OA211x2_ASAP7_75t_R _27661_ (.A1(net293),
    .A2(_08655_),
    .B(_09142_),
    .C(_09156_),
    .Y(_09157_));
 AO21x1_ASAP7_75t_R _27662_ (.A1(_08675_),
    .A2(_09139_),
    .B(_09157_),
    .Y(_02725_));
 NAND2x1_ASAP7_75t_R _27663_ (.A(net2323),
    .B(_08655_),
    .Y(_09158_));
 OA211x2_ASAP7_75t_R _27664_ (.A1(_05791_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09158_),
    .Y(_09159_));
 AOI21x1_ASAP7_75t_R _27665_ (.A1(_01672_),
    .A2(_09139_),
    .B(_09159_),
    .Y(_02726_));
 AO21x1_ASAP7_75t_R _27666_ (.A1(_05513_),
    .A2(_05950_),
    .B(_15103_),
    .Y(_09160_));
 OA211x2_ASAP7_75t_R _27667_ (.A1(net289),
    .A2(_08655_),
    .B(_09142_),
    .C(_09160_),
    .Y(_09161_));
 AO21x1_ASAP7_75t_R _27668_ (.A1(_08696_),
    .A2(_09139_),
    .B(_09161_),
    .Y(_02727_));
 NAND2x1_ASAP7_75t_R _27669_ (.A(_15167_),
    .B(_08655_),
    .Y(_09162_));
 OA211x2_ASAP7_75t_R _27670_ (.A1(_05793_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09162_),
    .Y(_09163_));
 AOI21x1_ASAP7_75t_R _27671_ (.A1(_01670_),
    .A2(_09139_),
    .B(_09163_),
    .Y(_02728_));
 OR2x2_ASAP7_75t_R _27672_ (.A(_05885_),
    .B(_08652_),
    .Y(_09164_));
 OA211x2_ASAP7_75t_R _27673_ (.A1(_00676_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09164_),
    .Y(_09165_));
 AOI21x1_ASAP7_75t_R _27674_ (.A1(_01669_),
    .A2(_09139_),
    .B(_09165_),
    .Y(_02729_));
 AO21x1_ASAP7_75t_R _27675_ (.A1(_05513_),
    .A2(_05950_),
    .B(_15279_),
    .Y(_09166_));
 OA211x2_ASAP7_75t_R _27676_ (.A1(net179),
    .A2(_08655_),
    .B(_09142_),
    .C(_09166_),
    .Y(_09167_));
 AO21x1_ASAP7_75t_R _27677_ (.A1(_08684_),
    .A2(_09139_),
    .B(_09167_),
    .Y(_02730_));
 AO21x1_ASAP7_75t_R _27678_ (.A1(_05513_),
    .A2(_05950_),
    .B(_15331_),
    .Y(_09168_));
 OA211x2_ASAP7_75t_R _27679_ (.A1(net2204),
    .A2(_08655_),
    .B(_09142_),
    .C(_09168_),
    .Y(_09169_));
 AO21x1_ASAP7_75t_R _27680_ (.A1(_08687_),
    .A2(_09139_),
    .B(_09169_),
    .Y(_02731_));
 NAND2x1_ASAP7_75t_R _27681_ (.A(net2312),
    .B(_08655_),
    .Y(_09170_));
 OA211x2_ASAP7_75t_R _27682_ (.A1(_05797_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09170_),
    .Y(_09171_));
 AOI21x1_ASAP7_75t_R _27683_ (.A1(_01666_),
    .A2(_09139_),
    .B(_09171_),
    .Y(_02732_));
 INVx1_ASAP7_75t_R _27684_ (.A(_01665_),
    .Y(_09172_));
 TAPCELL_ASAP7_75t_R PHY_633 ();
 AO21x1_ASAP7_75t_R _27686_ (.A1(_05513_),
    .A2(_05950_),
    .B(_14783_),
    .Y(_09174_));
 OA211x2_ASAP7_75t_R _27687_ (.A1(net262),
    .A2(_08655_),
    .B(_09142_),
    .C(_09174_),
    .Y(_09175_));
 AO21x1_ASAP7_75t_R _27688_ (.A1(_09172_),
    .A2(_09139_),
    .B(_09175_),
    .Y(_02733_));
 NAND2x1_ASAP7_75t_R _27689_ (.A(_14099_),
    .B(_08655_),
    .Y(_09176_));
 OA211x2_ASAP7_75t_R _27690_ (.A1(_05796_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09176_),
    .Y(_09177_));
 AOI21x1_ASAP7_75t_R _27691_ (.A1(_01664_),
    .A2(_09139_),
    .B(_09177_),
    .Y(_02734_));
 TAPCELL_ASAP7_75t_R PHY_632 ();
 AO21x1_ASAP7_75t_R _27693_ (.A1(_05513_),
    .A2(_05950_),
    .B(_15643_),
    .Y(_09179_));
 OA211x2_ASAP7_75t_R _27694_ (.A1(net154),
    .A2(_08655_),
    .B(_09142_),
    .C(_09179_),
    .Y(_09180_));
 AO21x1_ASAP7_75t_R _27695_ (.A1(_08703_),
    .A2(_09139_),
    .B(_09180_),
    .Y(_02735_));
 NAND2x1_ASAP7_75t_R _27696_ (.A(_15773_),
    .B(_08655_),
    .Y(_09181_));
 OA211x2_ASAP7_75t_R _27697_ (.A1(_15778_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09181_),
    .Y(_09182_));
 AOI21x1_ASAP7_75t_R _27698_ (.A1(_01662_),
    .A2(_09139_),
    .B(_09182_),
    .Y(_02736_));
 INVx1_ASAP7_75t_R _27699_ (.A(_01661_),
    .Y(_09183_));
 AO21x1_ASAP7_75t_R _27700_ (.A1(_05513_),
    .A2(_05950_),
    .B(_05957_),
    .Y(_09184_));
 OA211x2_ASAP7_75t_R _27701_ (.A1(net156),
    .A2(_08655_),
    .B(_09142_),
    .C(_09184_),
    .Y(_09185_));
 AO21x1_ASAP7_75t_R _27702_ (.A1(_09183_),
    .A2(_09139_),
    .B(_09185_),
    .Y(_02737_));
 NAND2x1_ASAP7_75t_R _27703_ (.A(_05795_),
    .B(_08652_),
    .Y(_09186_));
 OA211x2_ASAP7_75t_R _27704_ (.A1(_05823_),
    .A2(_08652_),
    .B(_09142_),
    .C(_09186_),
    .Y(_09187_));
 AO21x1_ASAP7_75t_R _27705_ (.A1(_08709_),
    .A2(_09139_),
    .B(_09187_),
    .Y(_02738_));
 AO21x1_ASAP7_75t_R _27706_ (.A1(_05513_),
    .A2(_05950_),
    .B(_16138_),
    .Y(_09188_));
 OA211x2_ASAP7_75t_R _27707_ (.A1(net259),
    .A2(_08655_),
    .B(_09142_),
    .C(_09188_),
    .Y(_09189_));
 AO21x1_ASAP7_75t_R _27708_ (.A1(_08712_),
    .A2(_09139_),
    .B(_09189_),
    .Y(_02739_));
 OR2x2_ASAP7_75t_R _27709_ (.A(_16261_),
    .B(_08652_),
    .Y(_09190_));
 OA211x2_ASAP7_75t_R _27710_ (.A1(_16263_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09190_),
    .Y(_09191_));
 AOI21x1_ASAP7_75t_R _27711_ (.A1(_01658_),
    .A2(_09139_),
    .B(_09191_),
    .Y(_02740_));
 INVx1_ASAP7_75t_R _27712_ (.A(_01657_),
    .Y(_09192_));
 AO21x1_ASAP7_75t_R _27713_ (.A1(_05513_),
    .A2(_05950_),
    .B(_16378_),
    .Y(_09193_));
 OA211x2_ASAP7_75t_R _27714_ (.A1(net261),
    .A2(_08655_),
    .B(_09142_),
    .C(_09193_),
    .Y(_09194_));
 AO21x1_ASAP7_75t_R _27715_ (.A1(_09192_),
    .A2(_09139_),
    .B(_09194_),
    .Y(_02741_));
 NAND2x1_ASAP7_75t_R _27716_ (.A(_05861_),
    .B(_08655_),
    .Y(_09195_));
 OA211x2_ASAP7_75t_R _27717_ (.A1(_16509_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09195_),
    .Y(_09196_));
 AOI21x1_ASAP7_75t_R _27718_ (.A1(_01656_),
    .A2(_09139_),
    .B(_09196_),
    .Y(_02742_));
 AO21x1_ASAP7_75t_R _27719_ (.A1(_05513_),
    .A2(_05950_),
    .B(_16617_),
    .Y(_09197_));
 OA211x2_ASAP7_75t_R _27720_ (.A1(net258),
    .A2(_08655_),
    .B(_09142_),
    .C(_09197_),
    .Y(_09198_));
 AO21x1_ASAP7_75t_R _27721_ (.A1(_08734_),
    .A2(_09139_),
    .B(_09198_),
    .Y(_02743_));
 INVx1_ASAP7_75t_R _27722_ (.A(_01654_),
    .Y(_09199_));
 AO21x1_ASAP7_75t_R _27723_ (.A1(_05513_),
    .A2(_05950_),
    .B(_05877_),
    .Y(_09200_));
 OA211x2_ASAP7_75t_R _27724_ (.A1(net163),
    .A2(_08655_),
    .B(_09142_),
    .C(_09200_),
    .Y(_09201_));
 AO21x1_ASAP7_75t_R _27725_ (.A1(_09199_),
    .A2(_09139_),
    .B(_09201_),
    .Y(_02744_));
 NAND2x1_ASAP7_75t_R _27726_ (.A(_04624_),
    .B(_08655_),
    .Y(_09202_));
 OA211x2_ASAP7_75t_R _27727_ (.A1(_06498_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09202_),
    .Y(_09203_));
 AOI21x1_ASAP7_75t_R _27728_ (.A1(_01653_),
    .A2(_09139_),
    .B(_09203_),
    .Y(_02745_));
 NAND2x1_ASAP7_75t_R _27729_ (.A(_05892_),
    .B(_08655_),
    .Y(_09204_));
 OA211x2_ASAP7_75t_R _27730_ (.A1(_04747_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09204_),
    .Y(_09205_));
 AOI21x1_ASAP7_75t_R _27731_ (.A1(_01652_),
    .A2(_09139_),
    .B(_09205_),
    .Y(_02746_));
 AO21x1_ASAP7_75t_R _27732_ (.A1(_05513_),
    .A2(_05950_),
    .B(_04854_),
    .Y(_09206_));
 OA211x2_ASAP7_75t_R _27733_ (.A1(net2172),
    .A2(_08655_),
    .B(_09142_),
    .C(_09206_),
    .Y(_09207_));
 AO21x1_ASAP7_75t_R _27734_ (.A1(_08719_),
    .A2(_09139_),
    .B(_09207_),
    .Y(_02747_));
 NAND2x1_ASAP7_75t_R _27735_ (.A(_04965_),
    .B(_08655_),
    .Y(_09208_));
 OA211x2_ASAP7_75t_R _27736_ (.A1(_04968_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09208_),
    .Y(_09209_));
 AOI21x1_ASAP7_75t_R _27737_ (.A1(_01650_),
    .A2(_09139_),
    .B(_09209_),
    .Y(_02748_));
 NAND2x1_ASAP7_75t_R _27738_ (.A(_05075_),
    .B(_08655_),
    .Y(_09210_));
 OA211x2_ASAP7_75t_R _27739_ (.A1(_06526_),
    .A2(_08655_),
    .B(_09142_),
    .C(_09210_),
    .Y(_09211_));
 AOI21x1_ASAP7_75t_R _27740_ (.A1(_01649_),
    .A2(_09139_),
    .B(_09211_),
    .Y(_02749_));
 AO21x1_ASAP7_75t_R _27741_ (.A1(_05513_),
    .A2(_05950_),
    .B(_05924_),
    .Y(_09212_));
 OA211x2_ASAP7_75t_R _27742_ (.A1(net169),
    .A2(_08655_),
    .B(_09142_),
    .C(_09212_),
    .Y(_09213_));
 AO21x1_ASAP7_75t_R _27743_ (.A1(_08724_),
    .A2(_09139_),
    .B(_09213_),
    .Y(_02750_));
 AND2x2_ASAP7_75t_R _27744_ (.A(_05936_),
    .B(_08655_),
    .Y(_09214_));
 AO21x1_ASAP7_75t_R _27745_ (.A1(net2139),
    .A2(_08652_),
    .B(_09214_),
    .Y(_09215_));
 OR2x2_ASAP7_75t_R _27746_ (.A(_09139_),
    .B(_09215_),
    .Y(_09216_));
 OA21x2_ASAP7_75t_R _27747_ (.A1(_08727_),
    .A2(_09142_),
    .B(_09216_),
    .Y(_02751_));
 INVx1_ASAP7_75t_R _27748_ (.A(_01646_),
    .Y(_09217_));
 AO21x1_ASAP7_75t_R _27749_ (.A1(_05513_),
    .A2(_05950_),
    .B(_05400_),
    .Y(_09218_));
 OA211x2_ASAP7_75t_R _27750_ (.A1(net172),
    .A2(_08655_),
    .B(_09142_),
    .C(_09218_),
    .Y(_09219_));
 AO21x1_ASAP7_75t_R _27751_ (.A1(_09217_),
    .A2(_09139_),
    .B(_09219_),
    .Y(_02752_));
 OA211x2_ASAP7_75t_R _27752_ (.A1(net173),
    .A2(_05966_),
    .B(_09142_),
    .C(_05513_),
    .Y(_09220_));
 AO21x1_ASAP7_75t_R _27753_ (.A1(_08742_),
    .A2(_09139_),
    .B(_09220_),
    .Y(_02753_));
 AND3x4_ASAP7_75t_R _27754_ (.A(_05781_),
    .B(_01357_),
    .C(_05777_),
    .Y(_09221_));
 TAPCELL_ASAP7_75t_R PHY_631 ();
 TAPCELL_ASAP7_75t_R PHY_630 ();
 OR2x4_ASAP7_75t_R _27757_ (.A(_01321_),
    .B(_05808_),
    .Y(_09224_));
 OA21x2_ASAP7_75t_R _27758_ (.A1(_08752_),
    .A2(_09224_),
    .B(_01323_),
    .Y(_09225_));
 NOR2x1_ASAP7_75t_R _27759_ (.A(_09221_),
    .B(_09225_),
    .Y(_02754_));
 OA21x2_ASAP7_75t_R _27760_ (.A1(_05808_),
    .A2(_08768_),
    .B(_01324_),
    .Y(_09226_));
 NOR2x1_ASAP7_75t_R _27761_ (.A(_09221_),
    .B(_09226_),
    .Y(_02755_));
 OR2x6_ASAP7_75t_R _27762_ (.A(_01326_),
    .B(_05808_),
    .Y(_09227_));
 TAPCELL_ASAP7_75t_R PHY_629 ();
 OA21x2_ASAP7_75t_R _27764_ (.A1(_08752_),
    .A2(_09227_),
    .B(_01325_),
    .Y(_09229_));
 NOR2x1_ASAP7_75t_R _27765_ (.A(_09221_),
    .B(_09229_),
    .Y(_02756_));
 TAPCELL_ASAP7_75t_R PHY_628 ();
 OR2x6_ASAP7_75t_R _27767_ (.A(_01320_),
    .B(_05808_),
    .Y(_09231_));
 TAPCELL_ASAP7_75t_R PHY_627 ();
 OAI22x1_ASAP7_75t_R _27769_ (.A1(_01327_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_08752_),
    .Y(_02757_));
 OA21x2_ASAP7_75t_R _27770_ (.A1(_08822_),
    .A2(_09224_),
    .B(_01328_),
    .Y(_09233_));
 NOR2x1_ASAP7_75t_R _27771_ (.A(_09221_),
    .B(_09233_),
    .Y(_02758_));
 OR3x1_ASAP7_75t_R _27772_ (.A(_05774_),
    .B(_05808_),
    .C(_08821_),
    .Y(_09234_));
 AOI21x1_ASAP7_75t_R _27773_ (.A1(_01329_),
    .A2(_09234_),
    .B(_09221_),
    .Y(_02759_));
 OAI22x1_ASAP7_75t_R _27774_ (.A1(_01330_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_08822_),
    .Y(_02760_));
 OAI22x1_ASAP7_75t_R _27775_ (.A1(_01331_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_08822_),
    .Y(_02761_));
 OA21x2_ASAP7_75t_R _27776_ (.A1(_08874_),
    .A2(_09224_),
    .B(_01332_),
    .Y(_09235_));
 NOR2x1_ASAP7_75t_R _27777_ (.A(_09221_),
    .B(_09235_),
    .Y(_02762_));
 OR4x1_ASAP7_75t_R _27778_ (.A(_01322_),
    .B(_05774_),
    .C(_05808_),
    .D(_08884_),
    .Y(_09236_));
 AOI21x1_ASAP7_75t_R _27779_ (.A1(_01333_),
    .A2(_09236_),
    .B(_09221_),
    .Y(_02763_));
 OAI22x1_ASAP7_75t_R _27780_ (.A1(_01334_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_08874_),
    .Y(_02764_));
 TAPCELL_ASAP7_75t_R PHY_626 ();
 OAI22x1_ASAP7_75t_R _27782_ (.A1(_01335_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_08874_),
    .Y(_02765_));
 OR4x2_ASAP7_75t_R _27783_ (.A(_01321_),
    .B(_17825_),
    .C(_05808_),
    .D(_08746_),
    .Y(_09238_));
 OAI22x1_ASAP7_75t_R _27784_ (.A1(_01336_),
    .A2(_09221_),
    .B1(_09238_),
    .B2(_08873_),
    .Y(_02766_));
 OA21x2_ASAP7_75t_R _27785_ (.A1(_05808_),
    .A2(_08926_),
    .B(_01337_),
    .Y(_09239_));
 NOR2x1_ASAP7_75t_R _27786_ (.A(_09221_),
    .B(_09239_),
    .Y(_02767_));
 OAI22x1_ASAP7_75t_R _27787_ (.A1(_01338_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_08942_),
    .Y(_02768_));
 OAI22x1_ASAP7_75t_R _27788_ (.A1(_01339_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_08942_),
    .Y(_02769_));
 OAI22x1_ASAP7_75t_R _27789_ (.A1(_01340_),
    .A2(_09221_),
    .B1(_09224_),
    .B2(_08964_),
    .Y(_02770_));
 OA21x2_ASAP7_75t_R _27790_ (.A1(_05808_),
    .A2(_08972_),
    .B(_01341_),
    .Y(_09240_));
 NOR2x1_ASAP7_75t_R _27791_ (.A(_09221_),
    .B(_09240_),
    .Y(_02771_));
 OAI22x1_ASAP7_75t_R _27792_ (.A1(_01342_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_08964_),
    .Y(_02772_));
 OAI22x1_ASAP7_75t_R _27793_ (.A1(_01343_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_08964_),
    .Y(_02773_));
 OAI22x1_ASAP7_75t_R _27794_ (.A1(_01344_),
    .A2(_09221_),
    .B1(_09238_),
    .B2(_09001_),
    .Y(_02774_));
 OAI22x1_ASAP7_75t_R _27795_ (.A1(_05808_),
    .A2(_09013_),
    .B1(_09221_),
    .B2(_01345_),
    .Y(_02775_));
 OAI22x1_ASAP7_75t_R _27796_ (.A1(_01346_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_09022_),
    .Y(_02776_));
 OAI22x1_ASAP7_75t_R _27797_ (.A1(_01347_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_09022_),
    .Y(_02777_));
 OAI22x1_ASAP7_75t_R _27798_ (.A1(_01348_),
    .A2(_09221_),
    .B1(_09224_),
    .B2(_09045_),
    .Y(_02778_));
 OR3x1_ASAP7_75t_R _27799_ (.A(_05808_),
    .B(_08884_),
    .C(_09054_),
    .Y(_09241_));
 AOI21x1_ASAP7_75t_R _27800_ (.A1(_01349_),
    .A2(_09241_),
    .B(_09221_),
    .Y(_02779_));
 OAI22x1_ASAP7_75t_R _27801_ (.A1(_01350_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_09045_),
    .Y(_02780_));
 OAI22x1_ASAP7_75t_R _27802_ (.A1(_01351_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_09045_),
    .Y(_02781_));
 OR3x1_ASAP7_75t_R _27803_ (.A(_01318_),
    .B(_01322_),
    .C(_09238_),
    .Y(_09242_));
 OAI21x1_ASAP7_75t_R _27804_ (.A1(_01352_),
    .A2(_09221_),
    .B(_09242_),
    .Y(_02782_));
 OR4x1_ASAP7_75t_R _27805_ (.A(_17825_),
    .B(_05808_),
    .C(_08746_),
    .D(_09054_),
    .Y(_09243_));
 AOI21x1_ASAP7_75t_R _27806_ (.A1(_01353_),
    .A2(_09243_),
    .B(_09221_),
    .Y(_02783_));
 OAI22x1_ASAP7_75t_R _27807_ (.A1(_01354_),
    .A2(_09221_),
    .B1(_09227_),
    .B2(_09083_),
    .Y(_02784_));
 OAI22x1_ASAP7_75t_R _27808_ (.A1(_01355_),
    .A2(_09221_),
    .B1(_09231_),
    .B2(_09083_),
    .Y(_02785_));
 OR4x2_ASAP7_75t_R _27809_ (.A(_05781_),
    .B(_05782_),
    .C(_05776_),
    .D(_05769_),
    .Y(_09244_));
 OR2x2_ASAP7_75t_R _27810_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_05777_),
    .Y(_09245_));
 OA21x2_ASAP7_75t_R _27811_ (.A1(_17818_),
    .A2(_09244_),
    .B(_09245_),
    .Y(_02786_));
 OA22x2_ASAP7_75t_R _27812_ (.A1(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .A2(_05777_),
    .B1(_09244_),
    .B2(_02290_),
    .Y(_02787_));
 OA22x2_ASAP7_75t_R _27813_ (.A1(_08872_),
    .A2(_05777_),
    .B1(_09244_),
    .B2(_02293_),
    .Y(_02788_));
 OA22x2_ASAP7_75t_R _27814_ (.A1(_08819_),
    .A2(_05777_),
    .B1(_08672_),
    .B2(_09244_),
    .Y(_02789_));
 OA21x2_ASAP7_75t_R _27815_ (.A1(_08669_),
    .A2(_09244_),
    .B(_05777_),
    .Y(_09246_));
 OR4x1_ASAP7_75t_R _27816_ (.A(_01318_),
    .B(_02291_),
    .C(_05771_),
    .D(_09244_),
    .Y(_09247_));
 OA21x2_ASAP7_75t_R _27817_ (.A1(_05773_),
    .A2(_09246_),
    .B(_09247_),
    .Y(_02790_));
 AND2x2_ASAP7_75t_R _27818_ (.A(_05759_),
    .B(net218),
    .Y(_09248_));
 AO21x1_ASAP7_75t_R _27819_ (.A1(_05555_),
    .A2(_05758_),
    .B(_09248_),
    .Y(_02791_));
 AND4x2_ASAP7_75t_R _27820_ (.A(_00279_),
    .B(_00175_),
    .C(_14828_),
    .D(_05759_),
    .Y(_09249_));
 AO21x1_ASAP7_75t_R _27821_ (.A1(_07816_),
    .A2(_05758_),
    .B(_09249_),
    .Y(_02792_));
 OR2x2_ASAP7_75t_R _27822_ (.A(_07051_),
    .B(_05759_),
    .Y(_09250_));
 OA21x2_ASAP7_75t_R _27823_ (.A1(net298),
    .A2(_05758_),
    .B(_09250_),
    .Y(_02793_));
 OR2x2_ASAP7_75t_R _27824_ (.A(_07039_),
    .B(_05759_),
    .Y(_09251_));
 OA21x2_ASAP7_75t_R _27825_ (.A1(net297),
    .A2(_05758_),
    .B(_09251_),
    .Y(_02794_));
 NAND2x1_ASAP7_75t_R _27826_ (.A(net3055),
    .B(_01609_),
    .Y(_09252_));
 NOR2x1_ASAP7_75t_R _27827_ (.A(net2732),
    .B(_09252_),
    .Y(_09253_));
 AO21x1_ASAP7_75t_R _27828_ (.A1(_01607_),
    .A2(_13446_),
    .B(_09253_),
    .Y(_09254_));
 OA22x2_ASAP7_75t_R _27829_ (.A1(_13444_),
    .A2(_05753_),
    .B1(_09254_),
    .B2(_01608_),
    .Y(_09255_));
 AND2x2_ASAP7_75t_R _27830_ (.A(_13448_),
    .B(_01608_),
    .Y(_09256_));
 AO32x2_ASAP7_75t_R _27831_ (.A1(_00277_),
    .A2(net2728),
    .A3(_09255_),
    .B1(_09256_),
    .B2(_09253_),
    .Y(_09257_));
 TAPCELL_ASAP7_75t_R PHY_625 ();
 TAPCELL_ASAP7_75t_R PHY_624 ();
 TAPCELL_ASAP7_75t_R PHY_623 ();
 NOR2x1_ASAP7_75t_R _27835_ (.A(_01641_),
    .B(_09257_),
    .Y(_09261_));
 AO21x1_ASAP7_75t_R _27836_ (.A1(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A2(_09257_),
    .B(_09261_),
    .Y(_02795_));
 NOR2x1_ASAP7_75t_R _27837_ (.A(_01640_),
    .B(_09257_),
    .Y(_09262_));
 AO21x1_ASAP7_75t_R _27838_ (.A1(\ex_block_i.alu_adder_result_ex_o[1] ),
    .A2(_09257_),
    .B(_09262_),
    .Y(_02796_));
 TAPCELL_ASAP7_75t_R PHY_622 ();
 NOR2x1_ASAP7_75t_R _27840_ (.A(_01639_),
    .B(_09257_),
    .Y(_09264_));
 AO21x1_ASAP7_75t_R _27841_ (.A1(net171),
    .A2(_09257_),
    .B(_09264_),
    .Y(_02797_));
 NOR2x1_ASAP7_75t_R _27842_ (.A(_01638_),
    .B(_09257_),
    .Y(_09265_));
 AO21x1_ASAP7_75t_R _27843_ (.A1(net293),
    .A2(_09257_),
    .B(_09265_),
    .Y(_02798_));
 NOR2x1_ASAP7_75t_R _27844_ (.A(_01637_),
    .B(_09257_),
    .Y(_09266_));
 AO21x1_ASAP7_75t_R _27845_ (.A1(net175),
    .A2(_09257_),
    .B(_09266_),
    .Y(_02799_));
 NOR2x1_ASAP7_75t_R _27846_ (.A(_01636_),
    .B(_09257_),
    .Y(_09267_));
 AO21x1_ASAP7_75t_R _27847_ (.A1(net289),
    .A2(_09257_),
    .B(_09267_),
    .Y(_02800_));
 NOR2x1_ASAP7_75t_R _27848_ (.A(_01635_),
    .B(_09257_),
    .Y(_09268_));
 AO21x1_ASAP7_75t_R _27849_ (.A1(net177),
    .A2(_09257_),
    .B(_09268_),
    .Y(_02801_));
 TAPCELL_ASAP7_75t_R PHY_621 ();
 NAND2x1_ASAP7_75t_R _27851_ (.A(_00676_),
    .B(_09257_),
    .Y(_09270_));
 OA21x2_ASAP7_75t_R _27852_ (.A1(_15224_),
    .A2(_09257_),
    .B(_09270_),
    .Y(_02802_));
 NAND2x1_ASAP7_75t_R _27853_ (.A(_05798_),
    .B(_09257_),
    .Y(_09271_));
 OA21x2_ASAP7_75t_R _27854_ (.A1(_15229_),
    .A2(_09257_),
    .B(_09271_),
    .Y(_02803_));
 NOR2x1_ASAP7_75t_R _27855_ (.A(_01632_),
    .B(_09257_),
    .Y(_09272_));
 AO21x1_ASAP7_75t_R _27856_ (.A1(net2205),
    .A2(_09257_),
    .B(_09272_),
    .Y(_02804_));
 NOR2x1_ASAP7_75t_R _27857_ (.A(_01631_),
    .B(_09257_),
    .Y(_09273_));
 AO21x1_ASAP7_75t_R _27858_ (.A1(net151),
    .A2(_09257_),
    .B(_09273_),
    .Y(_02805_));
 NOR2x1_ASAP7_75t_R _27859_ (.A(_01630_),
    .B(_09257_),
    .Y(_09274_));
 AO21x1_ASAP7_75t_R _27860_ (.A1(net262),
    .A2(_09257_),
    .B(_09274_),
    .Y(_02806_));
 TAPCELL_ASAP7_75t_R PHY_620 ();
 NOR2x1_ASAP7_75t_R _27862_ (.A(_01629_),
    .B(_09257_),
    .Y(_09276_));
 AO21x1_ASAP7_75t_R _27863_ (.A1(net153),
    .A2(_09257_),
    .B(_09276_),
    .Y(_02807_));
 NOR2x1_ASAP7_75t_R _27864_ (.A(_01628_),
    .B(_09257_),
    .Y(_09277_));
 AO21x1_ASAP7_75t_R _27865_ (.A1(net154),
    .A2(_09257_),
    .B(_09277_),
    .Y(_02808_));
 TAPCELL_ASAP7_75t_R PHY_619 ();
 NOR2x1_ASAP7_75t_R _27867_ (.A(_01627_),
    .B(_09257_),
    .Y(_09279_));
 AO21x1_ASAP7_75t_R _27868_ (.A1(net155),
    .A2(_09257_),
    .B(_09279_),
    .Y(_02809_));
 NAND2x1_ASAP7_75t_R _27869_ (.A(net260),
    .B(_09257_),
    .Y(_09280_));
 OA21x2_ASAP7_75t_R _27870_ (.A1(_15886_),
    .A2(_09257_),
    .B(_09280_),
    .Y(_02810_));
 INVx1_ASAP7_75t_R _27871_ (.A(_01625_),
    .Y(_09281_));
 NAND2x1_ASAP7_75t_R _27872_ (.A(_05795_),
    .B(_09257_),
    .Y(_09282_));
 OA21x2_ASAP7_75t_R _27873_ (.A1(_09281_),
    .A2(_09257_),
    .B(_09282_),
    .Y(_02811_));
 NOR2x1_ASAP7_75t_R _27874_ (.A(_01624_),
    .B(_09257_),
    .Y(_09283_));
 AO21x1_ASAP7_75t_R _27875_ (.A1(net259),
    .A2(_09257_),
    .B(_09283_),
    .Y(_02812_));
 NOR2x1_ASAP7_75t_R _27876_ (.A(_01623_),
    .B(_09257_),
    .Y(_09284_));
 AO21x1_ASAP7_75t_R _27877_ (.A1(net159),
    .A2(_09257_),
    .B(_09284_),
    .Y(_02813_));
 NOR2x1_ASAP7_75t_R _27878_ (.A(_01622_),
    .B(_09257_),
    .Y(_09285_));
 AO21x1_ASAP7_75t_R _27879_ (.A1(net261),
    .A2(_09257_),
    .B(_09285_),
    .Y(_02814_));
 NOR2x1_ASAP7_75t_R _27880_ (.A(_01621_),
    .B(_09257_),
    .Y(_09286_));
 AO21x1_ASAP7_75t_R _27881_ (.A1(net161),
    .A2(_09257_),
    .B(_09286_),
    .Y(_02815_));
 NOR2x1_ASAP7_75t_R _27882_ (.A(_01620_),
    .B(_09257_),
    .Y(_09287_));
 AO21x1_ASAP7_75t_R _27883_ (.A1(net258),
    .A2(_09257_),
    .B(_09287_),
    .Y(_02816_));
 NAND2x1_ASAP7_75t_R _27884_ (.A(_04517_),
    .B(_09257_),
    .Y(_09288_));
 OA21x2_ASAP7_75t_R _27885_ (.A1(_04515_),
    .A2(_09257_),
    .B(_09288_),
    .Y(_02817_));
 NOR2x1_ASAP7_75t_R _27886_ (.A(_01618_),
    .B(_09257_),
    .Y(_09289_));
 AO21x1_ASAP7_75t_R _27887_ (.A1(net2180),
    .A2(_09257_),
    .B(_09289_),
    .Y(_02818_));
 NOR2x1_ASAP7_75t_R _27888_ (.A(_01617_),
    .B(_09257_),
    .Y(_09290_));
 AO21x1_ASAP7_75t_R _27889_ (.A1(net165),
    .A2(_09257_),
    .B(_09290_),
    .Y(_02819_));
 NOR2x1_ASAP7_75t_R _27890_ (.A(_01616_),
    .B(_09257_),
    .Y(_09291_));
 AO21x1_ASAP7_75t_R _27891_ (.A1(net2174),
    .A2(_09257_),
    .B(_09291_),
    .Y(_02820_));
 INVx1_ASAP7_75t_R _27892_ (.A(_01615_),
    .Y(_09292_));
 NAND2x1_ASAP7_75t_R _27893_ (.A(_04968_),
    .B(_09257_),
    .Y(_09293_));
 OA21x2_ASAP7_75t_R _27894_ (.A1(_09292_),
    .A2(_09257_),
    .B(_09293_),
    .Y(_02821_));
 NOR2x1_ASAP7_75t_R _27895_ (.A(_01614_),
    .B(_09257_),
    .Y(_09294_));
 AO21x1_ASAP7_75t_R _27896_ (.A1(net2154),
    .A2(_09257_),
    .B(_09294_),
    .Y(_02822_));
 INVx1_ASAP7_75t_R _27897_ (.A(_01613_),
    .Y(_09295_));
 NAND2x1_ASAP7_75t_R _27898_ (.A(_05185_),
    .B(_09257_),
    .Y(_09296_));
 OA21x2_ASAP7_75t_R _27899_ (.A1(_09295_),
    .A2(_09257_),
    .B(_09296_),
    .Y(_02823_));
 NOR2x1_ASAP7_75t_R _27900_ (.A(_01612_),
    .B(_09257_),
    .Y(_09297_));
 AO21x1_ASAP7_75t_R _27901_ (.A1(net2140),
    .A2(_09257_),
    .B(_09297_),
    .Y(_02824_));
 NAND2x1_ASAP7_75t_R _27902_ (.A(_05404_),
    .B(_09257_),
    .Y(_09298_));
 OA21x2_ASAP7_75t_R _27903_ (.A1(_05402_),
    .A2(_09257_),
    .B(_09298_),
    .Y(_02825_));
 NOR2x1_ASAP7_75t_R _27904_ (.A(_01610_),
    .B(_09257_),
    .Y(_09299_));
 AO21x1_ASAP7_75t_R _27905_ (.A1(net173),
    .A2(_09257_),
    .B(_09299_),
    .Y(_02826_));
 AO21x1_ASAP7_75t_R _27906_ (.A1(net3055),
    .A2(_13509_),
    .B(_05754_),
    .Y(_09300_));
 INVx1_ASAP7_75t_R _27907_ (.A(net3030),
    .Y(_09301_));
 OA211x2_ASAP7_75t_R _27908_ (.A1(_13446_),
    .A2(_09300_),
    .B(_00277_),
    .C(net3031),
    .Y(_02827_));
 OR3x1_ASAP7_75t_R _27909_ (.A(_00281_),
    .B(_02537_),
    .C(_06189_),
    .Y(_09302_));
 OA211x2_ASAP7_75t_R _27910_ (.A1(_06114_),
    .A2(_05763_),
    .B(_09302_),
    .C(_01609_),
    .Y(_09303_));
 INVx1_ASAP7_75t_R _27911_ (.A(_09303_),
    .Y(_09304_));
 OA21x2_ASAP7_75t_R _27912_ (.A1(_13446_),
    .A2(_05753_),
    .B(net3030),
    .Y(_09305_));
 AO21x1_ASAP7_75t_R _27913_ (.A1(_05753_),
    .A2(_09303_),
    .B(_13509_),
    .Y(_09306_));
 AO32x1_ASAP7_75t_R _27914_ (.A1(_01608_),
    .A2(_09304_),
    .A3(_09305_),
    .B1(_09306_),
    .B2(net3031),
    .Y(_09307_));
 AND2x2_ASAP7_75t_R _27915_ (.A(_00277_),
    .B(_09307_),
    .Y(_02828_));
 NOR2x1_ASAP7_75t_R _27916_ (.A(_01608_),
    .B(_05757_),
    .Y(_09308_));
 INVx1_ASAP7_75t_R _27917_ (.A(net3055),
    .Y(_09309_));
 OA211x2_ASAP7_75t_R _27918_ (.A1(_09256_),
    .A2(_09308_),
    .B(net2805),
    .C(_01609_),
    .Y(_02829_));
 AND3x1_ASAP7_75t_R _27919_ (.A(_13448_),
    .B(net3055),
    .C(_01608_),
    .Y(_09310_));
 AO21x1_ASAP7_75t_R _27920_ (.A1(_00277_),
    .A2(_09300_),
    .B(_09310_),
    .Y(_09311_));
 AND2x2_ASAP7_75t_R _27921_ (.A(_01609_),
    .B(_09311_),
    .Y(_09312_));
 XOR2x2_ASAP7_75t_R _27922_ (.A(_00277_),
    .B(_01608_),
    .Y(_09313_));
 AND3x1_ASAP7_75t_R _27923_ (.A(net3036),
    .B(_09312_),
    .C(_09313_),
    .Y(_09314_));
 INVx1_ASAP7_75t_R _27924_ (.A(net2733),
    .Y(_09315_));
 OAI21x1_ASAP7_75t_R _27925_ (.A1(_01607_),
    .A2(_09312_),
    .B(net2734),
    .Y(_02830_));
 AOI21x1_ASAP7_75t_R _27926_ (.A1(net3031),
    .A2(_09252_),
    .B(_01608_),
    .Y(_09316_));
 OAI21x1_ASAP7_75t_R _27927_ (.A1(_09305_),
    .A2(_09316_),
    .B(_00277_),
    .Y(_09317_));
 AO32x1_ASAP7_75t_R _27928_ (.A1(_00277_),
    .A2(net3030),
    .A3(_09306_),
    .B1(_09317_),
    .B2(_18554_),
    .Y(_09318_));
 INVx1_ASAP7_75t_R _27929_ (.A(_09318_),
    .Y(_02831_));
 NAND2x2_ASAP7_75t_R _27930_ (.A(_06618_),
    .B(_06685_),
    .Y(_09319_));
 TAPCELL_ASAP7_75t_R PHY_618 ();
 TAPCELL_ASAP7_75t_R PHY_617 ();
 TAPCELL_ASAP7_75t_R PHY_616 ();
 TAPCELL_ASAP7_75t_R PHY_615 ();
 AND3x1_ASAP7_75t_R _27935_ (.A(_06676_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09324_));
 TAPCELL_ASAP7_75t_R PHY_614 ();
 TAPCELL_ASAP7_75t_R PHY_613 ();
 OAI22x1_ASAP7_75t_R _27938_ (.A1(net255),
    .A2(_06722_),
    .B1(_09324_),
    .B2(_00662_),
    .Y(_09327_));
 TAPCELL_ASAP7_75t_R PHY_612 ();
 AND3x1_ASAP7_75t_R _27940_ (.A(\ex_block_i.alu_adder_result_ex_o[1] ),
    .B(_14791_),
    .C(_14794_),
    .Y(_09329_));
 OAI22x1_ASAP7_75t_R _27941_ (.A1(_01944_),
    .A2(_06301_),
    .B1(_06308_),
    .B2(_00658_),
    .Y(_09330_));
 OR3x2_ASAP7_75t_R _27942_ (.A(_06273_),
    .B(_09329_),
    .C(_09330_),
    .Y(_09331_));
 OA21x2_ASAP7_75t_R _27943_ (.A1(_06296_),
    .A2(_09327_),
    .B(_09331_),
    .Y(_02832_));
 INVx1_ASAP7_75t_R _27944_ (.A(_00241_),
    .Y(_09332_));
 TAPCELL_ASAP7_75t_R PHY_611 ();
 TAPCELL_ASAP7_75t_R PHY_610 ();
 AO21x1_ASAP7_75t_R _27947_ (.A1(_06618_),
    .A2(_06685_),
    .B(_17754_),
    .Y(_09335_));
 OA211x2_ASAP7_75t_R _27948_ (.A1(_09332_),
    .A2(net255),
    .B(_09335_),
    .C(net300),
    .Y(_09336_));
 NOR2x1_ASAP7_75t_R _27949_ (.A(net3391),
    .B(_09336_),
    .Y(_02833_));
 TAPCELL_ASAP7_75t_R PHY_609 ();
 TAPCELL_ASAP7_75t_R PHY_608 ();
 AND3x1_ASAP7_75t_R _27952_ (.A(_02539_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09339_));
 AO21x1_ASAP7_75t_R _27953_ (.A1(_01606_),
    .A2(net255),
    .B(_09339_),
    .Y(_09340_));
 AOI21x1_ASAP7_75t_R _27954_ (.A1(net300),
    .A2(_09340_),
    .B(net3511),
    .Y(_02834_));
 INVx1_ASAP7_75t_R _27955_ (.A(_02538_),
    .Y(_09341_));
 AND3x1_ASAP7_75t_R _27956_ (.A(_09341_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09342_));
 XOR2x1_ASAP7_75t_R _27957_ (.A(_01605_),
    .Y(_09343_),
    .B(_09342_));
 AOI21x1_ASAP7_75t_R _27958_ (.A1(net300),
    .A2(_09343_),
    .B(net3503),
    .Y(_02835_));
 AND3x1_ASAP7_75t_R _27959_ (.A(_02541_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09344_));
 AO21x1_ASAP7_75t_R _27960_ (.A1(_01604_),
    .A2(net255),
    .B(_09344_),
    .Y(_09345_));
 AOI21x1_ASAP7_75t_R _27961_ (.A1(net300),
    .A2(_09345_),
    .B(_06352_),
    .Y(_02836_));
 INVx1_ASAP7_75t_R _27962_ (.A(_02540_),
    .Y(_09346_));
 AND3x1_ASAP7_75t_R _27963_ (.A(_09346_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09347_));
 XOR2x1_ASAP7_75t_R _27964_ (.A(_01603_),
    .Y(_09348_),
    .B(_09347_));
 AOI21x1_ASAP7_75t_R _27965_ (.A1(net300),
    .A2(_09348_),
    .B(_06362_),
    .Y(_02837_));
 NOR2x1_ASAP7_75t_R _27966_ (.A(net300),
    .B(_06376_),
    .Y(_09349_));
 INVx1_ASAP7_75t_R _27967_ (.A(_02543_),
    .Y(_09350_));
 TAPCELL_ASAP7_75t_R PHY_607 ();
 TAPCELL_ASAP7_75t_R PHY_606 ();
 AO21x1_ASAP7_75t_R _27970_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[7] ),
    .Y(_09353_));
 OA211x2_ASAP7_75t_R _27971_ (.A1(_09350_),
    .A2(net255),
    .B(_09353_),
    .C(net300),
    .Y(_09354_));
 OR2x2_ASAP7_75t_R _27972_ (.A(_09349_),
    .B(_09354_),
    .Y(_02838_));
 INVx1_ASAP7_75t_R _27973_ (.A(_02542_),
    .Y(_09355_));
 AND3x1_ASAP7_75t_R _27974_ (.A(_09355_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09356_));
 XOR2x1_ASAP7_75t_R _27975_ (.A(_01601_),
    .Y(_09357_),
    .B(_09356_));
 AOI21x1_ASAP7_75t_R _27976_ (.A1(net300),
    .A2(_09357_),
    .B(net3090),
    .Y(_02839_));
 AND3x1_ASAP7_75t_R _27977_ (.A(_02545_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09358_));
 AO21x1_ASAP7_75t_R _27978_ (.A1(_01600_),
    .A2(_09319_),
    .B(_09358_),
    .Y(_09359_));
 OAI21x1_ASAP7_75t_R _27979_ (.A1(net299),
    .A2(_09359_),
    .B(_06396_),
    .Y(_02840_));
 INVx1_ASAP7_75t_R _27980_ (.A(_02544_),
    .Y(_09360_));
 AND3x1_ASAP7_75t_R _27981_ (.A(_09360_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09361_));
 XOR2x1_ASAP7_75t_R _27982_ (.A(_01599_),
    .Y(_09362_),
    .B(_09361_));
 AOI21x1_ASAP7_75t_R _27983_ (.A1(net300),
    .A2(_09362_),
    .B(_06403_),
    .Y(_02841_));
 AND3x1_ASAP7_75t_R _27984_ (.A(_02547_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09363_));
 AO21x1_ASAP7_75t_R _27985_ (.A1(_01598_),
    .A2(_09319_),
    .B(_09363_),
    .Y(_09364_));
 OAI21x1_ASAP7_75t_R _27986_ (.A1(net299),
    .A2(_09364_),
    .B(_06416_),
    .Y(_02842_));
 INVx1_ASAP7_75t_R _27987_ (.A(_02546_),
    .Y(_09365_));
 AND3x1_ASAP7_75t_R _27988_ (.A(_09365_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09366_));
 XOR2x1_ASAP7_75t_R _27989_ (.A(_01597_),
    .Y(_09367_),
    .B(_09366_));
 AOI21x1_ASAP7_75t_R _27990_ (.A1(net301),
    .A2(_09367_),
    .B(_06425_),
    .Y(_02843_));
 INVx1_ASAP7_75t_R _27991_ (.A(_02549_),
    .Y(_09368_));
 AO21x1_ASAP7_75t_R _27992_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .Y(_09369_));
 OA211x2_ASAP7_75t_R _27993_ (.A1(_09368_),
    .A2(net255),
    .B(_09369_),
    .C(net300),
    .Y(_09370_));
 OR2x2_ASAP7_75t_R _27994_ (.A(_06433_),
    .B(_09370_),
    .Y(_02844_));
 INVx1_ASAP7_75t_R _27995_ (.A(_02548_),
    .Y(_09371_));
 AND3x1_ASAP7_75t_R _27996_ (.A(_09371_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09372_));
 XOR2x1_ASAP7_75t_R _27997_ (.A(_01595_),
    .Y(_09373_),
    .B(_09372_));
 AOI21x1_ASAP7_75t_R _27998_ (.A1(net301),
    .A2(_09373_),
    .B(net3168),
    .Y(_02845_));
 NOR2x1_ASAP7_75t_R _27999_ (.A(net300),
    .B(_06445_),
    .Y(_09374_));
 INVx1_ASAP7_75t_R _28000_ (.A(_02551_),
    .Y(_09375_));
 AO21x1_ASAP7_75t_R _28001_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[15] ),
    .Y(_09376_));
 OA211x2_ASAP7_75t_R _28002_ (.A1(_09375_),
    .A2(_09319_),
    .B(_09376_),
    .C(net300),
    .Y(_09377_));
 OR2x2_ASAP7_75t_R _28003_ (.A(_09374_),
    .B(_09377_),
    .Y(_02846_));
 INVx1_ASAP7_75t_R _28004_ (.A(_02550_),
    .Y(_09378_));
 AND3x1_ASAP7_75t_R _28005_ (.A(_09378_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09379_));
 XOR2x1_ASAP7_75t_R _28006_ (.A(_01593_),
    .Y(_09380_),
    .B(_09379_));
 AOI21x1_ASAP7_75t_R _28007_ (.A1(net301),
    .A2(_09380_),
    .B(_06455_),
    .Y(_02847_));
 NOR2x1_ASAP7_75t_R _28008_ (.A(net301),
    .B(_06461_),
    .Y(_09381_));
 INVx1_ASAP7_75t_R _28009_ (.A(_02553_),
    .Y(_09382_));
 AO21x1_ASAP7_75t_R _28010_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[17] ),
    .Y(_09383_));
 OA211x2_ASAP7_75t_R _28011_ (.A1(_09382_),
    .A2(_09319_),
    .B(_09383_),
    .C(net301),
    .Y(_09384_));
 OR2x2_ASAP7_75t_R _28012_ (.A(_09381_),
    .B(_09384_),
    .Y(_02848_));
 NOR2x1_ASAP7_75t_R _28013_ (.A(_02552_),
    .B(_09319_),
    .Y(_09385_));
 NAND2x1_ASAP7_75t_R _28014_ (.A(_01591_),
    .B(net301),
    .Y(_09386_));
 OR4x1_ASAP7_75t_R _28015_ (.A(_01591_),
    .B(_02552_),
    .C(net299),
    .D(_09319_),
    .Y(_09387_));
 INVx1_ASAP7_75t_R _28016_ (.A(_06469_),
    .Y(_09388_));
 OA211x2_ASAP7_75t_R _28017_ (.A1(_09385_),
    .A2(_09386_),
    .B(_09387_),
    .C(_09388_),
    .Y(_02849_));
 AND3x1_ASAP7_75t_R _28018_ (.A(_02555_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09389_));
 AO21x1_ASAP7_75t_R _28019_ (.A1(_01590_),
    .A2(_09319_),
    .B(_09389_),
    .Y(_09390_));
 AOI21x1_ASAP7_75t_R _28020_ (.A1(_06273_),
    .A2(_09390_),
    .B(_06475_),
    .Y(_02850_));
 NOR2x1_ASAP7_75t_R _28021_ (.A(_02554_),
    .B(_09319_),
    .Y(_09391_));
 NAND2x1_ASAP7_75t_R _28022_ (.A(_01589_),
    .B(_06273_),
    .Y(_09392_));
 OR4x1_ASAP7_75t_R _28023_ (.A(_01589_),
    .B(_02554_),
    .C(net299),
    .D(_09319_),
    .Y(_09393_));
 INVx1_ASAP7_75t_R _28024_ (.A(_06482_),
    .Y(_09394_));
 OA211x2_ASAP7_75t_R _28025_ (.A1(_09391_),
    .A2(_09392_),
    .B(_09393_),
    .C(_09394_),
    .Y(_02851_));
 AND3x1_ASAP7_75t_R _28026_ (.A(_02557_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09395_));
 AO21x1_ASAP7_75t_R _28027_ (.A1(_01588_),
    .A2(_09319_),
    .B(_09395_),
    .Y(_09396_));
 AOI21x1_ASAP7_75t_R _28028_ (.A1(_06273_),
    .A2(_09396_),
    .B(_06489_),
    .Y(_02852_));
 TAPCELL_ASAP7_75t_R PHY_605 ();
 NOR2x1_ASAP7_75t_R _28030_ (.A(_02556_),
    .B(_09319_),
    .Y(_09398_));
 TAPCELL_ASAP7_75t_R PHY_604 ();
 NAND2x1_ASAP7_75t_R _28032_ (.A(_01587_),
    .B(_06273_),
    .Y(_09400_));
 OR4x1_ASAP7_75t_R _28033_ (.A(_01587_),
    .B(_02556_),
    .C(net299),
    .D(_09319_),
    .Y(_09401_));
 INVx1_ASAP7_75t_R _28034_ (.A(_06495_),
    .Y(_09402_));
 OA211x2_ASAP7_75t_R _28035_ (.A1(_09398_),
    .A2(_09400_),
    .B(_09401_),
    .C(_09402_),
    .Y(_02853_));
 NOR2x1_ASAP7_75t_R _28036_ (.A(net301),
    .B(_06501_),
    .Y(_09403_));
 INVx1_ASAP7_75t_R _28037_ (.A(_02559_),
    .Y(_09404_));
 AO21x1_ASAP7_75t_R _28038_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[23] ),
    .Y(_09405_));
 OA211x2_ASAP7_75t_R _28039_ (.A1(_09404_),
    .A2(net255),
    .B(_09405_),
    .C(net301),
    .Y(_09406_));
 OR2x2_ASAP7_75t_R _28040_ (.A(_09403_),
    .B(_09406_),
    .Y(_02854_));
 INVx1_ASAP7_75t_R _28041_ (.A(_02558_),
    .Y(_09407_));
 AND3x1_ASAP7_75t_R _28042_ (.A(_09407_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09408_));
 XOR2x1_ASAP7_75t_R _28043_ (.A(_01585_),
    .Y(_09409_),
    .B(_09408_));
 AOI21x1_ASAP7_75t_R _28044_ (.A1(net301),
    .A2(_09409_),
    .B(_06508_),
    .Y(_02855_));
 NOR2x1_ASAP7_75t_R _28045_ (.A(_06273_),
    .B(_06515_),
    .Y(_09410_));
 INVx1_ASAP7_75t_R _28046_ (.A(_02561_),
    .Y(_09411_));
 AO21x1_ASAP7_75t_R _28047_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[25] ),
    .Y(_09412_));
 OA211x2_ASAP7_75t_R _28048_ (.A1(_09411_),
    .A2(net255),
    .B(_09412_),
    .C(_06273_),
    .Y(_09413_));
 OR2x2_ASAP7_75t_R _28049_ (.A(_09410_),
    .B(_09413_),
    .Y(_02856_));
 NOR2x1_ASAP7_75t_R _28050_ (.A(_02560_),
    .B(_09319_),
    .Y(_09414_));
 NAND2x1_ASAP7_75t_R _28051_ (.A(_01583_),
    .B(_06273_),
    .Y(_09415_));
 OR4x1_ASAP7_75t_R _28052_ (.A(_01583_),
    .B(_02560_),
    .C(net299),
    .D(_09319_),
    .Y(_09416_));
 INVx1_ASAP7_75t_R _28053_ (.A(_06523_),
    .Y(_09417_));
 OA211x2_ASAP7_75t_R _28054_ (.A1(_09414_),
    .A2(_09415_),
    .B(_09416_),
    .C(_09417_),
    .Y(_02857_));
 NOR2x1_ASAP7_75t_R _28055_ (.A(_06273_),
    .B(_06530_),
    .Y(_09418_));
 INVx1_ASAP7_75t_R _28056_ (.A(_02563_),
    .Y(_09419_));
 AO21x1_ASAP7_75t_R _28057_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_if_i[27] ),
    .Y(_09420_));
 OA211x2_ASAP7_75t_R _28058_ (.A1(_09419_),
    .A2(net255),
    .B(_09420_),
    .C(_06273_),
    .Y(_09421_));
 OR2x2_ASAP7_75t_R _28059_ (.A(_09418_),
    .B(_09421_),
    .Y(_02858_));
 NOR2x1_ASAP7_75t_R _28060_ (.A(_02562_),
    .B(net255),
    .Y(_09422_));
 NAND2x1_ASAP7_75t_R _28061_ (.A(_01581_),
    .B(_06273_),
    .Y(_09423_));
 OR4x1_ASAP7_75t_R _28062_ (.A(_01581_),
    .B(_02562_),
    .C(net299),
    .D(net255),
    .Y(_09424_));
 INVx1_ASAP7_75t_R _28063_ (.A(_06538_),
    .Y(_09425_));
 OA211x2_ASAP7_75t_R _28064_ (.A1(_09422_),
    .A2(_09423_),
    .B(_09424_),
    .C(_09425_),
    .Y(_02859_));
 AND3x1_ASAP7_75t_R _28065_ (.A(_02565_),
    .B(_06618_),
    .C(_06685_),
    .Y(_09426_));
 AO21x1_ASAP7_75t_R _28066_ (.A1(_01580_),
    .A2(net255),
    .B(_09426_),
    .Y(_09427_));
 AOI21x1_ASAP7_75t_R _28067_ (.A1(_06273_),
    .A2(_09427_),
    .B(_06544_),
    .Y(_02860_));
 NOR2x1_ASAP7_75t_R _28068_ (.A(_02564_),
    .B(net255),
    .Y(_09428_));
 NAND2x1_ASAP7_75t_R _28069_ (.A(_01579_),
    .B(_06273_),
    .Y(_09429_));
 OR4x1_ASAP7_75t_R _28070_ (.A(_01579_),
    .B(_02564_),
    .C(net299),
    .D(net255),
    .Y(_09430_));
 INVx1_ASAP7_75t_R _28071_ (.A(_06550_),
    .Y(_09431_));
 OA211x2_ASAP7_75t_R _28072_ (.A1(_09428_),
    .A2(_09429_),
    .B(_09430_),
    .C(_09431_),
    .Y(_02861_));
 OR3x1_ASAP7_75t_R _28073_ (.A(_01579_),
    .B(_01580_),
    .C(_06606_),
    .Y(_09432_));
 AO22x1_ASAP7_75t_R _28074_ (.A1(_06273_),
    .A2(net255),
    .B1(_09432_),
    .B2(net3065),
    .Y(_09433_));
 NOR2x1_ASAP7_75t_R _28075_ (.A(_01578_),
    .B(_09432_),
    .Y(_09434_));
 AO21x1_ASAP7_75t_R _28076_ (.A1(_06686_),
    .A2(_09434_),
    .B(net299),
    .Y(_09435_));
 AOI22x1_ASAP7_75t_R _28077_ (.A1(_01578_),
    .A2(_09433_),
    .B1(_09435_),
    .B2(net3065),
    .Y(_02862_));
 OR4x2_ASAP7_75t_R _28078_ (.A(_05563_),
    .B(_07928_),
    .C(_05589_),
    .D(_06997_),
    .Y(_09436_));
 AO221x1_ASAP7_75t_R _28079_ (.A1(_06938_),
    .A2(_07359_),
    .B1(_07699_),
    .B2(_05656_),
    .C(_06940_),
    .Y(_09437_));
 AND3x1_ASAP7_75t_R _28080_ (.A(_06941_),
    .B(_06971_),
    .C(_06972_),
    .Y(_09438_));
 AND3x1_ASAP7_75t_R _28081_ (.A(_14296_),
    .B(_06973_),
    .C(_05678_),
    .Y(_09439_));
 AND3x1_ASAP7_75t_R _28082_ (.A(_05588_),
    .B(_05663_),
    .C(_09439_),
    .Y(_09440_));
 OR5x1_ASAP7_75t_R _28083_ (.A(_06961_),
    .B(_06963_),
    .C(_06969_),
    .D(_09438_),
    .E(_09440_),
    .Y(_09441_));
 OR5x2_ASAP7_75t_R _28084_ (.A(_06958_),
    .B(_09437_),
    .C(_06944_),
    .D(_07700_),
    .E(_09441_),
    .Y(_09442_));
 AND3x4_ASAP7_75t_R _28085_ (.A(_02288_),
    .B(_05737_),
    .C(_05739_),
    .Y(_09443_));
 TAPCELL_ASAP7_75t_R PHY_603 ();
 NAND2x2_ASAP7_75t_R _28087_ (.A(_09442_),
    .B(_09443_),
    .Y(_09445_));
 NOR2x2_ASAP7_75t_R _28088_ (.A(_09436_),
    .B(_09445_),
    .Y(_09446_));
 TAPCELL_ASAP7_75t_R PHY_602 ();
 TAPCELL_ASAP7_75t_R PHY_601 ();
 NOR2x1_ASAP7_75t_R _28091_ (.A(_18332_),
    .B(_14714_),
    .Y(_09449_));
 AO21x1_ASAP7_75t_R _28092_ (.A1(net306),
    .A2(_18332_),
    .B(_09449_),
    .Y(_09450_));
 TAPCELL_ASAP7_75t_R PHY_600 ();
 AOI22x1_ASAP7_75t_R _28094_ (.A1(_18332_),
    .A2(_07381_),
    .B1(_09450_),
    .B2(net307),
    .Y(_09452_));
 TAPCELL_ASAP7_75t_R PHY_599 ();
 OR2x6_ASAP7_75t_R _28096_ (.A(_06935_),
    .B(_09446_),
    .Y(_09454_));
 TAPCELL_ASAP7_75t_R PHY_598 ();
 OAI21x1_ASAP7_75t_R _28098_ (.A1(_06229_),
    .A2(_06927_),
    .B(_06271_),
    .Y(_09456_));
 TAPCELL_ASAP7_75t_R PHY_597 ();
 OA21x2_ASAP7_75t_R _28100_ (.A1(_06229_),
    .A2(_06927_),
    .B(_06271_),
    .Y(_09458_));
 TAPCELL_ASAP7_75t_R PHY_596 ();
 AND2x2_ASAP7_75t_R _28102_ (.A(_01720_),
    .B(_09458_),
    .Y(_09460_));
 AO21x2_ASAP7_75t_R _28103_ (.A1(_00662_),
    .A2(_09456_),
    .B(_09460_),
    .Y(_09461_));
 OAI22x1_ASAP7_75t_R _28104_ (.A1(_00658_),
    .A2(_09454_),
    .B1(_09461_),
    .B2(_06932_),
    .Y(_09462_));
 AO21x1_ASAP7_75t_R _28105_ (.A1(_09446_),
    .A2(net3647),
    .B(_09462_),
    .Y(_02865_));
 NOR2x2_ASAP7_75t_R _28106_ (.A(_06935_),
    .B(_09446_),
    .Y(_09463_));
 TAPCELL_ASAP7_75t_R PHY_595 ();
 TAPCELL_ASAP7_75t_R PHY_594 ();
 TAPCELL_ASAP7_75t_R PHY_593 ();
 AND2x2_ASAP7_75t_R _28110_ (.A(_00162_),
    .B(_09458_),
    .Y(_09467_));
 AO21x2_ASAP7_75t_R _28111_ (.A1(_17754_),
    .A2(_09456_),
    .B(_09467_),
    .Y(_09468_));
 AND3x1_ASAP7_75t_R _28112_ (.A(_02289_),
    .B(_14854_),
    .C(_14923_),
    .Y(_09469_));
 AO21x1_ASAP7_75t_R _28113_ (.A1(_14713_),
    .A2(_18335_),
    .B(_09469_),
    .Y(_09470_));
 AND2x2_ASAP7_75t_R _28114_ (.A(_02286_),
    .B(_09470_),
    .Y(_09471_));
 AO21x1_ASAP7_75t_R _28115_ (.A1(_18336_),
    .A2(net3525),
    .B(_09471_),
    .Y(_09472_));
 AO22x1_ASAP7_75t_R _28116_ (.A1(_06935_),
    .A2(_09468_),
    .B1(net3526),
    .B2(_09446_),
    .Y(_09473_));
 AOI21x1_ASAP7_75t_R _28117_ (.A1(_01575_),
    .A2(_09463_),
    .B(net3527),
    .Y(_02866_));
 NAND2x1_ASAP7_75t_R _28118_ (.A(net306),
    .B(_18339_),
    .Y(_09474_));
 OA21x2_ASAP7_75t_R _28119_ (.A1(_14714_),
    .A2(_18339_),
    .B(_09474_),
    .Y(_09475_));
 INVx2_ASAP7_75t_R _28120_ (.A(_02286_),
    .Y(_09476_));
 OA22x2_ASAP7_75t_R _28121_ (.A1(_18341_),
    .A2(net3562),
    .B1(_09475_),
    .B2(_09476_),
    .Y(_09477_));
 TAPCELL_ASAP7_75t_R PHY_592 ();
 AND2x2_ASAP7_75t_R _28123_ (.A(_00170_),
    .B(_09458_),
    .Y(_09479_));
 AO21x2_ASAP7_75t_R _28124_ (.A1(_01606_),
    .A2(_09456_),
    .B(_09479_),
    .Y(_09480_));
 OAI22x1_ASAP7_75t_R _28125_ (.A1(_00081_),
    .A2(_09454_),
    .B1(_09480_),
    .B2(_06932_),
    .Y(_09481_));
 AO21x1_ASAP7_75t_R _28126_ (.A1(_09446_),
    .A2(net3563),
    .B(_09481_),
    .Y(_02867_));
 TAPCELL_ASAP7_75t_R PHY_591 ();
 NOR2x1_ASAP7_75t_R _28128_ (.A(_14714_),
    .B(_18344_),
    .Y(_09483_));
 AO21x1_ASAP7_75t_R _28129_ (.A1(net306),
    .A2(_18344_),
    .B(_09483_),
    .Y(_09484_));
 AO22x2_ASAP7_75t_R _28130_ (.A1(_18344_),
    .A2(net3385),
    .B1(_09484_),
    .B2(net307),
    .Y(_09485_));
 INVx3_ASAP7_75t_R _28131_ (.A(net3378),
    .Y(_09486_));
 AND2x2_ASAP7_75t_R _28132_ (.A(_00174_),
    .B(_09458_),
    .Y(_09487_));
 AO21x2_ASAP7_75t_R _28133_ (.A1(_01605_),
    .A2(_09456_),
    .B(_09487_),
    .Y(_09488_));
 OAI22x1_ASAP7_75t_R _28134_ (.A1(_00084_),
    .A2(_09454_),
    .B1(_09488_),
    .B2(_06932_),
    .Y(_09489_));
 AO21x1_ASAP7_75t_R _28135_ (.A1(_09446_),
    .A2(net3379),
    .B(_09489_),
    .Y(_02868_));
 AND2x2_ASAP7_75t_R _28136_ (.A(net306),
    .B(_18351_),
    .Y(_09490_));
 AO21x1_ASAP7_75t_R _28137_ (.A1(_14713_),
    .A2(_15115_),
    .B(_09490_),
    .Y(_09491_));
 TAPCELL_ASAP7_75t_R PHY_590 ();
 AOI22x1_ASAP7_75t_R _28139_ (.A1(_18351_),
    .A2(net3631),
    .B1(_09491_),
    .B2(net307),
    .Y(_09493_));
 TAPCELL_ASAP7_75t_R PHY_589 ();
 TAPCELL_ASAP7_75t_R PHY_588 ();
 TAPCELL_ASAP7_75t_R PHY_587 ();
 NAND2x1_ASAP7_75t_R _28143_ (.A(_00177_),
    .B(_09458_),
    .Y(_09497_));
 OA21x2_ASAP7_75t_R _28144_ (.A1(\cs_registers_i.pc_if_i[5] ),
    .A2(_09458_),
    .B(_09497_),
    .Y(_09498_));
 INVx1_ASAP7_75t_R _28145_ (.A(_00087_),
    .Y(_09499_));
 AO32x1_ASAP7_75t_R _28146_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09498_),
    .B1(_09463_),
    .B2(_09499_),
    .Y(_09500_));
 AO21x1_ASAP7_75t_R _28147_ (.A1(_09446_),
    .A2(net3632),
    .B(_09500_),
    .Y(_02869_));
 TAPCELL_ASAP7_75t_R PHY_586 ();
 AND2x2_ASAP7_75t_R _28149_ (.A(_14713_),
    .B(_15172_),
    .Y(_09502_));
 AO21x1_ASAP7_75t_R _28150_ (.A1(_02289_),
    .A2(_18356_),
    .B(_09502_),
    .Y(_09503_));
 AOI22x1_ASAP7_75t_R _28151_ (.A1(_18356_),
    .A2(_07706_),
    .B1(_09503_),
    .B2(_02286_),
    .Y(_09504_));
 NAND2x1_ASAP7_75t_R _28152_ (.A(_01603_),
    .B(_09456_),
    .Y(_09505_));
 OA21x2_ASAP7_75t_R _28153_ (.A1(_15169_),
    .A2(_09456_),
    .B(_09505_),
    .Y(_09506_));
 INVx1_ASAP7_75t_R _28154_ (.A(_00090_),
    .Y(_09507_));
 AO32x1_ASAP7_75t_R _28155_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09506_),
    .B1(_09463_),
    .B2(_09507_),
    .Y(_09508_));
 AO21x1_ASAP7_75t_R _28156_ (.A1(_09446_),
    .A2(_09504_),
    .B(_09508_),
    .Y(_02870_));
 AND2x2_ASAP7_75t_R _28157_ (.A(_14713_),
    .B(_15226_),
    .Y(_09509_));
 AO21x1_ASAP7_75t_R _28158_ (.A1(_02289_),
    .A2(_18361_),
    .B(_09509_),
    .Y(_09510_));
 TAPCELL_ASAP7_75t_R PHY_585 ();
 AOI22x1_ASAP7_75t_R _28160_ (.A1(_18361_),
    .A2(_07748_),
    .B1(_09510_),
    .B2(_02286_),
    .Y(_09512_));
 NAND2x1_ASAP7_75t_R _28161_ (.A(_00182_),
    .B(_09458_),
    .Y(_09513_));
 OA21x2_ASAP7_75t_R _28162_ (.A1(\cs_registers_i.pc_if_i[7] ),
    .A2(_09458_),
    .B(_09513_),
    .Y(_09514_));
 AO32x1_ASAP7_75t_R _28163_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09514_),
    .B1(_09463_),
    .B2(_06367_),
    .Y(_09515_));
 AO21x1_ASAP7_75t_R _28164_ (.A1(_09446_),
    .A2(net3654),
    .B(_09515_),
    .Y(_02871_));
 AND2x2_ASAP7_75t_R _28165_ (.A(_14713_),
    .B(_15280_),
    .Y(_09516_));
 AO21x1_ASAP7_75t_R _28166_ (.A1(net306),
    .A2(_18366_),
    .B(_09516_),
    .Y(_09517_));
 AOI22x1_ASAP7_75t_R _28167_ (.A1(_18366_),
    .A2(_07797_),
    .B1(_09517_),
    .B2(net307),
    .Y(_09518_));
 AND2x2_ASAP7_75t_R _28168_ (.A(_00186_),
    .B(_09458_),
    .Y(_09519_));
 AOI21x1_ASAP7_75t_R _28169_ (.A1(_01601_),
    .A2(_09456_),
    .B(_09519_),
    .Y(_09520_));
 AO32x1_ASAP7_75t_R _28170_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09520_),
    .B1(_09463_),
    .B2(_06382_),
    .Y(_09521_));
 AO21x1_ASAP7_75t_R _28171_ (.A1(_09446_),
    .A2(net3725),
    .B(_09521_),
    .Y(_02872_));
 AND2x2_ASAP7_75t_R _28172_ (.A(_14713_),
    .B(_15337_),
    .Y(_09522_));
 AO21x1_ASAP7_75t_R _28173_ (.A1(net306),
    .A2(_18371_),
    .B(_09522_),
    .Y(_09523_));
 AOI22x1_ASAP7_75t_R _28174_ (.A1(_18371_),
    .A2(_07853_),
    .B1(_09523_),
    .B2(net307),
    .Y(_09524_));
 NAND2x1_ASAP7_75t_R _28175_ (.A(_00189_),
    .B(_09458_),
    .Y(_09525_));
 OA21x2_ASAP7_75t_R _28176_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(_09458_),
    .B(_09525_),
    .Y(_09526_));
 INVx1_ASAP7_75t_R _28177_ (.A(_01572_),
    .Y(_09527_));
 AO32x1_ASAP7_75t_R _28178_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09526_),
    .B1(_09463_),
    .B2(_09527_),
    .Y(_09528_));
 AO21x1_ASAP7_75t_R _28179_ (.A1(_09446_),
    .A2(net3716),
    .B(_09528_),
    .Y(_02873_));
 AND2x2_ASAP7_75t_R _28180_ (.A(_14713_),
    .B(_15401_),
    .Y(_09529_));
 AO21x1_ASAP7_75t_R _28181_ (.A1(net306),
    .A2(_18376_),
    .B(_09529_),
    .Y(_09530_));
 AOI22x1_ASAP7_75t_R _28182_ (.A1(_18376_),
    .A2(_07884_),
    .B1(_09530_),
    .B2(_02286_),
    .Y(_09531_));
 NAND2x1_ASAP7_75t_R _28183_ (.A(_01599_),
    .B(_09456_),
    .Y(_09532_));
 OA21x2_ASAP7_75t_R _28184_ (.A1(_15398_),
    .A2(_09456_),
    .B(_09532_),
    .Y(_09533_));
 INVx1_ASAP7_75t_R _28185_ (.A(_01571_),
    .Y(_09534_));
 AO32x1_ASAP7_75t_R _28186_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09533_),
    .B1(_09463_),
    .B2(_09534_),
    .Y(_09535_));
 AO21x1_ASAP7_75t_R _28187_ (.A1(_09446_),
    .A2(net3736),
    .B(_09535_),
    .Y(_02874_));
 NOR2x1_ASAP7_75t_R _28188_ (.A(_14714_),
    .B(_18379_),
    .Y(_09536_));
 AO21x1_ASAP7_75t_R _28189_ (.A1(net306),
    .A2(_18379_),
    .B(_09536_),
    .Y(_09537_));
 AOI22x1_ASAP7_75t_R _28190_ (.A1(_18379_),
    .A2(_07935_),
    .B1(_09537_),
    .B2(net307),
    .Y(_09538_));
 TAPCELL_ASAP7_75t_R PHY_584 ();
 NAND2x1_ASAP7_75t_R _28192_ (.A(_00196_),
    .B(_09458_),
    .Y(_09540_));
 OA21x2_ASAP7_75t_R _28193_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(_09458_),
    .B(_09540_),
    .Y(_09541_));
 INVx1_ASAP7_75t_R _28194_ (.A(_01570_),
    .Y(_09542_));
 AO32x1_ASAP7_75t_R _28195_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09541_),
    .B1(_09463_),
    .B2(_09542_),
    .Y(_09543_));
 AO21x1_ASAP7_75t_R _28196_ (.A1(_09446_),
    .A2(_09538_),
    .B(_09543_),
    .Y(_02875_));
 TAPCELL_ASAP7_75t_R PHY_583 ();
 INVx1_ASAP7_75t_R _28198_ (.A(net306),
    .Y(_09545_));
 OR2x2_ASAP7_75t_R _28199_ (.A(_18385_),
    .B(_14714_),
    .Y(_09546_));
 OA21x2_ASAP7_75t_R _28200_ (.A1(_09545_),
    .A2(_18383_),
    .B(_09546_),
    .Y(_09547_));
 OA22x2_ASAP7_75t_R _28201_ (.A1(_18383_),
    .A2(_07982_),
    .B1(_09547_),
    .B2(_09476_),
    .Y(_09548_));
 TAPCELL_ASAP7_75t_R PHY_582 ();
 AND2x2_ASAP7_75t_R _28203_ (.A(_00199_),
    .B(_09458_),
    .Y(_09550_));
 AOI21x1_ASAP7_75t_R _28204_ (.A1(_01597_),
    .A2(_09456_),
    .B(_09550_),
    .Y(_09551_));
 INVx1_ASAP7_75t_R _28205_ (.A(_01569_),
    .Y(_09552_));
 AO32x1_ASAP7_75t_R _28206_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09551_),
    .B1(_09463_),
    .B2(_09552_),
    .Y(_09553_));
 AO21x1_ASAP7_75t_R _28207_ (.A1(_09446_),
    .A2(net3673),
    .B(_09553_),
    .Y(_02876_));
 NOR2x1_ASAP7_75t_R _28208_ (.A(_14714_),
    .B(_18390_),
    .Y(_09554_));
 AO21x1_ASAP7_75t_R _28209_ (.A1(net306),
    .A2(_18390_),
    .B(_09554_),
    .Y(_09555_));
 AOI22x1_ASAP7_75t_R _28210_ (.A1(_18390_),
    .A2(_08012_),
    .B1(_09555_),
    .B2(net307),
    .Y(_09556_));
 TAPCELL_ASAP7_75t_R PHY_581 ();
 TAPCELL_ASAP7_75t_R PHY_580 ();
 NAND2x1_ASAP7_75t_R _28213_ (.A(_00201_),
    .B(_09458_),
    .Y(_09559_));
 OA21x2_ASAP7_75t_R _28214_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(_09458_),
    .B(_09559_),
    .Y(_09560_));
 INVx1_ASAP7_75t_R _28215_ (.A(_01568_),
    .Y(_09561_));
 AO32x1_ASAP7_75t_R _28216_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09560_),
    .B1(_09463_),
    .B2(_09561_),
    .Y(_09562_));
 AO21x1_ASAP7_75t_R _28217_ (.A1(_09446_),
    .A2(net3707),
    .B(_09562_),
    .Y(_02877_));
 NAND2x1_ASAP7_75t_R _28218_ (.A(net306),
    .B(_18394_),
    .Y(_09563_));
 OR2x2_ASAP7_75t_R _28219_ (.A(_14714_),
    .B(_18394_),
    .Y(_09564_));
 AO21x1_ASAP7_75t_R _28220_ (.A1(_09563_),
    .A2(_09564_),
    .B(_09476_),
    .Y(_09565_));
 OA21x2_ASAP7_75t_R _28221_ (.A1(_18396_),
    .A2(_08065_),
    .B(_09565_),
    .Y(_09566_));
 TAPCELL_ASAP7_75t_R PHY_579 ();
 NAND2x1_ASAP7_75t_R _28223_ (.A(_01595_),
    .B(_09456_),
    .Y(_09568_));
 OA21x2_ASAP7_75t_R _28224_ (.A1(_15775_),
    .A2(_09456_),
    .B(_09568_),
    .Y(_09569_));
 TAPCELL_ASAP7_75t_R PHY_578 ();
 INVx1_ASAP7_75t_R _28226_ (.A(_01567_),
    .Y(_09571_));
 AO32x1_ASAP7_75t_R _28227_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09569_),
    .B1(_09463_),
    .B2(_09571_),
    .Y(_09572_));
 AO21x1_ASAP7_75t_R _28228_ (.A1(_09446_),
    .A2(net3541),
    .B(_09572_),
    .Y(_02878_));
 AND2x2_ASAP7_75t_R _28229_ (.A(_14713_),
    .B(_15887_),
    .Y(_09573_));
 AO21x1_ASAP7_75t_R _28230_ (.A1(net306),
    .A2(_18400_),
    .B(_09573_),
    .Y(_09574_));
 AOI22x1_ASAP7_75t_R _28231_ (.A1(_18400_),
    .A2(_08106_),
    .B1(_09574_),
    .B2(net307),
    .Y(_09575_));
 TAPCELL_ASAP7_75t_R PHY_577 ();
 TAPCELL_ASAP7_75t_R PHY_576 ();
 TAPCELL_ASAP7_75t_R PHY_575 ();
 NAND2x1_ASAP7_75t_R _28235_ (.A(_00206_),
    .B(_09458_),
    .Y(_09579_));
 OA21x2_ASAP7_75t_R _28236_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(_09458_),
    .B(_09579_),
    .Y(_09580_));
 INVx1_ASAP7_75t_R _28237_ (.A(_01566_),
    .Y(_09581_));
 AO32x1_ASAP7_75t_R _28238_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09580_),
    .B1(_09463_),
    .B2(_09581_),
    .Y(_09582_));
 AO21x1_ASAP7_75t_R _28239_ (.A1(_09446_),
    .A2(net3747),
    .B(_09582_),
    .Y(_02879_));
 AND2x2_ASAP7_75t_R _28240_ (.A(_14713_),
    .B(_16020_),
    .Y(_09583_));
 AO21x1_ASAP7_75t_R _28241_ (.A1(net306),
    .A2(_18404_),
    .B(_09583_),
    .Y(_09584_));
 AOI22x1_ASAP7_75t_R _28242_ (.A1(_18404_),
    .A2(_08142_),
    .B1(_09584_),
    .B2(net307),
    .Y(_09585_));
 AND2x2_ASAP7_75t_R _28243_ (.A(_00208_),
    .B(_09458_),
    .Y(_09586_));
 AOI21x1_ASAP7_75t_R _28244_ (.A1(_01593_),
    .A2(_09456_),
    .B(_09586_),
    .Y(_09587_));
 INVx1_ASAP7_75t_R _28245_ (.A(_01565_),
    .Y(_09588_));
 AO32x1_ASAP7_75t_R _28246_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09587_),
    .B1(_09463_),
    .B2(_09588_),
    .Y(_09589_));
 AO21x1_ASAP7_75t_R _28247_ (.A1(_09446_),
    .A2(net3604),
    .B(_09589_),
    .Y(_02880_));
 AND2x2_ASAP7_75t_R _28248_ (.A(_14713_),
    .B(_16145_),
    .Y(_09590_));
 AO21x1_ASAP7_75t_R _28249_ (.A1(net306),
    .A2(_18409_),
    .B(_09590_),
    .Y(_09591_));
 AOI22x1_ASAP7_75t_R _28250_ (.A1(_18409_),
    .A2(net3667),
    .B1(_09591_),
    .B2(net307),
    .Y(_09592_));
 TAPCELL_ASAP7_75t_R PHY_574 ();
 NAND2x1_ASAP7_75t_R _28252_ (.A(_00209_),
    .B(_09458_),
    .Y(_09594_));
 OA21x2_ASAP7_75t_R _28253_ (.A1(\cs_registers_i.pc_if_i[17] ),
    .A2(_09458_),
    .B(_09594_),
    .Y(_09595_));
 INVx1_ASAP7_75t_R _28254_ (.A(_01564_),
    .Y(_09596_));
 AO32x1_ASAP7_75t_R _28255_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09595_),
    .B1(_09463_),
    .B2(_09596_),
    .Y(_09597_));
 AO21x1_ASAP7_75t_R _28256_ (.A1(_09446_),
    .A2(net3660),
    .B(_09597_),
    .Y(_02881_));
 OR2x2_ASAP7_75t_R _28257_ (.A(_14714_),
    .B(_16262_),
    .Y(_09598_));
 OA21x2_ASAP7_75t_R _28258_ (.A1(_09545_),
    .A2(_18416_),
    .B(_09598_),
    .Y(_09599_));
 OAI22x1_ASAP7_75t_R _28259_ (.A1(_18416_),
    .A2(_08222_),
    .B1(_09599_),
    .B2(_09476_),
    .Y(_09600_));
 INVx3_ASAP7_75t_R _28260_ (.A(net3571),
    .Y(_09601_));
 AND2x2_ASAP7_75t_R _28261_ (.A(_00211_),
    .B(_09458_),
    .Y(_09602_));
 AOI21x1_ASAP7_75t_R _28262_ (.A1(_01591_),
    .A2(_09456_),
    .B(_09602_),
    .Y(_09603_));
 AO32x1_ASAP7_75t_R _28263_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09603_),
    .B1(_09463_),
    .B2(_06465_),
    .Y(_09604_));
 AO21x1_ASAP7_75t_R _28264_ (.A1(_09446_),
    .A2(net3557),
    .B(_09604_),
    .Y(_02882_));
 NOR2x1_ASAP7_75t_R _28265_ (.A(_14714_),
    .B(_16386_),
    .Y(_09605_));
 AO21x1_ASAP7_75t_R _28266_ (.A1(net306),
    .A2(_16386_),
    .B(_09605_),
    .Y(_09606_));
 AOI22x1_ASAP7_75t_R _28267_ (.A1(_16386_),
    .A2(net3720),
    .B1(_09606_),
    .B2(net307),
    .Y(_09607_));
 TAPCELL_ASAP7_75t_R PHY_573 ();
 NAND2x1_ASAP7_75t_R _28269_ (.A(_00212_),
    .B(_09458_),
    .Y(_09609_));
 OA21x2_ASAP7_75t_R _28270_ (.A1(\cs_registers_i.pc_if_i[19] ),
    .A2(_09458_),
    .B(_09609_),
    .Y(_09610_));
 INVx1_ASAP7_75t_R _28271_ (.A(_01562_),
    .Y(_09611_));
 AO32x1_ASAP7_75t_R _28272_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09610_),
    .B1(_09463_),
    .B2(_09611_),
    .Y(_09612_));
 AO21x1_ASAP7_75t_R _28273_ (.A1(_09446_),
    .A2(net3711),
    .B(_09612_),
    .Y(_02883_));
 NOR2x1_ASAP7_75t_R _28274_ (.A(_14714_),
    .B(_18424_),
    .Y(_09613_));
 AO21x1_ASAP7_75t_R _28275_ (.A1(net306),
    .A2(_18424_),
    .B(_09613_),
    .Y(_09614_));
 AO22x2_ASAP7_75t_R _28276_ (.A1(_18424_),
    .A2(net3681),
    .B1(_09614_),
    .B2(net307),
    .Y(_09615_));
 INVx4_ASAP7_75t_R _28277_ (.A(net3682),
    .Y(_09616_));
 AND2x2_ASAP7_75t_R _28278_ (.A(_00214_),
    .B(_09458_),
    .Y(_09617_));
 AOI21x1_ASAP7_75t_R _28279_ (.A1(_01589_),
    .A2(_09456_),
    .B(_09617_),
    .Y(_09618_));
 INVx1_ASAP7_75t_R _28280_ (.A(_01561_),
    .Y(_09619_));
 AO32x1_ASAP7_75t_R _28281_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09618_),
    .B1(_09463_),
    .B2(_09619_),
    .Y(_09620_));
 AO21x1_ASAP7_75t_R _28282_ (.A1(_09446_),
    .A2(net3683),
    .B(_09620_),
    .Y(_02884_));
 AND2x2_ASAP7_75t_R _28283_ (.A(_14713_),
    .B(_16620_),
    .Y(_09621_));
 AO21x1_ASAP7_75t_R _28284_ (.A1(net306),
    .A2(_18429_),
    .B(_09621_),
    .Y(_09622_));
 AOI22x1_ASAP7_75t_R _28285_ (.A1(_18429_),
    .A2(net3677),
    .B1(_09622_),
    .B2(_02286_),
    .Y(_09623_));
 TAPCELL_ASAP7_75t_R PHY_572 ();
 NAND2x1_ASAP7_75t_R _28287_ (.A(_00215_),
    .B(_09458_),
    .Y(_09625_));
 OA21x2_ASAP7_75t_R _28288_ (.A1(\cs_registers_i.pc_if_i[21] ),
    .A2(_09458_),
    .B(_09625_),
    .Y(_09626_));
 AO32x1_ASAP7_75t_R _28289_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09626_),
    .B1(_09463_),
    .B2(_06485_),
    .Y(_09627_));
 AO21x1_ASAP7_75t_R _28290_ (.A1(_09446_),
    .A2(net3678),
    .B(_09627_),
    .Y(_02885_));
 TAPCELL_ASAP7_75t_R PHY_571 ();
 AND2x2_ASAP7_75t_R _28292_ (.A(_14713_),
    .B(_04516_),
    .Y(_09629_));
 AO21x1_ASAP7_75t_R _28293_ (.A1(net306),
    .A2(_18435_),
    .B(_09629_),
    .Y(_09630_));
 AOI22x1_ASAP7_75t_R _28294_ (.A1(_18435_),
    .A2(net3690),
    .B1(_09630_),
    .B2(net307),
    .Y(_09631_));
 AND2x2_ASAP7_75t_R _28295_ (.A(_00217_),
    .B(_09458_),
    .Y(_09632_));
 AOI21x1_ASAP7_75t_R _28296_ (.A1(_01587_),
    .A2(_09456_),
    .B(_09632_),
    .Y(_09633_));
 AO32x1_ASAP7_75t_R _28297_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09633_),
    .B1(_09463_),
    .B2(_06492_),
    .Y(_09634_));
 AO21x1_ASAP7_75t_R _28298_ (.A1(_09446_),
    .A2(net3691),
    .B(_09634_),
    .Y(_02886_));
 AND2x2_ASAP7_75t_R _28299_ (.A(_14713_),
    .B(_04632_),
    .Y(_09635_));
 AO21x1_ASAP7_75t_R _28300_ (.A1(net306),
    .A2(_18440_),
    .B(_09635_),
    .Y(_09636_));
 AO22x2_ASAP7_75t_R _28301_ (.A1(_18440_),
    .A2(_08399_),
    .B1(_09636_),
    .B2(_02286_),
    .Y(_09637_));
 INVx5_ASAP7_75t_R _28302_ (.A(net3599),
    .Y(_09638_));
 NAND2x1_ASAP7_75t_R _28303_ (.A(_00218_),
    .B(_09458_),
    .Y(_09639_));
 OA21x2_ASAP7_75t_R _28304_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(_09458_),
    .B(_09639_),
    .Y(_09640_));
 INVx1_ASAP7_75t_R _28305_ (.A(_01558_),
    .Y(_09641_));
 AO32x1_ASAP7_75t_R _28306_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09640_),
    .B1(_09463_),
    .B2(_09641_),
    .Y(_09642_));
 AO21x1_ASAP7_75t_R _28307_ (.A1(_09446_),
    .A2(_09638_),
    .B(_09642_),
    .Y(_02887_));
 NOR2x2_ASAP7_75t_R _28308_ (.A(_18446_),
    .B(_08445_),
    .Y(_09643_));
 NOR2x1_ASAP7_75t_R _28309_ (.A(_14714_),
    .B(_18444_),
    .Y(_09644_));
 AO21x1_ASAP7_75t_R _28310_ (.A1(net306),
    .A2(_18444_),
    .B(_09644_),
    .Y(_09645_));
 AND2x4_ASAP7_75t_R _28311_ (.A(_02286_),
    .B(_09645_),
    .Y(_09646_));
 NOR2x2_ASAP7_75t_R _28312_ (.A(net3531),
    .B(_09646_),
    .Y(_09647_));
 AND2x2_ASAP7_75t_R _28313_ (.A(_00220_),
    .B(_09458_),
    .Y(_09648_));
 AO21x2_ASAP7_75t_R _28314_ (.A1(_01585_),
    .A2(_09456_),
    .B(_09648_),
    .Y(_09649_));
 OAI22x1_ASAP7_75t_R _28315_ (.A1(_01557_),
    .A2(_09454_),
    .B1(_09649_),
    .B2(_06932_),
    .Y(_09650_));
 AO21x1_ASAP7_75t_R _28316_ (.A1(_09446_),
    .A2(_09647_),
    .B(_09650_),
    .Y(_02888_));
 AND2x2_ASAP7_75t_R _28317_ (.A(_14713_),
    .B(_04857_),
    .Y(_09651_));
 AO21x1_ASAP7_75t_R _28318_ (.A1(net306),
    .A2(_18449_),
    .B(_09651_),
    .Y(_09652_));
 AOI22x1_ASAP7_75t_R _28319_ (.A1(_18449_),
    .A2(_08478_),
    .B1(_09652_),
    .B2(_02286_),
    .Y(_09653_));
 TAPCELL_ASAP7_75t_R PHY_570 ();
 NAND2x1_ASAP7_75t_R _28321_ (.A(_00221_),
    .B(_09458_),
    .Y(_09655_));
 OA21x2_ASAP7_75t_R _28322_ (.A1(\cs_registers_i.pc_if_i[25] ),
    .A2(_09458_),
    .B(_09655_),
    .Y(_09656_));
 INVx1_ASAP7_75t_R _28323_ (.A(_01556_),
    .Y(_09657_));
 AO32x1_ASAP7_75t_R _28324_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09656_),
    .B1(_09463_),
    .B2(_09657_),
    .Y(_09658_));
 AO21x1_ASAP7_75t_R _28325_ (.A1(_09446_),
    .A2(net3644),
    .B(_09658_),
    .Y(_02889_));
 AND2x2_ASAP7_75t_R _28326_ (.A(_14713_),
    .B(_04967_),
    .Y(_09659_));
 AO21x1_ASAP7_75t_R _28327_ (.A1(net306),
    .A2(_18455_),
    .B(_09659_),
    .Y(_09660_));
 AO22x2_ASAP7_75t_R _28328_ (.A1(_18455_),
    .A2(net3752),
    .B1(_09660_),
    .B2(_02286_),
    .Y(_09661_));
 INVx4_ASAP7_75t_R _28329_ (.A(_09661_),
    .Y(_09662_));
 AND2x2_ASAP7_75t_R _28330_ (.A(_00223_),
    .B(_09458_),
    .Y(_09663_));
 AOI21x1_ASAP7_75t_R _28331_ (.A1(_01583_),
    .A2(_09456_),
    .B(_09663_),
    .Y(_09664_));
 AO32x1_ASAP7_75t_R _28332_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09664_),
    .B1(_09463_),
    .B2(_06520_),
    .Y(_09665_));
 AO21x1_ASAP7_75t_R _28333_ (.A1(_09446_),
    .A2(_09662_),
    .B(_09665_),
    .Y(_02890_));
 AND2x2_ASAP7_75t_R _28334_ (.A(_14713_),
    .B(_05077_),
    .Y(_09666_));
 AO21x1_ASAP7_75t_R _28335_ (.A1(net306),
    .A2(_18460_),
    .B(_09666_),
    .Y(_09667_));
 AOI22x1_ASAP7_75t_R _28336_ (.A1(_18460_),
    .A2(_08535_),
    .B1(_09667_),
    .B2(net307),
    .Y(_09668_));
 TAPCELL_ASAP7_75t_R PHY_569 ();
 NAND2x1_ASAP7_75t_R _28338_ (.A(_00224_),
    .B(_09458_),
    .Y(_09670_));
 OA21x2_ASAP7_75t_R _28339_ (.A1(\cs_registers_i.pc_if_i[27] ),
    .A2(_09458_),
    .B(_09670_),
    .Y(_09671_));
 INVx1_ASAP7_75t_R _28340_ (.A(_01554_),
    .Y(_09672_));
 AO32x1_ASAP7_75t_R _28341_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09671_),
    .B1(_09463_),
    .B2(_09672_),
    .Y(_09673_));
 AO21x1_ASAP7_75t_R _28342_ (.A1(_09446_),
    .A2(net3594),
    .B(_09673_),
    .Y(_02891_));
 NOR2x1_ASAP7_75t_R _28343_ (.A(_14714_),
    .B(_05184_),
    .Y(_09674_));
 AO21x1_ASAP7_75t_R _28344_ (.A1(net306),
    .A2(_05184_),
    .B(_09674_),
    .Y(_09675_));
 AOI22x1_ASAP7_75t_R _28345_ (.A1(_05184_),
    .A2(net3742),
    .B1(_09675_),
    .B2(net307),
    .Y(_09676_));
 AND2x2_ASAP7_75t_R _28346_ (.A(_00226_),
    .B(_09458_),
    .Y(_09677_));
 AOI21x1_ASAP7_75t_R _28347_ (.A1(_01581_),
    .A2(_09456_),
    .B(_09677_),
    .Y(_09678_));
 INVx1_ASAP7_75t_R _28348_ (.A(_01553_),
    .Y(_09679_));
 AO32x1_ASAP7_75t_R _28349_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09678_),
    .B1(_09463_),
    .B2(_09679_),
    .Y(_09680_));
 AO21x1_ASAP7_75t_R _28350_ (.A1(_09446_),
    .A2(_09676_),
    .B(_09680_),
    .Y(_02892_));
 AND3x1_ASAP7_75t_R _28351_ (.A(_02289_),
    .B(_05292_),
    .C(_05294_),
    .Y(_09681_));
 AO21x1_ASAP7_75t_R _28352_ (.A1(_14713_),
    .A2(_18471_),
    .B(_09681_),
    .Y(_09682_));
 AOI22x1_ASAP7_75t_R _28353_ (.A1(_18469_),
    .A2(net3610),
    .B1(_09682_),
    .B2(_02286_),
    .Y(_09683_));
 TAPCELL_ASAP7_75t_R PHY_568 ();
 NAND2x1_ASAP7_75t_R _28355_ (.A(_00227_),
    .B(_09458_),
    .Y(_09685_));
 OA21x2_ASAP7_75t_R _28356_ (.A1(\cs_registers_i.pc_if_i[29] ),
    .A2(_09458_),
    .B(_09685_),
    .Y(_09686_));
 INVx1_ASAP7_75t_R _28357_ (.A(_01552_),
    .Y(_09687_));
 AO32x1_ASAP7_75t_R _28358_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09686_),
    .B1(_09463_),
    .B2(_09687_),
    .Y(_09688_));
 AO21x1_ASAP7_75t_R _28359_ (.A1(_09446_),
    .A2(net3611),
    .B(_09688_),
    .Y(_02893_));
 OR2x2_ASAP7_75t_R _28360_ (.A(_14714_),
    .B(_18474_),
    .Y(_09689_));
 OA21x2_ASAP7_75t_R _28361_ (.A1(_09545_),
    .A2(_18476_),
    .B(_09689_),
    .Y(_09690_));
 OA22x2_ASAP7_75t_R _28362_ (.A1(_18476_),
    .A2(net3697),
    .B1(_09690_),
    .B2(_09476_),
    .Y(_09691_));
 TAPCELL_ASAP7_75t_R PHY_567 ();
 NAND2x1_ASAP7_75t_R _28364_ (.A(_01579_),
    .B(_09456_),
    .Y(_09693_));
 OA21x2_ASAP7_75t_R _28365_ (.A1(_05401_),
    .A2(_09456_),
    .B(_09693_),
    .Y(_09694_));
 AO32x1_ASAP7_75t_R _28366_ (.A1(_06230_),
    .A2(_06931_),
    .A3(_09694_),
    .B1(_09463_),
    .B2(_06547_),
    .Y(_09695_));
 AO21x1_ASAP7_75t_R _28367_ (.A1(_09446_),
    .A2(net3698),
    .B(_09695_),
    .Y(_02894_));
 AND3x1_ASAP7_75t_R _28368_ (.A(_14713_),
    .B(_05457_),
    .C(_05511_),
    .Y(_09696_));
 AO21x1_ASAP7_75t_R _28369_ (.A1(_02289_),
    .A2(_17805_),
    .B(_09696_),
    .Y(_09697_));
 AOI22x1_ASAP7_75t_R _28370_ (.A1(_17805_),
    .A2(_08633_),
    .B1(_09697_),
    .B2(_02286_),
    .Y(_09698_));
 TAPCELL_ASAP7_75t_R PHY_566 ();
 AND2x2_ASAP7_75t_R _28372_ (.A(_00230_),
    .B(_09458_),
    .Y(_09700_));
 AO21x1_ASAP7_75t_R _28373_ (.A1(_01578_),
    .A2(_09456_),
    .B(_09700_),
    .Y(_09701_));
 OAI22x1_ASAP7_75t_R _28374_ (.A1(_01550_),
    .A2(_09454_),
    .B1(_09701_),
    .B2(_06932_),
    .Y(_09702_));
 AO21x1_ASAP7_75t_R _28375_ (.A1(_09446_),
    .A2(_09698_),
    .B(_09702_),
    .Y(_02895_));
 NAND2x2_ASAP7_75t_R _28376_ (.A(net301),
    .B(_06834_),
    .Y(_09703_));
 TAPCELL_ASAP7_75t_R PHY_565 ();
 AND3x1_ASAP7_75t_R _28378_ (.A(_01549_),
    .B(net300),
    .C(_06834_),
    .Y(_09705_));
 AOI21x1_ASAP7_75t_R _28379_ (.A1(_02596_),
    .A2(_09703_),
    .B(_09705_),
    .Y(_02896_));
 AND3x1_ASAP7_75t_R _28380_ (.A(_01548_),
    .B(net300),
    .C(_06834_),
    .Y(_09706_));
 AOI21x1_ASAP7_75t_R _28381_ (.A1(_02567_),
    .A2(_09703_),
    .B(_09706_),
    .Y(_02897_));
 AND3x1_ASAP7_75t_R _28382_ (.A(_01547_),
    .B(net300),
    .C(_06834_),
    .Y(_09707_));
 AOI21x1_ASAP7_75t_R _28383_ (.A1(_02569_),
    .A2(_09703_),
    .B(_09707_),
    .Y(_02898_));
 AND2x6_ASAP7_75t_R _28384_ (.A(net301),
    .B(_06834_),
    .Y(_09708_));
 TAPCELL_ASAP7_75t_R PHY_564 ();
 XOR2x1_ASAP7_75t_R _28386_ (.A(_02568_),
    .Y(_09710_),
    .B(_06353_));
 NAND2x1_ASAP7_75t_R _28387_ (.A(_01546_),
    .B(_09708_),
    .Y(_09711_));
 OA21x2_ASAP7_75t_R _28388_ (.A1(_09708_),
    .A2(_09710_),
    .B(_09711_),
    .Y(_02899_));
 AND3x1_ASAP7_75t_R _28389_ (.A(_01545_),
    .B(net300),
    .C(_06834_),
    .Y(_09712_));
 AOI21x1_ASAP7_75t_R _28390_ (.A1(_02571_),
    .A2(_09703_),
    .B(_09712_),
    .Y(_02900_));
 TAPCELL_ASAP7_75t_R PHY_563 ();
 XOR2x1_ASAP7_75t_R _28392_ (.A(_02570_),
    .Y(_09714_),
    .B(_06378_));
 NOR2x1_ASAP7_75t_R _28393_ (.A(_01544_),
    .B(_09703_),
    .Y(_09715_));
 AO21x1_ASAP7_75t_R _28394_ (.A1(_09703_),
    .A2(_09714_),
    .B(_09715_),
    .Y(_02901_));
 AND3x1_ASAP7_75t_R _28395_ (.A(_01543_),
    .B(net301),
    .C(_06834_),
    .Y(_09716_));
 AOI21x1_ASAP7_75t_R _28396_ (.A1(_02573_),
    .A2(_09703_),
    .B(_09716_),
    .Y(_02902_));
 XOR2x1_ASAP7_75t_R _28397_ (.A(_02572_),
    .Y(_09717_),
    .B(_06397_));
 NAND2x1_ASAP7_75t_R _28398_ (.A(_01542_),
    .B(_09708_),
    .Y(_09718_));
 OA21x2_ASAP7_75t_R _28399_ (.A1(_09708_),
    .A2(_09717_),
    .B(_09718_),
    .Y(_02903_));
 AND3x1_ASAP7_75t_R _28400_ (.A(_01541_),
    .B(net301),
    .C(_06834_),
    .Y(_09719_));
 AOI21x1_ASAP7_75t_R _28401_ (.A1(_02575_),
    .A2(_09703_),
    .B(_09719_),
    .Y(_02904_));
 XOR2x1_ASAP7_75t_R _28402_ (.A(_02574_),
    .Y(_09720_),
    .B(_06417_));
 NAND2x1_ASAP7_75t_R _28403_ (.A(_01540_),
    .B(_09708_),
    .Y(_09721_));
 OA21x2_ASAP7_75t_R _28404_ (.A1(_09708_),
    .A2(_09720_),
    .B(_09721_),
    .Y(_02905_));
 TAPCELL_ASAP7_75t_R PHY_562 ();
 AND3x1_ASAP7_75t_R _28406_ (.A(_01539_),
    .B(net301),
    .C(_06834_),
    .Y(_09723_));
 AOI21x1_ASAP7_75t_R _28407_ (.A1(_02577_),
    .A2(_09703_),
    .B(_09723_),
    .Y(_02906_));
 OR3x1_ASAP7_75t_R _28408_ (.A(_06354_),
    .B(_02576_),
    .C(_06565_),
    .Y(_09724_));
 XOR2x1_ASAP7_75t_R _28409_ (.A(_01538_),
    .Y(_09725_),
    .B(_09724_));
 XOR2x1_ASAP7_75t_R _28410_ (.A(_02576_),
    .Y(_09726_),
    .B(_06432_));
 AND2x2_ASAP7_75t_R _28411_ (.A(net299),
    .B(_09726_),
    .Y(_09727_));
 AO21x1_ASAP7_75t_R _28412_ (.A1(net300),
    .A2(_09725_),
    .B(_09727_),
    .Y(_02907_));
 AND3x1_ASAP7_75t_R _28413_ (.A(_01537_),
    .B(net301),
    .C(_06834_),
    .Y(_09728_));
 AOI21x1_ASAP7_75t_R _28414_ (.A1(_02579_),
    .A2(_09703_),
    .B(_09728_),
    .Y(_02908_));
 XOR2x1_ASAP7_75t_R _28415_ (.A(_02578_),
    .Y(_09729_),
    .B(_06447_));
 NOR2x1_ASAP7_75t_R _28416_ (.A(_01536_),
    .B(_09703_),
    .Y(_09730_));
 AO21x1_ASAP7_75t_R _28417_ (.A1(_09703_),
    .A2(_09729_),
    .B(_09730_),
    .Y(_02909_));
 AND3x1_ASAP7_75t_R _28418_ (.A(_01535_),
    .B(net301),
    .C(_06834_),
    .Y(_09731_));
 AOI21x1_ASAP7_75t_R _28419_ (.A1(_02581_),
    .A2(_09703_),
    .B(_09731_),
    .Y(_02910_));
 XOR2x1_ASAP7_75t_R _28420_ (.A(_02580_),
    .Y(_09732_),
    .B(_06463_));
 NOR2x1_ASAP7_75t_R _28421_ (.A(_01534_),
    .B(_09703_),
    .Y(_09733_));
 AO21x1_ASAP7_75t_R _28422_ (.A1(_09703_),
    .A2(_09732_),
    .B(_09733_),
    .Y(_02911_));
 AND3x1_ASAP7_75t_R _28423_ (.A(_01533_),
    .B(net301),
    .C(_06834_),
    .Y(_09734_));
 AOI21x1_ASAP7_75t_R _28424_ (.A1(_02583_),
    .A2(_09703_),
    .B(_09734_),
    .Y(_02912_));
 XNOR2x1_ASAP7_75t_R _28425_ (.B(_06476_),
    .Y(_09735_),
    .A(_02582_));
 NOR2x1_ASAP7_75t_R _28426_ (.A(_01532_),
    .B(_09703_),
    .Y(_09736_));
 AO21x1_ASAP7_75t_R _28427_ (.A1(_09703_),
    .A2(_09735_),
    .B(_09736_),
    .Y(_02913_));
 AND3x1_ASAP7_75t_R _28428_ (.A(_01531_),
    .B(net301),
    .C(_06834_),
    .Y(_09737_));
 AOI21x1_ASAP7_75t_R _28429_ (.A1(_02585_),
    .A2(_09703_),
    .B(_09737_),
    .Y(_02914_));
 XNOR2x1_ASAP7_75t_R _28430_ (.B(_06490_),
    .Y(_09738_),
    .A(_02584_));
 NOR2x1_ASAP7_75t_R _28431_ (.A(_01530_),
    .B(_09703_),
    .Y(_09739_));
 AO21x1_ASAP7_75t_R _28432_ (.A1(_09703_),
    .A2(_09738_),
    .B(_09739_),
    .Y(_02915_));
 AND3x1_ASAP7_75t_R _28433_ (.A(_01529_),
    .B(net301),
    .C(_06834_),
    .Y(_09740_));
 AOI21x1_ASAP7_75t_R _28434_ (.A1(_02587_),
    .A2(_09703_),
    .B(_09740_),
    .Y(_02916_));
 XNOR2x1_ASAP7_75t_R _28435_ (.B(_06503_),
    .Y(_09741_),
    .A(_02586_));
 NAND2x1_ASAP7_75t_R _28436_ (.A(_01528_),
    .B(_09708_),
    .Y(_09742_));
 OA21x2_ASAP7_75t_R _28437_ (.A1(_09708_),
    .A2(_09741_),
    .B(_09742_),
    .Y(_02917_));
 AND3x1_ASAP7_75t_R _28438_ (.A(_01527_),
    .B(net301),
    .C(_06834_),
    .Y(_09743_));
 AOI21x1_ASAP7_75t_R _28439_ (.A1(_02589_),
    .A2(_09703_),
    .B(_09743_),
    .Y(_02918_));
 XNOR2x1_ASAP7_75t_R _28440_ (.B(_06517_),
    .Y(_09744_),
    .A(_02588_));
 NAND2x1_ASAP7_75t_R _28441_ (.A(_01526_),
    .B(_09708_),
    .Y(_09745_));
 OA21x2_ASAP7_75t_R _28442_ (.A1(_09708_),
    .A2(_09744_),
    .B(_09745_),
    .Y(_02919_));
 AND3x1_ASAP7_75t_R _28443_ (.A(_01525_),
    .B(net301),
    .C(_06834_),
    .Y(_09746_));
 AOI21x1_ASAP7_75t_R _28444_ (.A1(_02591_),
    .A2(_09703_),
    .B(_09746_),
    .Y(_02920_));
 XNOR2x1_ASAP7_75t_R _28445_ (.B(_06532_),
    .Y(_09747_),
    .A(_02590_));
 NAND2x1_ASAP7_75t_R _28446_ (.A(_01524_),
    .B(_09708_),
    .Y(_09748_));
 OA21x2_ASAP7_75t_R _28447_ (.A1(_09708_),
    .A2(_09747_),
    .B(_09748_),
    .Y(_02921_));
 AND3x1_ASAP7_75t_R _28448_ (.A(_01523_),
    .B(net301),
    .C(_06834_),
    .Y(_09749_));
 AOI21x1_ASAP7_75t_R _28449_ (.A1(_02593_),
    .A2(_09703_),
    .B(_09749_),
    .Y(_02922_));
 XNOR2x1_ASAP7_75t_R _28450_ (.B(_06545_),
    .Y(_09750_),
    .A(_02592_));
 NAND2x1_ASAP7_75t_R _28451_ (.A(_01522_),
    .B(_09708_),
    .Y(_09751_));
 OA21x2_ASAP7_75t_R _28452_ (.A1(_09708_),
    .A2(_09750_),
    .B(_09751_),
    .Y(_02923_));
 AND3x1_ASAP7_75t_R _28453_ (.A(_01521_),
    .B(net301),
    .C(_06834_),
    .Y(_09752_));
 AOI21x1_ASAP7_75t_R _28454_ (.A1(_02595_),
    .A2(_09703_),
    .B(_09752_),
    .Y(_02924_));
 XNOR2x1_ASAP7_75t_R _28455_ (.B(_06557_),
    .Y(_09753_),
    .A(_02594_));
 NOR2x1_ASAP7_75t_R _28456_ (.A(_01520_),
    .B(_09703_),
    .Y(_09754_));
 AO21x1_ASAP7_75t_R _28457_ (.A1(_09703_),
    .A2(_09753_),
    .B(_09754_),
    .Y(_02925_));
 OR2x2_ASAP7_75t_R _28458_ (.A(_06981_),
    .B(_06983_),
    .Y(_09755_));
 AND4x2_ASAP7_75t_R _28459_ (.A(_00323_),
    .B(_05658_),
    .C(_00194_),
    .D(_09755_),
    .Y(_09756_));
 NAND2x2_ASAP7_75t_R _28460_ (.A(_14834_),
    .B(_09756_),
    .Y(_09757_));
 TAPCELL_ASAP7_75t_R PHY_561 ();
 TAPCELL_ASAP7_75t_R PHY_560 ();
 NOR2x1_ASAP7_75t_R _28463_ (.A(_07248_),
    .B(_09757_),
    .Y(_09760_));
 AO21x1_ASAP7_75t_R _28464_ (.A1(_13847_),
    .A2(_09757_),
    .B(_09760_),
    .Y(_02926_));
 TAPCELL_ASAP7_75t_R PHY_559 ();
 AND2x6_ASAP7_75t_R _28466_ (.A(_14834_),
    .B(_09756_),
    .Y(_09762_));
 TAPCELL_ASAP7_75t_R PHY_558 ();
 TAPCELL_ASAP7_75t_R PHY_557 ();
 AND2x2_ASAP7_75t_R _28469_ (.A(_13412_),
    .B(_09757_),
    .Y(_09765_));
 AO21x1_ASAP7_75t_R _28470_ (.A1(_07384_),
    .A2(_09762_),
    .B(_09765_),
    .Y(_02927_));
 TAPCELL_ASAP7_75t_R PHY_556 ();
 AND2x2_ASAP7_75t_R _28472_ (.A(_14165_),
    .B(_09757_),
    .Y(_09767_));
 AO21x1_ASAP7_75t_R _28473_ (.A1(_07472_),
    .A2(_09762_),
    .B(_09767_),
    .Y(_02928_));
 TAPCELL_ASAP7_75t_R PHY_555 ();
 TAPCELL_ASAP7_75t_R PHY_554 ();
 NOR2x1_ASAP7_75t_R _28476_ (.A(_00386_),
    .B(_09762_),
    .Y(_09770_));
 AO21x1_ASAP7_75t_R _28477_ (.A1(_07552_),
    .A2(_09762_),
    .B(_09770_),
    .Y(_02929_));
 TAPCELL_ASAP7_75t_R PHY_553 ();
 AND2x2_ASAP7_75t_R _28479_ (.A(_14258_),
    .B(_09757_),
    .Y(_09772_));
 AO21x1_ASAP7_75t_R _28480_ (.A1(_07608_),
    .A2(_09762_),
    .B(_09772_),
    .Y(_02930_));
 TAPCELL_ASAP7_75t_R PHY_552 ();
 AND2x2_ASAP7_75t_R _28482_ (.A(_14349_),
    .B(_09757_),
    .Y(_09774_));
 AO21x1_ASAP7_75t_R _28483_ (.A1(_07663_),
    .A2(_09762_),
    .B(_09774_),
    .Y(_02931_));
 TAPCELL_ASAP7_75t_R PHY_551 ();
 AND2x2_ASAP7_75t_R _28485_ (.A(_14388_),
    .B(_09757_),
    .Y(_09776_));
 AO21x1_ASAP7_75t_R _28486_ (.A1(_07709_),
    .A2(_09762_),
    .B(_09776_),
    .Y(_02932_));
 TAPCELL_ASAP7_75t_R PHY_550 ();
 AND2x2_ASAP7_75t_R _28488_ (.A(_14446_),
    .B(_09757_),
    .Y(_09778_));
 AO21x1_ASAP7_75t_R _28489_ (.A1(net252),
    .A2(_09762_),
    .B(_09778_),
    .Y(_02933_));
 TAPCELL_ASAP7_75t_R PHY_549 ();
 AND2x2_ASAP7_75t_R _28491_ (.A(_14504_),
    .B(_09757_),
    .Y(_09780_));
 AO21x1_ASAP7_75t_R _28492_ (.A1(net257),
    .A2(_09762_),
    .B(_09780_),
    .Y(_02934_));
 TAPCELL_ASAP7_75t_R PHY_548 ();
 AND2x2_ASAP7_75t_R _28494_ (.A(_14568_),
    .B(_09757_),
    .Y(_09782_));
 AO21x1_ASAP7_75t_R _28495_ (.A1(net256),
    .A2(_09762_),
    .B(_09782_),
    .Y(_02935_));
 TAPCELL_ASAP7_75t_R PHY_547 ();
 NOR2x1_ASAP7_75t_R _28497_ (.A(_00596_),
    .B(_09762_),
    .Y(_09784_));
 AO21x1_ASAP7_75t_R _28498_ (.A1(_07903_),
    .A2(_09762_),
    .B(_09784_),
    .Y(_02936_));
 TAPCELL_ASAP7_75t_R PHY_546 ();
 TAPCELL_ASAP7_75t_R PHY_545 ();
 AND2x2_ASAP7_75t_R _28501_ (.A(_14672_),
    .B(_09757_),
    .Y(_09787_));
 AO21x1_ASAP7_75t_R _28502_ (.A1(_07948_),
    .A2(_09762_),
    .B(_09787_),
    .Y(_02937_));
 TAPCELL_ASAP7_75t_R PHY_544 ();
 NOR2x1_ASAP7_75t_R _28504_ (.A(_00325_),
    .B(_09762_),
    .Y(_09789_));
 AO21x1_ASAP7_75t_R _28505_ (.A1(_07985_),
    .A2(_09762_),
    .B(_09789_),
    .Y(_02938_));
 TAPCELL_ASAP7_75t_R PHY_543 ();
 NOR2x1_ASAP7_75t_R _28507_ (.A(_00688_),
    .B(_09762_),
    .Y(_09791_));
 AO21x1_ASAP7_75t_R _28508_ (.A1(net251),
    .A2(_09762_),
    .B(_09791_),
    .Y(_02939_));
 TAPCELL_ASAP7_75t_R PHY_542 ();
 NOR2x1_ASAP7_75t_R _28510_ (.A(_00720_),
    .B(_09762_),
    .Y(_09793_));
 AO21x1_ASAP7_75t_R _28511_ (.A1(_08068_),
    .A2(_09762_),
    .B(_09793_),
    .Y(_02940_));
 TAPCELL_ASAP7_75t_R PHY_541 ();
 NOR2x1_ASAP7_75t_R _28513_ (.A(_00753_),
    .B(_09762_),
    .Y(_09795_));
 AO21x1_ASAP7_75t_R _28514_ (.A1(_08110_),
    .A2(_09762_),
    .B(_09795_),
    .Y(_02941_));
 TAPCELL_ASAP7_75t_R PHY_540 ();
 NOR2x1_ASAP7_75t_R _28516_ (.A(_00786_),
    .B(_09762_),
    .Y(_09797_));
 AO21x1_ASAP7_75t_R _28517_ (.A1(_08151_),
    .A2(_09762_),
    .B(_09797_),
    .Y(_02942_));
 TAPCELL_ASAP7_75t_R PHY_539 ();
 NOR2x1_ASAP7_75t_R _28519_ (.A(_00819_),
    .B(_09762_),
    .Y(_09799_));
 AO21x1_ASAP7_75t_R _28520_ (.A1(_08190_),
    .A2(_09762_),
    .B(_09799_),
    .Y(_02943_));
 TAPCELL_ASAP7_75t_R PHY_538 ();
 NOR2x1_ASAP7_75t_R _28522_ (.A(_00851_),
    .B(_09762_),
    .Y(_09801_));
 AO21x1_ASAP7_75t_R _28523_ (.A1(_08225_),
    .A2(_09762_),
    .B(_09801_),
    .Y(_02944_));
 TAPCELL_ASAP7_75t_R PHY_537 ();
 NOR2x1_ASAP7_75t_R _28525_ (.A(_00884_),
    .B(_09762_),
    .Y(_09803_));
 AO21x1_ASAP7_75t_R _28526_ (.A1(_08263_),
    .A2(_09762_),
    .B(_09803_),
    .Y(_02945_));
 TAPCELL_ASAP7_75t_R PHY_536 ();
 AND2x2_ASAP7_75t_R _28528_ (.A(_16393_),
    .B(_09757_),
    .Y(_09805_));
 AO21x1_ASAP7_75t_R _28529_ (.A1(_08294_),
    .A2(_09762_),
    .B(_09805_),
    .Y(_02946_));
 TAPCELL_ASAP7_75t_R PHY_535 ();
 TAPCELL_ASAP7_75t_R PHY_534 ();
 NOR2x1_ASAP7_75t_R _28532_ (.A(_00949_),
    .B(_09762_),
    .Y(_09808_));
 AO21x1_ASAP7_75t_R _28533_ (.A1(_08328_),
    .A2(_09762_),
    .B(_09808_),
    .Y(_02947_));
 TAPCELL_ASAP7_75t_R PHY_533 ();
 NOR2x1_ASAP7_75t_R _28535_ (.A(_00981_),
    .B(_09762_),
    .Y(_09810_));
 AO21x1_ASAP7_75t_R _28536_ (.A1(_08360_),
    .A2(_09762_),
    .B(_09810_),
    .Y(_02948_));
 TAPCELL_ASAP7_75t_R PHY_532 ();
 NOR2x1_ASAP7_75t_R _28538_ (.A(_01015_),
    .B(_09762_),
    .Y(_09812_));
 AO21x1_ASAP7_75t_R _28539_ (.A1(_08406_),
    .A2(_09762_),
    .B(_09812_),
    .Y(_02949_));
 TAPCELL_ASAP7_75t_R PHY_531 ();
 NOR2x1_ASAP7_75t_R _28541_ (.A(_01047_),
    .B(_09762_),
    .Y(_09814_));
 AO21x1_ASAP7_75t_R _28542_ (.A1(_08450_),
    .A2(_09762_),
    .B(_09814_),
    .Y(_02950_));
 TAPCELL_ASAP7_75t_R PHY_530 ();
 AND2x2_ASAP7_75t_R _28544_ (.A(_04748_),
    .B(_09757_),
    .Y(_09816_));
 AO21x1_ASAP7_75t_R _28545_ (.A1(_08481_),
    .A2(_09762_),
    .B(_09816_),
    .Y(_02951_));
 TAPCELL_ASAP7_75t_R PHY_529 ();
 NOR2x1_ASAP7_75t_R _28547_ (.A(_01112_),
    .B(_09762_),
    .Y(_09818_));
 AO21x1_ASAP7_75t_R _28548_ (.A1(_08509_),
    .A2(_09762_),
    .B(_09818_),
    .Y(_02952_));
 TAPCELL_ASAP7_75t_R PHY_528 ();
 NOR2x1_ASAP7_75t_R _28550_ (.A(_01146_),
    .B(_09762_),
    .Y(_09820_));
 AO21x1_ASAP7_75t_R _28551_ (.A1(_08537_),
    .A2(_09762_),
    .B(_09820_),
    .Y(_02953_));
 TAPCELL_ASAP7_75t_R PHY_527 ();
 NOR2x1_ASAP7_75t_R _28553_ (.A(_01178_),
    .B(_09762_),
    .Y(_09822_));
 AO21x1_ASAP7_75t_R _28554_ (.A1(_08563_),
    .A2(_09762_),
    .B(_09822_),
    .Y(_02954_));
 TAPCELL_ASAP7_75t_R PHY_526 ();
 NOR2x1_ASAP7_75t_R _28556_ (.A(_01212_),
    .B(_09762_),
    .Y(_09824_));
 AO21x1_ASAP7_75t_R _28557_ (.A1(net250),
    .A2(_09762_),
    .B(_09824_),
    .Y(_02955_));
 TAPCELL_ASAP7_75t_R PHY_525 ();
 AND2x2_ASAP7_75t_R _28559_ (.A(_05302_),
    .B(_09757_),
    .Y(_09826_));
 AO21x1_ASAP7_75t_R _28560_ (.A1(net2329),
    .A2(_09762_),
    .B(_09826_),
    .Y(_02956_));
 TAPCELL_ASAP7_75t_R PHY_524 ();
 AND2x2_ASAP7_75t_R _28562_ (.A(_08648_),
    .B(_09762_),
    .Y(_09828_));
 AOI21x1_ASAP7_75t_R _28563_ (.A1(_01278_),
    .A2(_09757_),
    .B(_09828_),
    .Y(_02957_));
 OR3x4_ASAP7_75t_R _28564_ (.A(_00184_),
    .B(_14293_),
    .C(_06984_),
    .Y(_09829_));
 TAPCELL_ASAP7_75t_R PHY_523 ();
 NOR2x2_ASAP7_75t_R _28566_ (.A(_06936_),
    .B(_09829_),
    .Y(_09831_));
 TAPCELL_ASAP7_75t_R PHY_522 ();
 TAPCELL_ASAP7_75t_R PHY_521 ();
 NAND2x1_ASAP7_75t_R _28569_ (.A(_07248_),
    .B(_09831_),
    .Y(_09834_));
 OA21x2_ASAP7_75t_R _28570_ (.A1(_13903_),
    .A2(_09831_),
    .B(_09834_),
    .Y(_02958_));
 NOR2x1_ASAP7_75t_R _28571_ (.A(_00248_),
    .B(_09831_),
    .Y(_09835_));
 AO21x1_ASAP7_75t_R _28572_ (.A1(_07384_),
    .A2(_09831_),
    .B(_09835_),
    .Y(_02959_));
 NOR2x1_ASAP7_75t_R _28573_ (.A(_00356_),
    .B(net287),
    .Y(_09836_));
 AO21x1_ASAP7_75t_R _28574_ (.A1(_07472_),
    .A2(net287),
    .B(_09836_),
    .Y(_02960_));
 NOR2x1_ASAP7_75t_R _28575_ (.A(_00387_),
    .B(_09831_),
    .Y(_09837_));
 AO21x1_ASAP7_75t_R _28576_ (.A1(_07552_),
    .A2(_09831_),
    .B(_09837_),
    .Y(_02961_));
 NOR2x1_ASAP7_75t_R _28577_ (.A(_00417_),
    .B(net287),
    .Y(_09838_));
 AO21x1_ASAP7_75t_R _28578_ (.A1(_07608_),
    .A2(net287),
    .B(_09838_),
    .Y(_02962_));
 NOR2x1_ASAP7_75t_R _28579_ (.A(_00447_),
    .B(net287),
    .Y(_09839_));
 AO21x1_ASAP7_75t_R _28580_ (.A1(_07663_),
    .A2(net287),
    .B(_09839_),
    .Y(_02963_));
 NOR2x1_ASAP7_75t_R _28581_ (.A(_00477_),
    .B(net287),
    .Y(_09840_));
 AO21x1_ASAP7_75t_R _28582_ (.A1(_07709_),
    .A2(net287),
    .B(_09840_),
    .Y(_02964_));
 TAPCELL_ASAP7_75t_R PHY_520 ();
 NOR2x1_ASAP7_75t_R _28584_ (.A(_00507_),
    .B(_09831_),
    .Y(_09842_));
 AO21x1_ASAP7_75t_R _28585_ (.A1(net252),
    .A2(net287),
    .B(_09842_),
    .Y(_02965_));
 NOR2x1_ASAP7_75t_R _28586_ (.A(_00537_),
    .B(net287),
    .Y(_09843_));
 AO21x1_ASAP7_75t_R _28587_ (.A1(net257),
    .A2(net287),
    .B(_09843_),
    .Y(_02966_));
 TAPCELL_ASAP7_75t_R PHY_519 ();
 NOR2x1_ASAP7_75t_R _28589_ (.A(_00567_),
    .B(_09831_),
    .Y(_09845_));
 AO21x1_ASAP7_75t_R _28590_ (.A1(net256),
    .A2(_09831_),
    .B(_09845_),
    .Y(_02967_));
 NOR2x1_ASAP7_75t_R _28591_ (.A(_00597_),
    .B(net287),
    .Y(_09846_));
 AO21x1_ASAP7_75t_R _28592_ (.A1(_07903_),
    .A2(net287),
    .B(_09846_),
    .Y(_02968_));
 NOR2x1_ASAP7_75t_R _28593_ (.A(_00627_),
    .B(net287),
    .Y(_09847_));
 AO21x1_ASAP7_75t_R _28594_ (.A1(_07948_),
    .A2(net287),
    .B(_09847_),
    .Y(_02969_));
 NOR2x1_ASAP7_75t_R _28595_ (.A(_00326_),
    .B(net287),
    .Y(_09848_));
 AO21x1_ASAP7_75t_R _28596_ (.A1(_07985_),
    .A2(net287),
    .B(_09848_),
    .Y(_02970_));
 NOR2x1_ASAP7_75t_R _28597_ (.A(_00689_),
    .B(_09831_),
    .Y(_09849_));
 AO21x1_ASAP7_75t_R _28598_ (.A1(net251),
    .A2(_09831_),
    .B(_09849_),
    .Y(_02971_));
 NOR2x1_ASAP7_75t_R _28599_ (.A(_00721_),
    .B(net287),
    .Y(_09850_));
 AO21x1_ASAP7_75t_R _28600_ (.A1(_08068_),
    .A2(net287),
    .B(_09850_),
    .Y(_02972_));
 NOR2x1_ASAP7_75t_R _28601_ (.A(_00754_),
    .B(_09831_),
    .Y(_09851_));
 AO21x1_ASAP7_75t_R _28602_ (.A1(_08110_),
    .A2(_09831_),
    .B(_09851_),
    .Y(_02973_));
 NOR2x1_ASAP7_75t_R _28603_ (.A(_00787_),
    .B(net287),
    .Y(_09852_));
 AO21x1_ASAP7_75t_R _28604_ (.A1(_08151_),
    .A2(net287),
    .B(_09852_),
    .Y(_02974_));
 TAPCELL_ASAP7_75t_R PHY_518 ();
 NOR2x1_ASAP7_75t_R _28606_ (.A(_00820_),
    .B(net287),
    .Y(_09854_));
 AO21x1_ASAP7_75t_R _28607_ (.A1(_08190_),
    .A2(net287),
    .B(_09854_),
    .Y(_02975_));
 NOR2x1_ASAP7_75t_R _28608_ (.A(_00852_),
    .B(_09831_),
    .Y(_09855_));
 AO21x1_ASAP7_75t_R _28609_ (.A1(_08225_),
    .A2(_09831_),
    .B(_09855_),
    .Y(_02976_));
 TAPCELL_ASAP7_75t_R PHY_517 ();
 NOR2x1_ASAP7_75t_R _28611_ (.A(_00885_),
    .B(net287),
    .Y(_09857_));
 AO21x1_ASAP7_75t_R _28612_ (.A1(_08263_),
    .A2(net287),
    .B(_09857_),
    .Y(_02977_));
 NOR2x1_ASAP7_75t_R _28613_ (.A(_00917_),
    .B(_09831_),
    .Y(_09858_));
 AO21x1_ASAP7_75t_R _28614_ (.A1(_08294_),
    .A2(_09831_),
    .B(_09858_),
    .Y(_02978_));
 NOR2x1_ASAP7_75t_R _28615_ (.A(_00950_),
    .B(net287),
    .Y(_09859_));
 AO21x1_ASAP7_75t_R _28616_ (.A1(_08328_),
    .A2(net287),
    .B(_09859_),
    .Y(_02979_));
 NOR2x1_ASAP7_75t_R _28617_ (.A(_00982_),
    .B(_09831_),
    .Y(_09860_));
 AO21x1_ASAP7_75t_R _28618_ (.A1(_08360_),
    .A2(_09831_),
    .B(_09860_),
    .Y(_02980_));
 NOR2x1_ASAP7_75t_R _28619_ (.A(_01016_),
    .B(_09831_),
    .Y(_09861_));
 AO21x1_ASAP7_75t_R _28620_ (.A1(_08406_),
    .A2(_09831_),
    .B(_09861_),
    .Y(_02981_));
 NOR2x1_ASAP7_75t_R _28621_ (.A(_01048_),
    .B(_09831_),
    .Y(_09862_));
 AO21x1_ASAP7_75t_R _28622_ (.A1(_08450_),
    .A2(_09831_),
    .B(_09862_),
    .Y(_02982_));
 NOR2x1_ASAP7_75t_R _28623_ (.A(_01081_),
    .B(net287),
    .Y(_09863_));
 AO21x1_ASAP7_75t_R _28624_ (.A1(_08481_),
    .A2(net287),
    .B(_09863_),
    .Y(_02983_));
 NOR2x1_ASAP7_75t_R _28625_ (.A(_01113_),
    .B(net287),
    .Y(_09864_));
 AO21x1_ASAP7_75t_R _28626_ (.A1(_08509_),
    .A2(net287),
    .B(_09864_),
    .Y(_02984_));
 NOR2x1_ASAP7_75t_R _28627_ (.A(_01147_),
    .B(net287),
    .Y(_09865_));
 AO21x1_ASAP7_75t_R _28628_ (.A1(_08537_),
    .A2(net287),
    .B(_09865_),
    .Y(_02985_));
 NOR2x1_ASAP7_75t_R _28629_ (.A(_01179_),
    .B(_09831_),
    .Y(_09866_));
 AO21x1_ASAP7_75t_R _28630_ (.A1(_08563_),
    .A2(_09831_),
    .B(_09866_),
    .Y(_02986_));
 NOR2x1_ASAP7_75t_R _28631_ (.A(_01213_),
    .B(net287),
    .Y(_09867_));
 AO21x1_ASAP7_75t_R _28632_ (.A1(net250),
    .A2(net287),
    .B(_09867_),
    .Y(_02987_));
 NOR2x1_ASAP7_75t_R _28633_ (.A(_01245_),
    .B(_09831_),
    .Y(_09868_));
 AO21x1_ASAP7_75t_R _28634_ (.A1(net2330),
    .A2(_09831_),
    .B(_09868_),
    .Y(_02988_));
 NAND2x1_ASAP7_75t_R _28635_ (.A(_08648_),
    .B(_09831_),
    .Y(_09869_));
 OA21x2_ASAP7_75t_R _28636_ (.A1(_05478_),
    .A2(_09831_),
    .B(_09869_),
    .Y(_02989_));
 INVx1_ASAP7_75t_R _28637_ (.A(_00295_),
    .Y(_09870_));
 AND2x2_ASAP7_75t_R _28638_ (.A(_00323_),
    .B(_09755_),
    .Y(_09871_));
 AND2x6_ASAP7_75t_R _28639_ (.A(_14176_),
    .B(_00191_),
    .Y(_09872_));
 AND4x2_ASAP7_75t_R _28640_ (.A(_00184_),
    .B(_00194_),
    .C(_09871_),
    .D(_09872_),
    .Y(_09873_));
 TAPCELL_ASAP7_75t_R PHY_516 ();
 TAPCELL_ASAP7_75t_R PHY_515 ();
 TAPCELL_ASAP7_75t_R PHY_514 ();
 NAND2x1_ASAP7_75t_R _28644_ (.A(_07248_),
    .B(_09873_),
    .Y(_09877_));
 OA21x2_ASAP7_75t_R _28645_ (.A1(_09870_),
    .A2(_09873_),
    .B(_09877_),
    .Y(_02990_));
 NOR2x1_ASAP7_75t_R _28646_ (.A(_00249_),
    .B(_09873_),
    .Y(_09878_));
 AO21x1_ASAP7_75t_R _28647_ (.A1(_07384_),
    .A2(_09873_),
    .B(_09878_),
    .Y(_02991_));
 NOR2x1_ASAP7_75t_R _28648_ (.A(_00357_),
    .B(net285),
    .Y(_09879_));
 AO21x1_ASAP7_75t_R _28649_ (.A1(_07472_),
    .A2(net285),
    .B(_09879_),
    .Y(_02992_));
 NOR2x1_ASAP7_75t_R _28650_ (.A(_00388_),
    .B(_09873_),
    .Y(_09880_));
 AO21x1_ASAP7_75t_R _28651_ (.A1(_07552_),
    .A2(_09873_),
    .B(_09880_),
    .Y(_02993_));
 NOR2x1_ASAP7_75t_R _28652_ (.A(_00418_),
    .B(net285),
    .Y(_09881_));
 AO21x1_ASAP7_75t_R _28653_ (.A1(_07608_),
    .A2(net285),
    .B(_09881_),
    .Y(_02994_));
 NOR2x1_ASAP7_75t_R _28654_ (.A(_00448_),
    .B(net285),
    .Y(_09882_));
 AO21x1_ASAP7_75t_R _28655_ (.A1(_07663_),
    .A2(net285),
    .B(_09882_),
    .Y(_02995_));
 NOR2x1_ASAP7_75t_R _28656_ (.A(_00478_),
    .B(net285),
    .Y(_09883_));
 AO21x1_ASAP7_75t_R _28657_ (.A1(_07709_),
    .A2(net285),
    .B(_09883_),
    .Y(_02996_));
 TAPCELL_ASAP7_75t_R PHY_513 ();
 NOR2x1_ASAP7_75t_R _28659_ (.A(_00508_),
    .B(net286),
    .Y(_09885_));
 AO21x1_ASAP7_75t_R _28660_ (.A1(net252),
    .A2(net286),
    .B(_09885_),
    .Y(_02997_));
 NOR2x1_ASAP7_75t_R _28661_ (.A(_00538_),
    .B(net285),
    .Y(_09886_));
 AO21x1_ASAP7_75t_R _28662_ (.A1(net257),
    .A2(net285),
    .B(_09886_),
    .Y(_02998_));
 TAPCELL_ASAP7_75t_R PHY_512 ();
 NOR2x1_ASAP7_75t_R _28664_ (.A(_00568_),
    .B(net286),
    .Y(_09888_));
 AO21x1_ASAP7_75t_R _28665_ (.A1(net256),
    .A2(net286),
    .B(_09888_),
    .Y(_02999_));
 NOR2x1_ASAP7_75t_R _28666_ (.A(_00598_),
    .B(net285),
    .Y(_09889_));
 AO21x1_ASAP7_75t_R _28667_ (.A1(_07903_),
    .A2(net285),
    .B(_09889_),
    .Y(_03000_));
 NOR2x1_ASAP7_75t_R _28668_ (.A(_00628_),
    .B(net285),
    .Y(_09890_));
 AO21x1_ASAP7_75t_R _28669_ (.A1(_07948_),
    .A2(net285),
    .B(_09890_),
    .Y(_03001_));
 NOR2x1_ASAP7_75t_R _28670_ (.A(_00327_),
    .B(net285),
    .Y(_09891_));
 AO21x1_ASAP7_75t_R _28671_ (.A1(_07985_),
    .A2(net285),
    .B(_09891_),
    .Y(_03002_));
 NOR2x1_ASAP7_75t_R _28672_ (.A(_00690_),
    .B(net286),
    .Y(_09892_));
 AO21x1_ASAP7_75t_R _28673_ (.A1(net251),
    .A2(net286),
    .B(_09892_),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _28674_ (.A(_00722_),
    .B(net285),
    .Y(_09893_));
 AO21x1_ASAP7_75t_R _28675_ (.A1(_08068_),
    .A2(net285),
    .B(_09893_),
    .Y(_03004_));
 NOR2x1_ASAP7_75t_R _28676_ (.A(_00755_),
    .B(_09873_),
    .Y(_09894_));
 AO21x1_ASAP7_75t_R _28677_ (.A1(_08110_),
    .A2(_09873_),
    .B(_09894_),
    .Y(_03005_));
 NOR2x1_ASAP7_75t_R _28678_ (.A(_00788_),
    .B(net285),
    .Y(_09895_));
 AO21x1_ASAP7_75t_R _28679_ (.A1(_08151_),
    .A2(net285),
    .B(_09895_),
    .Y(_03006_));
 TAPCELL_ASAP7_75t_R PHY_511 ();
 NOR2x1_ASAP7_75t_R _28681_ (.A(_00821_),
    .B(net285),
    .Y(_09897_));
 AO21x1_ASAP7_75t_R _28682_ (.A1(_08190_),
    .A2(net285),
    .B(_09897_),
    .Y(_03007_));
 NOR2x1_ASAP7_75t_R _28683_ (.A(_00853_),
    .B(_09873_),
    .Y(_09898_));
 AO21x1_ASAP7_75t_R _28684_ (.A1(_08225_),
    .A2(_09873_),
    .B(_09898_),
    .Y(_03008_));
 TAPCELL_ASAP7_75t_R PHY_510 ();
 NOR2x1_ASAP7_75t_R _28686_ (.A(_00886_),
    .B(net285),
    .Y(_09900_));
 AO21x1_ASAP7_75t_R _28687_ (.A1(_08263_),
    .A2(net285),
    .B(_09900_),
    .Y(_03009_));
 NOR2x1_ASAP7_75t_R _28688_ (.A(_00918_),
    .B(_09873_),
    .Y(_09901_));
 AO21x1_ASAP7_75t_R _28689_ (.A1(_08294_),
    .A2(_09873_),
    .B(_09901_),
    .Y(_03010_));
 NOR2x1_ASAP7_75t_R _28690_ (.A(_00951_),
    .B(net285),
    .Y(_09902_));
 AO21x1_ASAP7_75t_R _28691_ (.A1(_08328_),
    .A2(net285),
    .B(_09902_),
    .Y(_03011_));
 NOR2x1_ASAP7_75t_R _28692_ (.A(_00983_),
    .B(_09873_),
    .Y(_09903_));
 AO21x1_ASAP7_75t_R _28693_ (.A1(_08360_),
    .A2(_09873_),
    .B(_09903_),
    .Y(_03012_));
 NOR2x1_ASAP7_75t_R _28694_ (.A(_01017_),
    .B(net286),
    .Y(_09904_));
 AO21x1_ASAP7_75t_R _28695_ (.A1(_08406_),
    .A2(net286),
    .B(_09904_),
    .Y(_03013_));
 NOR2x1_ASAP7_75t_R _28696_ (.A(_01049_),
    .B(_09873_),
    .Y(_09905_));
 AO21x1_ASAP7_75t_R _28697_ (.A1(_08450_),
    .A2(_09873_),
    .B(_09905_),
    .Y(_03014_));
 NOR2x1_ASAP7_75t_R _28698_ (.A(_01082_),
    .B(net285),
    .Y(_09906_));
 AO21x1_ASAP7_75t_R _28699_ (.A1(_08481_),
    .A2(net285),
    .B(_09906_),
    .Y(_03015_));
 NOR2x1_ASAP7_75t_R _28700_ (.A(_01114_),
    .B(net286),
    .Y(_09907_));
 AO21x1_ASAP7_75t_R _28701_ (.A1(_08509_),
    .A2(net286),
    .B(_09907_),
    .Y(_03016_));
 NOR2x1_ASAP7_75t_R _28702_ (.A(_01148_),
    .B(net286),
    .Y(_09908_));
 AO21x1_ASAP7_75t_R _28703_ (.A1(_08537_),
    .A2(net286),
    .B(_09908_),
    .Y(_03017_));
 NOR2x1_ASAP7_75t_R _28704_ (.A(_01180_),
    .B(net286),
    .Y(_09909_));
 AO21x1_ASAP7_75t_R _28705_ (.A1(_08563_),
    .A2(net286),
    .B(_09909_),
    .Y(_03018_));
 NOR2x1_ASAP7_75t_R _28706_ (.A(_01214_),
    .B(net285),
    .Y(_09910_));
 AO21x1_ASAP7_75t_R _28707_ (.A1(_08593_),
    .A2(net285),
    .B(_09910_),
    .Y(_03019_));
 NOR2x1_ASAP7_75t_R _28708_ (.A(_01246_),
    .B(net286),
    .Y(_09911_));
 AO21x1_ASAP7_75t_R _28709_ (.A1(net2329),
    .A2(net286),
    .B(_09911_),
    .Y(_03020_));
 INVx1_ASAP7_75t_R _28710_ (.A(_01280_),
    .Y(_09912_));
 NAND2x1_ASAP7_75t_R _28711_ (.A(_08648_),
    .B(net286),
    .Y(_09913_));
 OA21x2_ASAP7_75t_R _28712_ (.A1(_09912_),
    .A2(net286),
    .B(_09913_),
    .Y(_03021_));
 NAND2x2_ASAP7_75t_R _28713_ (.A(_14176_),
    .B(_00191_),
    .Y(_09914_));
 NOR2x2_ASAP7_75t_R _28714_ (.A(_06985_),
    .B(_09914_),
    .Y(_09915_));
 TAPCELL_ASAP7_75t_R PHY_509 ();
 TAPCELL_ASAP7_75t_R PHY_508 ();
 OR3x1_ASAP7_75t_R _28717_ (.A(_06985_),
    .B(_07248_),
    .C(_09914_),
    .Y(_09918_));
 OAI21x1_ASAP7_75t_R _28718_ (.A1(_00296_),
    .A2(_09915_),
    .B(_09918_),
    .Y(_03022_));
 TAPCELL_ASAP7_75t_R PHY_507 ();
 NOR2x1_ASAP7_75t_R _28720_ (.A(_00250_),
    .B(_09915_),
    .Y(_09920_));
 AO21x1_ASAP7_75t_R _28721_ (.A1(_07384_),
    .A2(_09915_),
    .B(_09920_),
    .Y(_03023_));
 NOR2x1_ASAP7_75t_R _28722_ (.A(_00358_),
    .B(net283),
    .Y(_09921_));
 AO21x1_ASAP7_75t_R _28723_ (.A1(_07472_),
    .A2(net283),
    .B(_09921_),
    .Y(_03024_));
 NOR2x1_ASAP7_75t_R _28724_ (.A(_00389_),
    .B(_09915_),
    .Y(_09922_));
 AO21x1_ASAP7_75t_R _28725_ (.A1(_07552_),
    .A2(_09915_),
    .B(_09922_),
    .Y(_03025_));
 NOR2x1_ASAP7_75t_R _28726_ (.A(_00419_),
    .B(net283),
    .Y(_09923_));
 AO21x1_ASAP7_75t_R _28727_ (.A1(_07608_),
    .A2(net283),
    .B(_09923_),
    .Y(_03026_));
 NOR2x1_ASAP7_75t_R _28728_ (.A(_00449_),
    .B(net283),
    .Y(_09924_));
 AO21x1_ASAP7_75t_R _28729_ (.A1(_07663_),
    .A2(net283),
    .B(_09924_),
    .Y(_03027_));
 NOR2x1_ASAP7_75t_R _28730_ (.A(_00479_),
    .B(net283),
    .Y(_09925_));
 AO21x1_ASAP7_75t_R _28731_ (.A1(_07709_),
    .A2(net283),
    .B(_09925_),
    .Y(_03028_));
 NOR2x1_ASAP7_75t_R _28732_ (.A(_00509_),
    .B(net283),
    .Y(_09926_));
 AO21x1_ASAP7_75t_R _28733_ (.A1(net252),
    .A2(net283),
    .B(_09926_),
    .Y(_03029_));
 NOR2x1_ASAP7_75t_R _28734_ (.A(_00539_),
    .B(net283),
    .Y(_09927_));
 AO21x1_ASAP7_75t_R _28735_ (.A1(net257),
    .A2(net283),
    .B(_09927_),
    .Y(_03030_));
 TAPCELL_ASAP7_75t_R PHY_506 ();
 TAPCELL_ASAP7_75t_R PHY_505 ();
 NOR2x1_ASAP7_75t_R _28738_ (.A(_00569_),
    .B(net284),
    .Y(_09930_));
 AO21x1_ASAP7_75t_R _28739_ (.A1(net256),
    .A2(net284),
    .B(_09930_),
    .Y(_03031_));
 NOR2x1_ASAP7_75t_R _28740_ (.A(_00599_),
    .B(net283),
    .Y(_09931_));
 AO21x1_ASAP7_75t_R _28741_ (.A1(_07903_),
    .A2(net283),
    .B(_09931_),
    .Y(_03032_));
 NOR2x1_ASAP7_75t_R _28742_ (.A(_00629_),
    .B(net283),
    .Y(_09932_));
 AO21x1_ASAP7_75t_R _28743_ (.A1(_07948_),
    .A2(net283),
    .B(_09932_),
    .Y(_03033_));
 NOR2x1_ASAP7_75t_R _28744_ (.A(_00328_),
    .B(net283),
    .Y(_09933_));
 AO21x1_ASAP7_75t_R _28745_ (.A1(_07985_),
    .A2(net283),
    .B(_09933_),
    .Y(_03034_));
 NOR2x1_ASAP7_75t_R _28746_ (.A(_00691_),
    .B(net284),
    .Y(_09934_));
 AO21x1_ASAP7_75t_R _28747_ (.A1(_08026_),
    .A2(net284),
    .B(_09934_),
    .Y(_03035_));
 NOR2x1_ASAP7_75t_R _28748_ (.A(_00723_),
    .B(net284),
    .Y(_09935_));
 AO21x1_ASAP7_75t_R _28749_ (.A1(_08068_),
    .A2(net284),
    .B(_09935_),
    .Y(_03036_));
 NOR2x1_ASAP7_75t_R _28750_ (.A(_00756_),
    .B(_09915_),
    .Y(_09936_));
 AO21x1_ASAP7_75t_R _28751_ (.A1(_08110_),
    .A2(_09915_),
    .B(_09936_),
    .Y(_03037_));
 NOR2x1_ASAP7_75t_R _28752_ (.A(_00789_),
    .B(net283),
    .Y(_09937_));
 AO21x1_ASAP7_75t_R _28753_ (.A1(_08151_),
    .A2(net283),
    .B(_09937_),
    .Y(_03038_));
 NOR2x1_ASAP7_75t_R _28754_ (.A(_00822_),
    .B(net283),
    .Y(_09938_));
 AO21x1_ASAP7_75t_R _28755_ (.A1(_08190_),
    .A2(net283),
    .B(_09938_),
    .Y(_03039_));
 NOR2x1_ASAP7_75t_R _28756_ (.A(_00854_),
    .B(_09915_),
    .Y(_09939_));
 AO21x1_ASAP7_75t_R _28757_ (.A1(_08225_),
    .A2(_09915_),
    .B(_09939_),
    .Y(_03040_));
 TAPCELL_ASAP7_75t_R PHY_504 ();
 TAPCELL_ASAP7_75t_R PHY_503 ();
 NOR2x1_ASAP7_75t_R _28760_ (.A(_00887_),
    .B(net283),
    .Y(_09942_));
 AO21x1_ASAP7_75t_R _28761_ (.A1(_08263_),
    .A2(net283),
    .B(_09942_),
    .Y(_03041_));
 NOR2x1_ASAP7_75t_R _28762_ (.A(_00919_),
    .B(_09915_),
    .Y(_09943_));
 AO21x1_ASAP7_75t_R _28763_ (.A1(_08294_),
    .A2(_09915_),
    .B(_09943_),
    .Y(_03042_));
 NOR2x1_ASAP7_75t_R _28764_ (.A(_00952_),
    .B(net283),
    .Y(_09944_));
 AO21x1_ASAP7_75t_R _28765_ (.A1(_08328_),
    .A2(net283),
    .B(_09944_),
    .Y(_03043_));
 NOR2x1_ASAP7_75t_R _28766_ (.A(_00984_),
    .B(_09915_),
    .Y(_09945_));
 AO21x1_ASAP7_75t_R _28767_ (.A1(_08360_),
    .A2(_09915_),
    .B(_09945_),
    .Y(_03044_));
 NOR2x1_ASAP7_75t_R _28768_ (.A(_01018_),
    .B(net284),
    .Y(_09946_));
 AO21x1_ASAP7_75t_R _28769_ (.A1(_08406_),
    .A2(net284),
    .B(_09946_),
    .Y(_03045_));
 NOR2x1_ASAP7_75t_R _28770_ (.A(_01050_),
    .B(_09915_),
    .Y(_09947_));
 AO21x1_ASAP7_75t_R _28771_ (.A1(_08450_),
    .A2(_09915_),
    .B(_09947_),
    .Y(_03046_));
 NOR2x1_ASAP7_75t_R _28772_ (.A(_01083_),
    .B(net283),
    .Y(_09948_));
 AO21x1_ASAP7_75t_R _28773_ (.A1(_08481_),
    .A2(net283),
    .B(_09948_),
    .Y(_03047_));
 NOR2x1_ASAP7_75t_R _28774_ (.A(_01115_),
    .B(net284),
    .Y(_09949_));
 AO21x1_ASAP7_75t_R _28775_ (.A1(_08509_),
    .A2(net284),
    .B(_09949_),
    .Y(_03048_));
 NOR2x1_ASAP7_75t_R _28776_ (.A(_01149_),
    .B(net284),
    .Y(_09950_));
 AO21x1_ASAP7_75t_R _28777_ (.A1(_08537_),
    .A2(net284),
    .B(_09950_),
    .Y(_03049_));
 NOR2x1_ASAP7_75t_R _28778_ (.A(_01181_),
    .B(net284),
    .Y(_09951_));
 AO21x1_ASAP7_75t_R _28779_ (.A1(_08563_),
    .A2(net284),
    .B(_09951_),
    .Y(_03050_));
 NOR2x1_ASAP7_75t_R _28780_ (.A(_01215_),
    .B(net283),
    .Y(_09952_));
 AO21x1_ASAP7_75t_R _28781_ (.A1(net250),
    .A2(net283),
    .B(_09952_),
    .Y(_03051_));
 NOR2x1_ASAP7_75t_R _28782_ (.A(_01247_),
    .B(net284),
    .Y(_09953_));
 AO21x1_ASAP7_75t_R _28783_ (.A1(net2330),
    .A2(net284),
    .B(_09953_),
    .Y(_03052_));
 OR3x1_ASAP7_75t_R _28784_ (.A(_06985_),
    .B(_08648_),
    .C(_09914_),
    .Y(_09954_));
 OAI21x1_ASAP7_75t_R _28785_ (.A1(_01281_),
    .A2(net284),
    .B(_09954_),
    .Y(_03053_));
 NAND2x2_ASAP7_75t_R _28786_ (.A(_09756_),
    .B(_09872_),
    .Y(_09955_));
 TAPCELL_ASAP7_75t_R PHY_502 ();
 NOR2x1_ASAP7_75t_R _28788_ (.A(_07248_),
    .B(_09955_),
    .Y(_09957_));
 AO21x1_ASAP7_75t_R _28789_ (.A1(_13934_),
    .A2(_09955_),
    .B(_09957_),
    .Y(_03054_));
 AND2x6_ASAP7_75t_R _28790_ (.A(_09756_),
    .B(_09872_),
    .Y(_09958_));
 TAPCELL_ASAP7_75t_R PHY_501 ();
 AND2x2_ASAP7_75t_R _28792_ (.A(_13654_),
    .B(_09955_),
    .Y(_09960_));
 AO21x1_ASAP7_75t_R _28793_ (.A1(_07384_),
    .A2(_09958_),
    .B(_09960_),
    .Y(_03055_));
 AND2x2_ASAP7_75t_R _28794_ (.A(_14878_),
    .B(_09955_),
    .Y(_09961_));
 AO21x1_ASAP7_75t_R _28795_ (.A1(_07472_),
    .A2(_09958_),
    .B(_09961_),
    .Y(_03056_));
 AND2x2_ASAP7_75t_R _28796_ (.A(_14928_),
    .B(_09955_),
    .Y(_09962_));
 AO21x1_ASAP7_75t_R _28797_ (.A1(_07552_),
    .A2(_09958_),
    .B(_09962_),
    .Y(_03057_));
 AND2x2_ASAP7_75t_R _28798_ (.A(_15013_),
    .B(_09955_),
    .Y(_09963_));
 AO21x1_ASAP7_75t_R _28799_ (.A1(_07608_),
    .A2(_09958_),
    .B(_09963_),
    .Y(_03058_));
 AND2x2_ASAP7_75t_R _28800_ (.A(_15065_),
    .B(_09955_),
    .Y(_09964_));
 AO21x1_ASAP7_75t_R _28801_ (.A1(_07663_),
    .A2(_09958_),
    .B(_09964_),
    .Y(_03059_));
 TAPCELL_ASAP7_75t_R PHY_500 ();
 AND2x2_ASAP7_75t_R _28803_ (.A(_14380_),
    .B(_09955_),
    .Y(_09966_));
 AO21x1_ASAP7_75t_R _28804_ (.A1(_07709_),
    .A2(_09958_),
    .B(_09966_),
    .Y(_03060_));
 AND2x2_ASAP7_75t_R _28805_ (.A(_14439_),
    .B(_09955_),
    .Y(_09967_));
 AO21x1_ASAP7_75t_R _28806_ (.A1(net252),
    .A2(_09958_),
    .B(_09967_),
    .Y(_03061_));
 AND2x2_ASAP7_75t_R _28807_ (.A(_15245_),
    .B(_09955_),
    .Y(_09968_));
 AO21x1_ASAP7_75t_R _28808_ (.A1(net257),
    .A2(_09958_),
    .B(_09968_),
    .Y(_03062_));
 AND2x2_ASAP7_75t_R _28809_ (.A(_15297_),
    .B(_09955_),
    .Y(_09969_));
 AO21x1_ASAP7_75t_R _28810_ (.A1(net256),
    .A2(_09958_),
    .B(_09969_),
    .Y(_03063_));
 AND2x2_ASAP7_75t_R _28811_ (.A(_14621_),
    .B(_09955_),
    .Y(_09970_));
 AO21x1_ASAP7_75t_R _28812_ (.A1(_07903_),
    .A2(_09958_),
    .B(_09970_),
    .Y(_03064_));
 TAPCELL_ASAP7_75t_R PHY_499 ();
 AND2x2_ASAP7_75t_R _28814_ (.A(_14734_),
    .B(_09955_),
    .Y(_09972_));
 AO21x1_ASAP7_75t_R _28815_ (.A1(_07948_),
    .A2(_09958_),
    .B(_09972_),
    .Y(_03065_));
 TAPCELL_ASAP7_75t_R PHY_498 ();
 AND3x1_ASAP7_75t_R _28817_ (.A(_07961_),
    .B(_07984_),
    .C(_09958_),
    .Y(_09974_));
 AO21x1_ASAP7_75t_R _28818_ (.A1(_14019_),
    .A2(_09955_),
    .B(_09974_),
    .Y(_03066_));
 AND2x2_ASAP7_75t_R _28819_ (.A(_15523_),
    .B(_09955_),
    .Y(_09975_));
 AO21x1_ASAP7_75t_R _28820_ (.A1(net251),
    .A2(_09958_),
    .B(_09975_),
    .Y(_03067_));
 AND2x2_ASAP7_75t_R _28821_ (.A(_15679_),
    .B(_09955_),
    .Y(_09976_));
 AO21x1_ASAP7_75t_R _28822_ (.A1(_08068_),
    .A2(_09958_),
    .B(_09976_),
    .Y(_03068_));
 AND2x2_ASAP7_75t_R _28823_ (.A(_15795_),
    .B(_09955_),
    .Y(_09977_));
 AO21x1_ASAP7_75t_R _28824_ (.A1(_08110_),
    .A2(_09958_),
    .B(_09977_),
    .Y(_03069_));
 AND2x2_ASAP7_75t_R _28825_ (.A(_15917_),
    .B(_09955_),
    .Y(_09978_));
 AO21x1_ASAP7_75t_R _28826_ (.A1(_08151_),
    .A2(_09958_),
    .B(_09978_),
    .Y(_03070_));
 TAPCELL_ASAP7_75t_R PHY_497 ();
 AND2x2_ASAP7_75t_R _28828_ (.A(_16046_),
    .B(_09955_),
    .Y(_09980_));
 AO21x1_ASAP7_75t_R _28829_ (.A1(_08190_),
    .A2(_09958_),
    .B(_09980_),
    .Y(_03071_));
 AND2x2_ASAP7_75t_R _28830_ (.A(_16165_),
    .B(_09955_),
    .Y(_09981_));
 AO21x1_ASAP7_75t_R _28831_ (.A1(_08225_),
    .A2(_09958_),
    .B(_09981_),
    .Y(_03072_));
 AND2x2_ASAP7_75t_R _28832_ (.A(_16318_),
    .B(_09955_),
    .Y(_09982_));
 AO21x1_ASAP7_75t_R _28833_ (.A1(_08263_),
    .A2(_09958_),
    .B(_09982_),
    .Y(_03073_));
 AND2x2_ASAP7_75t_R _28834_ (.A(_16410_),
    .B(_09955_),
    .Y(_09983_));
 AO21x1_ASAP7_75t_R _28835_ (.A1(_08294_),
    .A2(_09958_),
    .B(_09983_),
    .Y(_03074_));
 AND2x2_ASAP7_75t_R _28836_ (.A(_16531_),
    .B(_09955_),
    .Y(_09984_));
 AO21x1_ASAP7_75t_R _28837_ (.A1(_08328_),
    .A2(_09958_),
    .B(_09984_),
    .Y(_03075_));
 AND2x2_ASAP7_75t_R _28838_ (.A(_16635_),
    .B(_09955_),
    .Y(_09985_));
 AO21x1_ASAP7_75t_R _28839_ (.A1(_08360_),
    .A2(_09958_),
    .B(_09985_),
    .Y(_03076_));
 AND2x2_ASAP7_75t_R _28840_ (.A(_04532_),
    .B(_09955_),
    .Y(_09986_));
 AO21x1_ASAP7_75t_R _28841_ (.A1(_08406_),
    .A2(_09958_),
    .B(_09986_),
    .Y(_03077_));
 AND2x2_ASAP7_75t_R _28842_ (.A(_04652_),
    .B(_09955_),
    .Y(_09987_));
 AO21x1_ASAP7_75t_R _28843_ (.A1(_08450_),
    .A2(_09958_),
    .B(_09987_),
    .Y(_03078_));
 AND2x2_ASAP7_75t_R _28844_ (.A(_04764_),
    .B(_09955_),
    .Y(_09988_));
 AO21x1_ASAP7_75t_R _28845_ (.A1(_08481_),
    .A2(_09958_),
    .B(_09988_),
    .Y(_03079_));
 AND2x2_ASAP7_75t_R _28846_ (.A(_04868_),
    .B(_09955_),
    .Y(_09989_));
 AO21x1_ASAP7_75t_R _28847_ (.A1(_08509_),
    .A2(_09958_),
    .B(_09989_),
    .Y(_03080_));
 AND2x2_ASAP7_75t_R _28848_ (.A(_04983_),
    .B(_09955_),
    .Y(_09990_));
 AO21x1_ASAP7_75t_R _28849_ (.A1(_08537_),
    .A2(_09958_),
    .B(_09990_),
    .Y(_03081_));
 AND2x2_ASAP7_75t_R _28850_ (.A(_05092_),
    .B(_09955_),
    .Y(_09991_));
 AO21x1_ASAP7_75t_R _28851_ (.A1(_08563_),
    .A2(_09958_),
    .B(_09991_),
    .Y(_03082_));
 AND2x2_ASAP7_75t_R _28852_ (.A(_05200_),
    .B(_09955_),
    .Y(_09992_));
 AO21x1_ASAP7_75t_R _28853_ (.A1(_08593_),
    .A2(_09958_),
    .B(_09992_),
    .Y(_03083_));
 AND2x2_ASAP7_75t_R _28854_ (.A(_05311_),
    .B(_09955_),
    .Y(_09993_));
 AO21x1_ASAP7_75t_R _28855_ (.A1(net2329),
    .A2(_09958_),
    .B(_09993_),
    .Y(_03084_));
 TAPCELL_ASAP7_75t_R PHY_496 ();
 NOR2x1_ASAP7_75t_R _28857_ (.A(_08648_),
    .B(_09955_),
    .Y(_09995_));
 AO21x1_ASAP7_75t_R _28858_ (.A1(_05433_),
    .A2(_09955_),
    .B(_09995_),
    .Y(_03085_));
 NOR2x2_ASAP7_75t_R _28859_ (.A(_09829_),
    .B(_09914_),
    .Y(_09996_));
 TAPCELL_ASAP7_75t_R PHY_495 ();
 TAPCELL_ASAP7_75t_R PHY_494 ();
 NAND2x1_ASAP7_75t_R _28862_ (.A(_07248_),
    .B(_09996_),
    .Y(_09999_));
 OA21x2_ASAP7_75t_R _28863_ (.A1(_13927_),
    .A2(_09996_),
    .B(_09999_),
    .Y(_03086_));
 NOR2x1_ASAP7_75t_R _28864_ (.A(_00252_),
    .B(_09996_),
    .Y(_10000_));
 AO21x1_ASAP7_75t_R _28865_ (.A1(_07384_),
    .A2(_09996_),
    .B(_10000_),
    .Y(_03087_));
 NOR2x1_ASAP7_75t_R _28866_ (.A(_00360_),
    .B(net281),
    .Y(_10001_));
 AO21x1_ASAP7_75t_R _28867_ (.A1(_07472_),
    .A2(net281),
    .B(_10001_),
    .Y(_03088_));
 NOR2x1_ASAP7_75t_R _28868_ (.A(_00391_),
    .B(_09996_),
    .Y(_10002_));
 AO21x1_ASAP7_75t_R _28869_ (.A1(_07552_),
    .A2(_09996_),
    .B(_10002_),
    .Y(_03089_));
 NOR2x1_ASAP7_75t_R _28870_ (.A(_00421_),
    .B(net281),
    .Y(_10003_));
 AO21x1_ASAP7_75t_R _28871_ (.A1(_07608_),
    .A2(net281),
    .B(_10003_),
    .Y(_03090_));
 NOR2x1_ASAP7_75t_R _28872_ (.A(_00451_),
    .B(net281),
    .Y(_10004_));
 AO21x1_ASAP7_75t_R _28873_ (.A1(_07663_),
    .A2(net281),
    .B(_10004_),
    .Y(_03091_));
 NOR2x1_ASAP7_75t_R _28874_ (.A(_00481_),
    .B(net281),
    .Y(_10005_));
 AO21x1_ASAP7_75t_R _28875_ (.A1(_07709_),
    .A2(net281),
    .B(_10005_),
    .Y(_03092_));
 TAPCELL_ASAP7_75t_R PHY_493 ();
 NOR2x1_ASAP7_75t_R _28877_ (.A(_00511_),
    .B(net282),
    .Y(_10007_));
 AO21x1_ASAP7_75t_R _28878_ (.A1(net252),
    .A2(net282),
    .B(_10007_),
    .Y(_03093_));
 NOR2x1_ASAP7_75t_R _28879_ (.A(_00541_),
    .B(net282),
    .Y(_10008_));
 AO21x1_ASAP7_75t_R _28880_ (.A1(net257),
    .A2(net282),
    .B(_10008_),
    .Y(_03094_));
 TAPCELL_ASAP7_75t_R PHY_492 ();
 NOR2x1_ASAP7_75t_R _28882_ (.A(_00571_),
    .B(net282),
    .Y(_10010_));
 AO21x1_ASAP7_75t_R _28883_ (.A1(net256),
    .A2(net282),
    .B(_10010_),
    .Y(_03095_));
 NOR2x1_ASAP7_75t_R _28884_ (.A(_00601_),
    .B(net281),
    .Y(_10011_));
 AO21x1_ASAP7_75t_R _28885_ (.A1(_07903_),
    .A2(net281),
    .B(_10011_),
    .Y(_03096_));
 NOR2x1_ASAP7_75t_R _28886_ (.A(_00631_),
    .B(net281),
    .Y(_10012_));
 AO21x1_ASAP7_75t_R _28887_ (.A1(_07948_),
    .A2(net281),
    .B(_10012_),
    .Y(_03097_));
 NOR2x1_ASAP7_75t_R _28888_ (.A(_00330_),
    .B(net281),
    .Y(_10013_));
 AO21x1_ASAP7_75t_R _28889_ (.A1(_07985_),
    .A2(net281),
    .B(_10013_),
    .Y(_03098_));
 NOR2x1_ASAP7_75t_R _28890_ (.A(_00693_),
    .B(net282),
    .Y(_10014_));
 AO21x1_ASAP7_75t_R _28891_ (.A1(_08026_),
    .A2(net282),
    .B(_10014_),
    .Y(_03099_));
 NOR2x1_ASAP7_75t_R _28892_ (.A(_00725_),
    .B(net281),
    .Y(_10015_));
 AO21x1_ASAP7_75t_R _28893_ (.A1(_08068_),
    .A2(net281),
    .B(_10015_),
    .Y(_03100_));
 NOR2x1_ASAP7_75t_R _28894_ (.A(_00758_),
    .B(_09996_),
    .Y(_10016_));
 AO21x1_ASAP7_75t_R _28895_ (.A1(_08110_),
    .A2(_09996_),
    .B(_10016_),
    .Y(_03101_));
 NOR2x1_ASAP7_75t_R _28896_ (.A(_00791_),
    .B(net281),
    .Y(_10017_));
 AO21x1_ASAP7_75t_R _28897_ (.A1(_08151_),
    .A2(net281),
    .B(_10017_),
    .Y(_03102_));
 TAPCELL_ASAP7_75t_R PHY_491 ();
 NOR2x1_ASAP7_75t_R _28899_ (.A(_00824_),
    .B(net281),
    .Y(_10019_));
 AO21x1_ASAP7_75t_R _28900_ (.A1(_08190_),
    .A2(net281),
    .B(_10019_),
    .Y(_03103_));
 NOR2x1_ASAP7_75t_R _28901_ (.A(_00856_),
    .B(_09996_),
    .Y(_10020_));
 AO21x1_ASAP7_75t_R _28902_ (.A1(_08225_),
    .A2(_09996_),
    .B(_10020_),
    .Y(_03104_));
 TAPCELL_ASAP7_75t_R PHY_490 ();
 NOR2x1_ASAP7_75t_R _28904_ (.A(_00889_),
    .B(net281),
    .Y(_10022_));
 AO21x1_ASAP7_75t_R _28905_ (.A1(_08263_),
    .A2(net281),
    .B(_10022_),
    .Y(_03105_));
 NOR2x1_ASAP7_75t_R _28906_ (.A(_00921_),
    .B(_09996_),
    .Y(_10023_));
 AO21x1_ASAP7_75t_R _28907_ (.A1(_08294_),
    .A2(_09996_),
    .B(_10023_),
    .Y(_03106_));
 NOR2x1_ASAP7_75t_R _28908_ (.A(_00954_),
    .B(net281),
    .Y(_10024_));
 AO21x1_ASAP7_75t_R _28909_ (.A1(_08328_),
    .A2(net281),
    .B(_10024_),
    .Y(_03107_));
 NOR2x1_ASAP7_75t_R _28910_ (.A(_00986_),
    .B(_09996_),
    .Y(_10025_));
 AO21x1_ASAP7_75t_R _28911_ (.A1(_08360_),
    .A2(_09996_),
    .B(_10025_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _28912_ (.A(_01020_),
    .B(net282),
    .Y(_10026_));
 AO21x1_ASAP7_75t_R _28913_ (.A1(_08406_),
    .A2(net282),
    .B(_10026_),
    .Y(_03109_));
 NOR2x1_ASAP7_75t_R _28914_ (.A(_01052_),
    .B(_09996_),
    .Y(_10027_));
 AO21x1_ASAP7_75t_R _28915_ (.A1(_08450_),
    .A2(_09996_),
    .B(_10027_),
    .Y(_03110_));
 NOR2x1_ASAP7_75t_R _28916_ (.A(_01085_),
    .B(net281),
    .Y(_10028_));
 AO21x1_ASAP7_75t_R _28917_ (.A1(_08481_),
    .A2(net281),
    .B(_10028_),
    .Y(_03111_));
 NOR2x1_ASAP7_75t_R _28918_ (.A(_01117_),
    .B(net281),
    .Y(_10029_));
 AO21x1_ASAP7_75t_R _28919_ (.A1(_08509_),
    .A2(net281),
    .B(_10029_),
    .Y(_03112_));
 NOR2x1_ASAP7_75t_R _28920_ (.A(_01151_),
    .B(net282),
    .Y(_10030_));
 AO21x1_ASAP7_75t_R _28921_ (.A1(_08537_),
    .A2(net282),
    .B(_10030_),
    .Y(_03113_));
 NOR2x1_ASAP7_75t_R _28922_ (.A(_01183_),
    .B(net282),
    .Y(_10031_));
 AO21x1_ASAP7_75t_R _28923_ (.A1(_08563_),
    .A2(net282),
    .B(_10031_),
    .Y(_03114_));
 NOR2x1_ASAP7_75t_R _28924_ (.A(_01217_),
    .B(net281),
    .Y(_10032_));
 AO21x1_ASAP7_75t_R _28925_ (.A1(net250),
    .A2(net281),
    .B(_10032_),
    .Y(_03115_));
 NOR2x1_ASAP7_75t_R _28926_ (.A(_01249_),
    .B(net282),
    .Y(_10033_));
 AO21x1_ASAP7_75t_R _28927_ (.A1(net2330),
    .A2(net282),
    .B(_10033_),
    .Y(_03116_));
 NAND2x1_ASAP7_75t_R _28928_ (.A(_08648_),
    .B(net282),
    .Y(_10034_));
 OA21x2_ASAP7_75t_R _28929_ (.A1(_05436_),
    .A2(net282),
    .B(_10034_),
    .Y(_03117_));
 INVx1_ASAP7_75t_R _28930_ (.A(_00299_),
    .Y(_10035_));
 AND2x6_ASAP7_75t_R _28931_ (.A(_00187_),
    .B(_14182_),
    .Y(_10036_));
 AND4x2_ASAP7_75t_R _28932_ (.A(_00184_),
    .B(_00194_),
    .C(_09871_),
    .D(_10036_),
    .Y(_10037_));
 TAPCELL_ASAP7_75t_R PHY_489 ();
 TAPCELL_ASAP7_75t_R PHY_488 ();
 TAPCELL_ASAP7_75t_R PHY_487 ();
 NAND2x1_ASAP7_75t_R _28936_ (.A(_07248_),
    .B(_10037_),
    .Y(_10041_));
 OA21x2_ASAP7_75t_R _28937_ (.A1(_10035_),
    .A2(_10037_),
    .B(_10041_),
    .Y(_03118_));
 NOR2x1_ASAP7_75t_R _28938_ (.A(_00253_),
    .B(_10037_),
    .Y(_10042_));
 AO21x1_ASAP7_75t_R _28939_ (.A1(_07384_),
    .A2(_10037_),
    .B(_10042_),
    .Y(_03119_));
 NOR2x1_ASAP7_75t_R _28940_ (.A(_00361_),
    .B(net279),
    .Y(_10043_));
 AO21x1_ASAP7_75t_R _28941_ (.A1(_07472_),
    .A2(net279),
    .B(_10043_),
    .Y(_03120_));
 NOR2x1_ASAP7_75t_R _28942_ (.A(_00392_),
    .B(_10037_),
    .Y(_10044_));
 AO21x1_ASAP7_75t_R _28943_ (.A1(_07552_),
    .A2(_10037_),
    .B(_10044_),
    .Y(_03121_));
 NOR2x1_ASAP7_75t_R _28944_ (.A(_00422_),
    .B(net279),
    .Y(_10045_));
 AO21x1_ASAP7_75t_R _28945_ (.A1(_07608_),
    .A2(net279),
    .B(_10045_),
    .Y(_03122_));
 NOR2x1_ASAP7_75t_R _28946_ (.A(_00452_),
    .B(net279),
    .Y(_10046_));
 AO21x1_ASAP7_75t_R _28947_ (.A1(_07663_),
    .A2(net279),
    .B(_10046_),
    .Y(_03123_));
 NOR2x1_ASAP7_75t_R _28948_ (.A(_00482_),
    .B(net279),
    .Y(_10047_));
 AO21x1_ASAP7_75t_R _28949_ (.A1(_07709_),
    .A2(net279),
    .B(_10047_),
    .Y(_03124_));
 TAPCELL_ASAP7_75t_R PHY_486 ();
 NOR2x1_ASAP7_75t_R _28951_ (.A(_00512_),
    .B(net280),
    .Y(_10049_));
 AO21x1_ASAP7_75t_R _28952_ (.A1(net252),
    .A2(net280),
    .B(_10049_),
    .Y(_03125_));
 NOR2x1_ASAP7_75t_R _28953_ (.A(_00542_),
    .B(net280),
    .Y(_10050_));
 AO21x1_ASAP7_75t_R _28954_ (.A1(net257),
    .A2(net280),
    .B(_10050_),
    .Y(_03126_));
 TAPCELL_ASAP7_75t_R PHY_485 ();
 NOR2x1_ASAP7_75t_R _28956_ (.A(_00572_),
    .B(_10037_),
    .Y(_10052_));
 AO21x1_ASAP7_75t_R _28957_ (.A1(net256),
    .A2(_10037_),
    .B(_10052_),
    .Y(_03127_));
 NOR2x1_ASAP7_75t_R _28958_ (.A(_00602_),
    .B(net279),
    .Y(_10053_));
 AO21x1_ASAP7_75t_R _28959_ (.A1(_07903_),
    .A2(net279),
    .B(_10053_),
    .Y(_03128_));
 NOR2x1_ASAP7_75t_R _28960_ (.A(_00632_),
    .B(net279),
    .Y(_10054_));
 AO21x1_ASAP7_75t_R _28961_ (.A1(_07948_),
    .A2(net279),
    .B(_10054_),
    .Y(_03129_));
 NOR2x1_ASAP7_75t_R _28962_ (.A(_00331_),
    .B(net279),
    .Y(_10055_));
 AO21x1_ASAP7_75t_R _28963_ (.A1(_07985_),
    .A2(net279),
    .B(_10055_),
    .Y(_03130_));
 NOR2x1_ASAP7_75t_R _28964_ (.A(_00694_),
    .B(net280),
    .Y(_10056_));
 AO21x1_ASAP7_75t_R _28965_ (.A1(net251),
    .A2(net280),
    .B(_10056_),
    .Y(_03131_));
 NOR2x1_ASAP7_75t_R _28966_ (.A(_00726_),
    .B(net280),
    .Y(_10057_));
 AO21x1_ASAP7_75t_R _28967_ (.A1(_08068_),
    .A2(net280),
    .B(_10057_),
    .Y(_03132_));
 NOR2x1_ASAP7_75t_R _28968_ (.A(_00759_),
    .B(_10037_),
    .Y(_10058_));
 AO21x1_ASAP7_75t_R _28969_ (.A1(_08110_),
    .A2(_10037_),
    .B(_10058_),
    .Y(_03133_));
 NOR2x1_ASAP7_75t_R _28970_ (.A(_00792_),
    .B(net280),
    .Y(_10059_));
 AO21x1_ASAP7_75t_R _28971_ (.A1(_08151_),
    .A2(net280),
    .B(_10059_),
    .Y(_03134_));
 TAPCELL_ASAP7_75t_R PHY_484 ();
 NOR2x1_ASAP7_75t_R _28973_ (.A(_00825_),
    .B(net280),
    .Y(_10061_));
 AO21x1_ASAP7_75t_R _28974_ (.A1(_08190_),
    .A2(net280),
    .B(_10061_),
    .Y(_03135_));
 NOR2x1_ASAP7_75t_R _28975_ (.A(_00857_),
    .B(_10037_),
    .Y(_10062_));
 AO21x1_ASAP7_75t_R _28976_ (.A1(_08225_),
    .A2(_10037_),
    .B(_10062_),
    .Y(_03136_));
 TAPCELL_ASAP7_75t_R PHY_483 ();
 NOR2x1_ASAP7_75t_R _28978_ (.A(_00890_),
    .B(net279),
    .Y(_10064_));
 AO21x1_ASAP7_75t_R _28979_ (.A1(_08263_),
    .A2(net279),
    .B(_10064_),
    .Y(_03137_));
 NOR2x1_ASAP7_75t_R _28980_ (.A(_00922_),
    .B(_10037_),
    .Y(_10065_));
 AO21x1_ASAP7_75t_R _28981_ (.A1(_08294_),
    .A2(_10037_),
    .B(_10065_),
    .Y(_03138_));
 NOR2x1_ASAP7_75t_R _28982_ (.A(_00955_),
    .B(net279),
    .Y(_10066_));
 AO21x1_ASAP7_75t_R _28983_ (.A1(_08328_),
    .A2(net279),
    .B(_10066_),
    .Y(_03139_));
 NOR2x1_ASAP7_75t_R _28984_ (.A(_00987_),
    .B(_10037_),
    .Y(_10067_));
 AO21x1_ASAP7_75t_R _28985_ (.A1(_08360_),
    .A2(_10037_),
    .B(_10067_),
    .Y(_03140_));
 NOR2x1_ASAP7_75t_R _28986_ (.A(_01021_),
    .B(net280),
    .Y(_10068_));
 AO21x1_ASAP7_75t_R _28987_ (.A1(_08406_),
    .A2(net280),
    .B(_10068_),
    .Y(_03141_));
 NOR2x1_ASAP7_75t_R _28988_ (.A(_01053_),
    .B(_10037_),
    .Y(_10069_));
 AO21x1_ASAP7_75t_R _28989_ (.A1(_08450_),
    .A2(_10037_),
    .B(_10069_),
    .Y(_03142_));
 NOR2x1_ASAP7_75t_R _28990_ (.A(_01086_),
    .B(net279),
    .Y(_10070_));
 AO21x1_ASAP7_75t_R _28991_ (.A1(_08481_),
    .A2(net279),
    .B(_10070_),
    .Y(_03143_));
 NOR2x1_ASAP7_75t_R _28992_ (.A(_01118_),
    .B(net280),
    .Y(_10071_));
 AO21x1_ASAP7_75t_R _28993_ (.A1(_08509_),
    .A2(net280),
    .B(_10071_),
    .Y(_03144_));
 NOR2x1_ASAP7_75t_R _28994_ (.A(_01152_),
    .B(net280),
    .Y(_10072_));
 AO21x1_ASAP7_75t_R _28995_ (.A1(_08537_),
    .A2(net280),
    .B(_10072_),
    .Y(_03145_));
 NOR2x1_ASAP7_75t_R _28996_ (.A(_01184_),
    .B(net280),
    .Y(_10073_));
 AO21x1_ASAP7_75t_R _28997_ (.A1(_08563_),
    .A2(net280),
    .B(_10073_),
    .Y(_03146_));
 NOR2x1_ASAP7_75t_R _28998_ (.A(_01218_),
    .B(net279),
    .Y(_10074_));
 AO21x1_ASAP7_75t_R _28999_ (.A1(net250),
    .A2(net279),
    .B(_10074_),
    .Y(_03147_));
 NOR2x1_ASAP7_75t_R _29000_ (.A(_01250_),
    .B(net280),
    .Y(_10075_));
 AO21x1_ASAP7_75t_R _29001_ (.A1(net2329),
    .A2(net280),
    .B(_10075_),
    .Y(_03148_));
 NAND2x1_ASAP7_75t_R _29002_ (.A(_08648_),
    .B(net279),
    .Y(_10076_));
 OA21x2_ASAP7_75t_R _29003_ (.A1(_05464_),
    .A2(net280),
    .B(_10076_),
    .Y(_03149_));
 NAND2x2_ASAP7_75t_R _29004_ (.A(_00187_),
    .B(_14182_),
    .Y(_10077_));
 NOR2x2_ASAP7_75t_R _29005_ (.A(_06985_),
    .B(_10077_),
    .Y(_10078_));
 TAPCELL_ASAP7_75t_R PHY_482 ();
 OR3x1_ASAP7_75t_R _29007_ (.A(_06985_),
    .B(_07248_),
    .C(_10077_),
    .Y(_10080_));
 OAI21x1_ASAP7_75t_R _29008_ (.A1(_00300_),
    .A2(_10078_),
    .B(_10080_),
    .Y(_03150_));
 TAPCELL_ASAP7_75t_R PHY_481 ();
 NOR2x1_ASAP7_75t_R _29010_ (.A(_00254_),
    .B(_10078_),
    .Y(_10082_));
 AO21x1_ASAP7_75t_R _29011_ (.A1(_07384_),
    .A2(_10078_),
    .B(_10082_),
    .Y(_03151_));
 NOR2x1_ASAP7_75t_R _29012_ (.A(_00362_),
    .B(net277),
    .Y(_10083_));
 AO21x1_ASAP7_75t_R _29013_ (.A1(_07472_),
    .A2(net277),
    .B(_10083_),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _29014_ (.A(_00393_),
    .B(_10078_),
    .Y(_10084_));
 AO21x1_ASAP7_75t_R _29015_ (.A1(_07552_),
    .A2(_10078_),
    .B(_10084_),
    .Y(_03153_));
 NOR2x1_ASAP7_75t_R _29016_ (.A(_00423_),
    .B(net277),
    .Y(_10085_));
 AO21x1_ASAP7_75t_R _29017_ (.A1(_07608_),
    .A2(net277),
    .B(_10085_),
    .Y(_03154_));
 NOR2x1_ASAP7_75t_R _29018_ (.A(_00453_),
    .B(net277),
    .Y(_10086_));
 AO21x1_ASAP7_75t_R _29019_ (.A1(_07663_),
    .A2(net277),
    .B(_10086_),
    .Y(_03155_));
 NOR2x1_ASAP7_75t_R _29020_ (.A(_00483_),
    .B(net277),
    .Y(_10087_));
 AO21x1_ASAP7_75t_R _29021_ (.A1(_07709_),
    .A2(net277),
    .B(_10087_),
    .Y(_03156_));
 NOR2x1_ASAP7_75t_R _29022_ (.A(_00513_),
    .B(net278),
    .Y(_10088_));
 AO21x1_ASAP7_75t_R _29023_ (.A1(net252),
    .A2(net278),
    .B(_10088_),
    .Y(_03157_));
 NOR2x1_ASAP7_75t_R _29024_ (.A(_00543_),
    .B(net278),
    .Y(_10089_));
 AO21x1_ASAP7_75t_R _29025_ (.A1(net257),
    .A2(net278),
    .B(_10089_),
    .Y(_03158_));
 TAPCELL_ASAP7_75t_R PHY_480 ();
 TAPCELL_ASAP7_75t_R PHY_479 ();
 NOR2x1_ASAP7_75t_R _29028_ (.A(_00573_),
    .B(_10078_),
    .Y(_10092_));
 AO21x1_ASAP7_75t_R _29029_ (.A1(net256),
    .A2(_10078_),
    .B(_10092_),
    .Y(_03159_));
 NOR2x1_ASAP7_75t_R _29030_ (.A(_00603_),
    .B(net277),
    .Y(_10093_));
 AO21x1_ASAP7_75t_R _29031_ (.A1(_07903_),
    .A2(net277),
    .B(_10093_),
    .Y(_03160_));
 NOR2x1_ASAP7_75t_R _29032_ (.A(_00633_),
    .B(net277),
    .Y(_10094_));
 AO21x1_ASAP7_75t_R _29033_ (.A1(_07948_),
    .A2(net277),
    .B(_10094_),
    .Y(_03161_));
 NOR2x1_ASAP7_75t_R _29034_ (.A(_00332_),
    .B(net277),
    .Y(_10095_));
 AO21x1_ASAP7_75t_R _29035_ (.A1(_07985_),
    .A2(net277),
    .B(_10095_),
    .Y(_03162_));
 NOR2x1_ASAP7_75t_R _29036_ (.A(_00695_),
    .B(net278),
    .Y(_10096_));
 AO21x1_ASAP7_75t_R _29037_ (.A1(net251),
    .A2(net278),
    .B(_10096_),
    .Y(_03163_));
 NOR2x1_ASAP7_75t_R _29038_ (.A(_00727_),
    .B(net277),
    .Y(_10097_));
 AO21x1_ASAP7_75t_R _29039_ (.A1(_08068_),
    .A2(net277),
    .B(_10097_),
    .Y(_03164_));
 NOR2x1_ASAP7_75t_R _29040_ (.A(_00760_),
    .B(_10078_),
    .Y(_10098_));
 AO21x1_ASAP7_75t_R _29041_ (.A1(_08110_),
    .A2(_10078_),
    .B(_10098_),
    .Y(_03165_));
 NOR2x1_ASAP7_75t_R _29042_ (.A(_00793_),
    .B(net277),
    .Y(_10099_));
 AO21x1_ASAP7_75t_R _29043_ (.A1(_08151_),
    .A2(net277),
    .B(_10099_),
    .Y(_03166_));
 NOR2x1_ASAP7_75t_R _29044_ (.A(_00826_),
    .B(net277),
    .Y(_10100_));
 AO21x1_ASAP7_75t_R _29045_ (.A1(_08190_),
    .A2(net277),
    .B(_10100_),
    .Y(_03167_));
 NOR2x1_ASAP7_75t_R _29046_ (.A(_00858_),
    .B(_10078_),
    .Y(_10101_));
 AO21x1_ASAP7_75t_R _29047_ (.A1(_08225_),
    .A2(_10078_),
    .B(_10101_),
    .Y(_03168_));
 TAPCELL_ASAP7_75t_R PHY_478 ();
 TAPCELL_ASAP7_75t_R PHY_477 ();
 NOR2x1_ASAP7_75t_R _29050_ (.A(_00891_),
    .B(net277),
    .Y(_10104_));
 AO21x1_ASAP7_75t_R _29051_ (.A1(_08263_),
    .A2(net277),
    .B(_10104_),
    .Y(_03169_));
 NOR2x1_ASAP7_75t_R _29052_ (.A(_00923_),
    .B(_10078_),
    .Y(_10105_));
 AO21x1_ASAP7_75t_R _29053_ (.A1(_08294_),
    .A2(_10078_),
    .B(_10105_),
    .Y(_03170_));
 NOR2x1_ASAP7_75t_R _29054_ (.A(_00956_),
    .B(net277),
    .Y(_10106_));
 AO21x1_ASAP7_75t_R _29055_ (.A1(_08328_),
    .A2(net277),
    .B(_10106_),
    .Y(_03171_));
 NOR2x1_ASAP7_75t_R _29056_ (.A(_00988_),
    .B(_10078_),
    .Y(_10107_));
 AO21x1_ASAP7_75t_R _29057_ (.A1(_08360_),
    .A2(_10078_),
    .B(_10107_),
    .Y(_03172_));
 NOR2x1_ASAP7_75t_R _29058_ (.A(_01022_),
    .B(net278),
    .Y(_10108_));
 AO21x1_ASAP7_75t_R _29059_ (.A1(_08406_),
    .A2(net278),
    .B(_10108_),
    .Y(_03173_));
 NOR2x1_ASAP7_75t_R _29060_ (.A(_01054_),
    .B(_10078_),
    .Y(_10109_));
 AO21x1_ASAP7_75t_R _29061_ (.A1(_08450_),
    .A2(_10078_),
    .B(_10109_),
    .Y(_03174_));
 NOR2x1_ASAP7_75t_R _29062_ (.A(_01087_),
    .B(net277),
    .Y(_10110_));
 AO21x1_ASAP7_75t_R _29063_ (.A1(_08481_),
    .A2(net277),
    .B(_10110_),
    .Y(_03175_));
 NOR2x1_ASAP7_75t_R _29064_ (.A(_01119_),
    .B(net277),
    .Y(_10111_));
 AO21x1_ASAP7_75t_R _29065_ (.A1(_08509_),
    .A2(net277),
    .B(_10111_),
    .Y(_03176_));
 NOR2x1_ASAP7_75t_R _29066_ (.A(_01153_),
    .B(net278),
    .Y(_10112_));
 AO21x1_ASAP7_75t_R _29067_ (.A1(_08537_),
    .A2(net278),
    .B(_10112_),
    .Y(_03177_));
 NOR2x1_ASAP7_75t_R _29068_ (.A(_01185_),
    .B(net278),
    .Y(_10113_));
 AO21x1_ASAP7_75t_R _29069_ (.A1(_08563_),
    .A2(net278),
    .B(_10113_),
    .Y(_03178_));
 NOR2x1_ASAP7_75t_R _29070_ (.A(_01219_),
    .B(net277),
    .Y(_10114_));
 AO21x1_ASAP7_75t_R _29071_ (.A1(net250),
    .A2(net277),
    .B(_10114_),
    .Y(_03179_));
 NOR2x1_ASAP7_75t_R _29072_ (.A(_01251_),
    .B(net278),
    .Y(_10115_));
 AO21x1_ASAP7_75t_R _29073_ (.A1(net2329),
    .A2(net278),
    .B(_10115_),
    .Y(_03180_));
 OR3x1_ASAP7_75t_R _29074_ (.A(_06985_),
    .B(_08648_),
    .C(_10077_),
    .Y(_10116_));
 OAI21x1_ASAP7_75t_R _29075_ (.A1(_01285_),
    .A2(net278),
    .B(_10116_),
    .Y(_03181_));
 NAND2x2_ASAP7_75t_R _29076_ (.A(_09756_),
    .B(_10036_),
    .Y(_10117_));
 TAPCELL_ASAP7_75t_R PHY_476 ();
 NOR2x1_ASAP7_75t_R _29078_ (.A(_07248_),
    .B(_10117_),
    .Y(_10119_));
 AO21x1_ASAP7_75t_R _29079_ (.A1(_13823_),
    .A2(_10117_),
    .B(_10119_),
    .Y(_03182_));
 AND2x6_ASAP7_75t_R _29080_ (.A(_09756_),
    .B(_10036_),
    .Y(_10120_));
 TAPCELL_ASAP7_75t_R PHY_475 ();
 AND2x2_ASAP7_75t_R _29082_ (.A(_13385_),
    .B(_10117_),
    .Y(_10122_));
 AO21x1_ASAP7_75t_R _29083_ (.A1(_07384_),
    .A2(_10120_),
    .B(_10122_),
    .Y(_03183_));
 AND2x2_ASAP7_75t_R _29084_ (.A(_14140_),
    .B(_10117_),
    .Y(_10123_));
 AO21x1_ASAP7_75t_R _29085_ (.A1(_07472_),
    .A2(_10120_),
    .B(_10123_),
    .Y(_03184_));
 AND2x2_ASAP7_75t_R _29086_ (.A(_14214_),
    .B(_10117_),
    .Y(_10124_));
 AO21x1_ASAP7_75t_R _29087_ (.A1(_07552_),
    .A2(_10120_),
    .B(_10124_),
    .Y(_03185_));
 AND2x2_ASAP7_75t_R _29088_ (.A(_15032_),
    .B(_10117_),
    .Y(_10125_));
 AO21x1_ASAP7_75t_R _29089_ (.A1(_07608_),
    .A2(_10120_),
    .B(_10125_),
    .Y(_03186_));
 AND2x2_ASAP7_75t_R _29090_ (.A(_14333_),
    .B(_10117_),
    .Y(_10126_));
 AO21x1_ASAP7_75t_R _29091_ (.A1(_07663_),
    .A2(_10120_),
    .B(_10126_),
    .Y(_03187_));
 AND2x2_ASAP7_75t_R _29092_ (.A(_14369_),
    .B(_10117_),
    .Y(_10127_));
 AO21x1_ASAP7_75t_R _29093_ (.A1(_07709_),
    .A2(_10120_),
    .B(_10127_),
    .Y(_03188_));
 TAPCELL_ASAP7_75t_R PHY_474 ();
 AND2x2_ASAP7_75t_R _29095_ (.A(_14428_),
    .B(_10117_),
    .Y(_10129_));
 AO21x1_ASAP7_75t_R _29096_ (.A1(net252),
    .A2(_10120_),
    .B(_10129_),
    .Y(_03189_));
 AND2x2_ASAP7_75t_R _29097_ (.A(_14490_),
    .B(_10117_),
    .Y(_10130_));
 AO21x1_ASAP7_75t_R _29098_ (.A1(net257),
    .A2(_10120_),
    .B(_10130_),
    .Y(_03190_));
 AND2x2_ASAP7_75t_R _29099_ (.A(_14552_),
    .B(_10117_),
    .Y(_10131_));
 AO21x1_ASAP7_75t_R _29100_ (.A1(net256),
    .A2(_10120_),
    .B(_10131_),
    .Y(_03191_));
 AND2x2_ASAP7_75t_R _29101_ (.A(_15377_),
    .B(_10117_),
    .Y(_10132_));
 AO21x1_ASAP7_75t_R _29102_ (.A1(_07903_),
    .A2(_10120_),
    .B(_10132_),
    .Y(_03192_));
 TAPCELL_ASAP7_75t_R PHY_473 ();
 AND2x2_ASAP7_75t_R _29104_ (.A(_14654_),
    .B(_10117_),
    .Y(_10134_));
 AO21x1_ASAP7_75t_R _29105_ (.A1(_07948_),
    .A2(_10120_),
    .B(_10134_),
    .Y(_03193_));
 AND2x2_ASAP7_75t_R _29106_ (.A(_14052_),
    .B(_10117_),
    .Y(_10135_));
 AO21x1_ASAP7_75t_R _29107_ (.A1(_07985_),
    .A2(_10120_),
    .B(_10135_),
    .Y(_03194_));
 AND2x2_ASAP7_75t_R _29108_ (.A(_15541_),
    .B(_10117_),
    .Y(_10136_));
 AO21x1_ASAP7_75t_R _29109_ (.A1(net251),
    .A2(_10120_),
    .B(_10136_),
    .Y(_03195_));
 AND2x2_ASAP7_75t_R _29110_ (.A(_15666_),
    .B(_10117_),
    .Y(_10137_));
 AO21x1_ASAP7_75t_R _29111_ (.A1(_08068_),
    .A2(_10120_),
    .B(_10137_),
    .Y(_03196_));
 TAPCELL_ASAP7_75t_R PHY_472 ();
 AND2x2_ASAP7_75t_R _29113_ (.A(_15787_),
    .B(_10117_),
    .Y(_10139_));
 AO21x1_ASAP7_75t_R _29114_ (.A1(_08110_),
    .A2(_10120_),
    .B(_10139_),
    .Y(_03197_));
 AND2x2_ASAP7_75t_R _29115_ (.A(_15904_),
    .B(_10117_),
    .Y(_10140_));
 AO21x1_ASAP7_75t_R _29116_ (.A1(_08151_),
    .A2(_10120_),
    .B(_10140_),
    .Y(_03198_));
 TAPCELL_ASAP7_75t_R PHY_471 ();
 AND2x2_ASAP7_75t_R _29118_ (.A(_16028_),
    .B(_10117_),
    .Y(_10142_));
 AO21x1_ASAP7_75t_R _29119_ (.A1(_08190_),
    .A2(_10120_),
    .B(_10142_),
    .Y(_03199_));
 AND2x2_ASAP7_75t_R _29120_ (.A(_16156_),
    .B(_10117_),
    .Y(_10143_));
 AO21x1_ASAP7_75t_R _29121_ (.A1(_08225_),
    .A2(_10120_),
    .B(_10143_),
    .Y(_03200_));
 AND2x2_ASAP7_75t_R _29122_ (.A(_16302_),
    .B(_10117_),
    .Y(_10144_));
 AO21x1_ASAP7_75t_R _29123_ (.A1(_08263_),
    .A2(_10120_),
    .B(_10144_),
    .Y(_03201_));
 AND2x2_ASAP7_75t_R _29124_ (.A(_16401_),
    .B(_10117_),
    .Y(_10145_));
 AO21x1_ASAP7_75t_R _29125_ (.A1(_08294_),
    .A2(_10120_),
    .B(_10145_),
    .Y(_03202_));
 TAPCELL_ASAP7_75t_R PHY_470 ();
 AND2x2_ASAP7_75t_R _29127_ (.A(_16516_),
    .B(_10117_),
    .Y(_10147_));
 AO21x1_ASAP7_75t_R _29128_ (.A1(_08328_),
    .A2(_10120_),
    .B(_10147_),
    .Y(_03203_));
 TAPCELL_ASAP7_75t_R PHY_469 ();
 AND2x2_ASAP7_75t_R _29130_ (.A(_16627_),
    .B(_10117_),
    .Y(_10149_));
 AO21x1_ASAP7_75t_R _29131_ (.A1(_08360_),
    .A2(_10120_),
    .B(_10149_),
    .Y(_03204_));
 AND2x2_ASAP7_75t_R _29132_ (.A(_04524_),
    .B(_10117_),
    .Y(_10150_));
 AO21x1_ASAP7_75t_R _29133_ (.A1(_08406_),
    .A2(_10120_),
    .B(_10150_),
    .Y(_03205_));
 TAPCELL_ASAP7_75t_R PHY_468 ();
 AND2x2_ASAP7_75t_R _29135_ (.A(_04644_),
    .B(_10117_),
    .Y(_10152_));
 AO21x1_ASAP7_75t_R _29136_ (.A1(_08450_),
    .A2(_10120_),
    .B(_10152_),
    .Y(_03206_));
 AND2x2_ASAP7_75t_R _29137_ (.A(_04756_),
    .B(_10117_),
    .Y(_10153_));
 AO21x1_ASAP7_75t_R _29138_ (.A1(_08481_),
    .A2(_10120_),
    .B(_10153_),
    .Y(_03207_));
 TAPCELL_ASAP7_75t_R PHY_467 ();
 AND2x2_ASAP7_75t_R _29140_ (.A(_04879_),
    .B(_10117_),
    .Y(_10155_));
 AO21x1_ASAP7_75t_R _29141_ (.A1(_08509_),
    .A2(_10120_),
    .B(_10155_),
    .Y(_03208_));
 AND2x2_ASAP7_75t_R _29142_ (.A(_04975_),
    .B(_10117_),
    .Y(_10156_));
 AO21x1_ASAP7_75t_R _29143_ (.A1(_08537_),
    .A2(_10120_),
    .B(_10156_),
    .Y(_03209_));
 AND2x2_ASAP7_75t_R _29144_ (.A(_05084_),
    .B(_10117_),
    .Y(_10157_));
 AO21x1_ASAP7_75t_R _29145_ (.A1(_08563_),
    .A2(_10120_),
    .B(_10157_),
    .Y(_03210_));
 AND2x2_ASAP7_75t_R _29146_ (.A(_05192_),
    .B(_10117_),
    .Y(_10158_));
 AO21x1_ASAP7_75t_R _29147_ (.A1(net250),
    .A2(_10120_),
    .B(_10158_),
    .Y(_03211_));
 TAPCELL_ASAP7_75t_R PHY_466 ();
 AND2x2_ASAP7_75t_R _29149_ (.A(_05298_),
    .B(_10117_),
    .Y(_10160_));
 AO21x1_ASAP7_75t_R _29150_ (.A1(net2329),
    .A2(_10120_),
    .B(_10160_),
    .Y(_03212_));
 NOR2x1_ASAP7_75t_R _29151_ (.A(_08648_),
    .B(_10117_),
    .Y(_10161_));
 AO21x1_ASAP7_75t_R _29152_ (.A1(_05426_),
    .A2(_10117_),
    .B(_10161_),
    .Y(_03213_));
 NOR2x2_ASAP7_75t_R _29153_ (.A(_09829_),
    .B(_10077_),
    .Y(_10162_));
 TAPCELL_ASAP7_75t_R PHY_465 ();
 TAPCELL_ASAP7_75t_R PHY_464 ();
 NAND2x1_ASAP7_75t_R _29156_ (.A(_07248_),
    .B(net276),
    .Y(_10165_));
 OA21x2_ASAP7_75t_R _29157_ (.A1(_13828_),
    .A2(net276),
    .B(_10165_),
    .Y(_03214_));
 TAPCELL_ASAP7_75t_R PHY_463 ();
 NOR2x1_ASAP7_75t_R _29159_ (.A(_00256_),
    .B(net276),
    .Y(_10167_));
 AO21x1_ASAP7_75t_R _29160_ (.A1(_07384_),
    .A2(net276),
    .B(_10167_),
    .Y(_03215_));
 NOR2x1_ASAP7_75t_R _29161_ (.A(_00364_),
    .B(net275),
    .Y(_10168_));
 AO21x1_ASAP7_75t_R _29162_ (.A1(_07472_),
    .A2(net275),
    .B(_10168_),
    .Y(_03216_));
 NOR2x1_ASAP7_75t_R _29163_ (.A(_00395_),
    .B(net276),
    .Y(_10169_));
 AO21x1_ASAP7_75t_R _29164_ (.A1(_07552_),
    .A2(net276),
    .B(_10169_),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _29165_ (.A(_00425_),
    .B(net275),
    .Y(_10170_));
 AO21x1_ASAP7_75t_R _29166_ (.A1(_07608_),
    .A2(net275),
    .B(_10170_),
    .Y(_03218_));
 TAPCELL_ASAP7_75t_R PHY_462 ();
 NOR2x1_ASAP7_75t_R _29168_ (.A(_00455_),
    .B(net275),
    .Y(_10172_));
 AO21x1_ASAP7_75t_R _29169_ (.A1(_07663_),
    .A2(net275),
    .B(_10172_),
    .Y(_03219_));
 NOR2x1_ASAP7_75t_R _29170_ (.A(_00485_),
    .B(net275),
    .Y(_10173_));
 AO21x1_ASAP7_75t_R _29171_ (.A1(_07709_),
    .A2(net275),
    .B(_10173_),
    .Y(_03220_));
 TAPCELL_ASAP7_75t_R PHY_461 ();
 NOR2x1_ASAP7_75t_R _29173_ (.A(_00515_),
    .B(_10162_),
    .Y(_10175_));
 AO21x1_ASAP7_75t_R _29174_ (.A1(net252),
    .A2(_10162_),
    .B(_10175_),
    .Y(_03221_));
 TAPCELL_ASAP7_75t_R PHY_460 ();
 NOR2x1_ASAP7_75t_R _29176_ (.A(_00545_),
    .B(_10162_),
    .Y(_10177_));
 AO21x1_ASAP7_75t_R _29177_ (.A1(net257),
    .A2(_10162_),
    .B(_10177_),
    .Y(_03222_));
 TAPCELL_ASAP7_75t_R PHY_459 ();
 NOR2x1_ASAP7_75t_R _29179_ (.A(_00575_),
    .B(net276),
    .Y(_10179_));
 AO21x1_ASAP7_75t_R _29180_ (.A1(net256),
    .A2(net276),
    .B(_10179_),
    .Y(_03223_));
 NOR2x1_ASAP7_75t_R _29181_ (.A(_00605_),
    .B(net275),
    .Y(_10180_));
 AO21x1_ASAP7_75t_R _29182_ (.A1(_07903_),
    .A2(net275),
    .B(_10180_),
    .Y(_03224_));
 NOR2x1_ASAP7_75t_R _29183_ (.A(_00635_),
    .B(net275),
    .Y(_10181_));
 AO21x1_ASAP7_75t_R _29184_ (.A1(_07948_),
    .A2(net275),
    .B(_10181_),
    .Y(_03225_));
 TAPCELL_ASAP7_75t_R PHY_458 ();
 NOR2x1_ASAP7_75t_R _29186_ (.A(_00334_),
    .B(net275),
    .Y(_10183_));
 AO21x1_ASAP7_75t_R _29187_ (.A1(_07985_),
    .A2(net275),
    .B(_10183_),
    .Y(_03226_));
 TAPCELL_ASAP7_75t_R PHY_457 ();
 NOR2x1_ASAP7_75t_R _29189_ (.A(_00697_),
    .B(net276),
    .Y(_10185_));
 AO21x1_ASAP7_75t_R _29190_ (.A1(net251),
    .A2(net276),
    .B(_10185_),
    .Y(_03227_));
 NOR2x1_ASAP7_75t_R _29191_ (.A(_00729_),
    .B(net275),
    .Y(_10186_));
 AO21x1_ASAP7_75t_R _29192_ (.A1(_08068_),
    .A2(net275),
    .B(_10186_),
    .Y(_03228_));
 NOR2x1_ASAP7_75t_R _29193_ (.A(_00762_),
    .B(net276),
    .Y(_10187_));
 AO21x1_ASAP7_75t_R _29194_ (.A1(_08110_),
    .A2(net276),
    .B(_10187_),
    .Y(_03229_));
 TAPCELL_ASAP7_75t_R PHY_456 ();
 NOR2x1_ASAP7_75t_R _29196_ (.A(_00795_),
    .B(net275),
    .Y(_10189_));
 AO21x1_ASAP7_75t_R _29197_ (.A1(_08151_),
    .A2(net275),
    .B(_10189_),
    .Y(_03230_));
 TAPCELL_ASAP7_75t_R PHY_455 ();
 NOR2x1_ASAP7_75t_R _29199_ (.A(_00828_),
    .B(net275),
    .Y(_10191_));
 AO21x1_ASAP7_75t_R _29200_ (.A1(_08190_),
    .A2(net275),
    .B(_10191_),
    .Y(_03231_));
 TAPCELL_ASAP7_75t_R PHY_454 ();
 NOR2x1_ASAP7_75t_R _29202_ (.A(_00860_),
    .B(net276),
    .Y(_10193_));
 AO21x1_ASAP7_75t_R _29203_ (.A1(_08225_),
    .A2(net276),
    .B(_10193_),
    .Y(_03232_));
 TAPCELL_ASAP7_75t_R PHY_453 ();
 NOR2x1_ASAP7_75t_R _29205_ (.A(_00893_),
    .B(net275),
    .Y(_10195_));
 AO21x1_ASAP7_75t_R _29206_ (.A1(_08263_),
    .A2(net275),
    .B(_10195_),
    .Y(_03233_));
 TAPCELL_ASAP7_75t_R PHY_452 ();
 NOR2x1_ASAP7_75t_R _29208_ (.A(_00925_),
    .B(net276),
    .Y(_10197_));
 AO21x1_ASAP7_75t_R _29209_ (.A1(_08294_),
    .A2(net276),
    .B(_10197_),
    .Y(_03234_));
 NOR2x1_ASAP7_75t_R _29210_ (.A(_00958_),
    .B(net275),
    .Y(_10198_));
 AO21x1_ASAP7_75t_R _29211_ (.A1(_08328_),
    .A2(net275),
    .B(_10198_),
    .Y(_03235_));
 NOR2x1_ASAP7_75t_R _29212_ (.A(_00990_),
    .B(net276),
    .Y(_10199_));
 AO21x1_ASAP7_75t_R _29213_ (.A1(_08360_),
    .A2(net276),
    .B(_10199_),
    .Y(_03236_));
 TAPCELL_ASAP7_75t_R PHY_451 ();
 NOR2x1_ASAP7_75t_R _29215_ (.A(_01024_),
    .B(net276),
    .Y(_10201_));
 AO21x1_ASAP7_75t_R _29216_ (.A1(_08406_),
    .A2(net276),
    .B(_10201_),
    .Y(_03237_));
 NOR2x1_ASAP7_75t_R _29217_ (.A(_01056_),
    .B(net276),
    .Y(_10202_));
 AO21x1_ASAP7_75t_R _29218_ (.A1(_08450_),
    .A2(net276),
    .B(_10202_),
    .Y(_03238_));
 NOR2x1_ASAP7_75t_R _29219_ (.A(_01089_),
    .B(net275),
    .Y(_10203_));
 AO21x1_ASAP7_75t_R _29220_ (.A1(_08481_),
    .A2(net275),
    .B(_10203_),
    .Y(_03239_));
 NOR2x1_ASAP7_75t_R _29221_ (.A(_01121_),
    .B(net275),
    .Y(_10204_));
 AO21x1_ASAP7_75t_R _29222_ (.A1(_08509_),
    .A2(net275),
    .B(_10204_),
    .Y(_03240_));
 NOR2x1_ASAP7_75t_R _29223_ (.A(_01155_),
    .B(_10162_),
    .Y(_10205_));
 AO21x1_ASAP7_75t_R _29224_ (.A1(_08537_),
    .A2(_10162_),
    .B(_10205_),
    .Y(_03241_));
 TAPCELL_ASAP7_75t_R PHY_450 ();
 NOR2x1_ASAP7_75t_R _29226_ (.A(_01187_),
    .B(_10162_),
    .Y(_10207_));
 AO21x1_ASAP7_75t_R _29227_ (.A1(_08563_),
    .A2(_10162_),
    .B(_10207_),
    .Y(_03242_));
 TAPCELL_ASAP7_75t_R PHY_449 ();
 NOR2x1_ASAP7_75t_R _29229_ (.A(_01221_),
    .B(net275),
    .Y(_10209_));
 AO21x1_ASAP7_75t_R _29230_ (.A1(net250),
    .A2(net275),
    .B(_10209_),
    .Y(_03243_));
 NOR2x1_ASAP7_75t_R _29231_ (.A(_01253_),
    .B(net276),
    .Y(_10210_));
 AO21x1_ASAP7_75t_R _29232_ (.A1(net2329),
    .A2(net276),
    .B(_10210_),
    .Y(_03244_));
 NAND2x1_ASAP7_75t_R _29233_ (.A(_08648_),
    .B(_10162_),
    .Y(_10211_));
 OA21x2_ASAP7_75t_R _29234_ (.A1(_05423_),
    .A2(_10162_),
    .B(_10211_),
    .Y(_03245_));
 INVx1_ASAP7_75t_R _29235_ (.A(_00303_),
    .Y(_10212_));
 NOR2x2_ASAP7_75t_R _29236_ (.A(_00187_),
    .B(_00191_),
    .Y(_10213_));
 AND4x2_ASAP7_75t_R _29237_ (.A(_00184_),
    .B(_00194_),
    .C(_09871_),
    .D(_10213_),
    .Y(_10214_));
 TAPCELL_ASAP7_75t_R PHY_448 ();
 TAPCELL_ASAP7_75t_R PHY_447 ();
 TAPCELL_ASAP7_75t_R PHY_446 ();
 NAND2x1_ASAP7_75t_R _29241_ (.A(_07248_),
    .B(_10214_),
    .Y(_10218_));
 OA21x2_ASAP7_75t_R _29242_ (.A1(_10212_),
    .A2(_10214_),
    .B(_10218_),
    .Y(_03246_));
 NOR2x1_ASAP7_75t_R _29243_ (.A(_00257_),
    .B(net274),
    .Y(_10219_));
 AO21x1_ASAP7_75t_R _29244_ (.A1(_07384_),
    .A2(net274),
    .B(_10219_),
    .Y(_03247_));
 TAPCELL_ASAP7_75t_R PHY_445 ();
 NOR2x1_ASAP7_75t_R _29246_ (.A(_00365_),
    .B(net273),
    .Y(_10221_));
 AO21x1_ASAP7_75t_R _29247_ (.A1(_07472_),
    .A2(net273),
    .B(_10221_),
    .Y(_03248_));
 TAPCELL_ASAP7_75t_R PHY_444 ();
 NOR2x1_ASAP7_75t_R _29249_ (.A(_00396_),
    .B(_10214_),
    .Y(_10223_));
 AO21x1_ASAP7_75t_R _29250_ (.A1(_07552_),
    .A2(_10214_),
    .B(_10223_),
    .Y(_03249_));
 TAPCELL_ASAP7_75t_R PHY_443 ();
 NOR2x1_ASAP7_75t_R _29252_ (.A(_00426_),
    .B(net273),
    .Y(_10225_));
 AO21x1_ASAP7_75t_R _29253_ (.A1(_07608_),
    .A2(net273),
    .B(_10225_),
    .Y(_03250_));
 NOR2x1_ASAP7_75t_R _29254_ (.A(_00456_),
    .B(net273),
    .Y(_10226_));
 AO21x1_ASAP7_75t_R _29255_ (.A1(_07663_),
    .A2(net273),
    .B(_10226_),
    .Y(_03251_));
 TAPCELL_ASAP7_75t_R PHY_442 ();
 NOR2x1_ASAP7_75t_R _29257_ (.A(_00486_),
    .B(net273),
    .Y(_10228_));
 AO21x1_ASAP7_75t_R _29258_ (.A1(_07709_),
    .A2(net273),
    .B(_10228_),
    .Y(_03252_));
 TAPCELL_ASAP7_75t_R PHY_441 ();
 TAPCELL_ASAP7_75t_R PHY_440 ();
 NOR2x1_ASAP7_75t_R _29261_ (.A(_00516_),
    .B(net274),
    .Y(_10231_));
 AO21x1_ASAP7_75t_R _29262_ (.A1(net252),
    .A2(net274),
    .B(_10231_),
    .Y(_03253_));
 NOR2x1_ASAP7_75t_R _29263_ (.A(_00546_),
    .B(net274),
    .Y(_10232_));
 AO21x1_ASAP7_75t_R _29264_ (.A1(net257),
    .A2(net274),
    .B(_10232_),
    .Y(_03254_));
 TAPCELL_ASAP7_75t_R PHY_439 ();
 TAPCELL_ASAP7_75t_R PHY_438 ();
 NOR2x1_ASAP7_75t_R _29267_ (.A(_00576_),
    .B(_10214_),
    .Y(_10235_));
 AO21x1_ASAP7_75t_R _29268_ (.A1(net256),
    .A2(_10214_),
    .B(_10235_),
    .Y(_03255_));
 TAPCELL_ASAP7_75t_R PHY_437 ();
 NOR2x1_ASAP7_75t_R _29270_ (.A(_00606_),
    .B(net273),
    .Y(_10237_));
 AO21x1_ASAP7_75t_R _29271_ (.A1(_07903_),
    .A2(net273),
    .B(_10237_),
    .Y(_03256_));
 TAPCELL_ASAP7_75t_R PHY_436 ();
 NOR2x1_ASAP7_75t_R _29273_ (.A(_00636_),
    .B(net273),
    .Y(_10239_));
 AO21x1_ASAP7_75t_R _29274_ (.A1(_07948_),
    .A2(net273),
    .B(_10239_),
    .Y(_03257_));
 NOR2x1_ASAP7_75t_R _29275_ (.A(_00335_),
    .B(net273),
    .Y(_10240_));
 AO21x1_ASAP7_75t_R _29276_ (.A1(_07985_),
    .A2(net273),
    .B(_10240_),
    .Y(_03258_));
 NOR2x1_ASAP7_75t_R _29277_ (.A(_00698_),
    .B(net274),
    .Y(_10241_));
 AO21x1_ASAP7_75t_R _29278_ (.A1(_08026_),
    .A2(net274),
    .B(_10241_),
    .Y(_03259_));
 TAPCELL_ASAP7_75t_R PHY_435 ();
 NOR2x1_ASAP7_75t_R _29280_ (.A(_00730_),
    .B(net274),
    .Y(_10243_));
 AO21x1_ASAP7_75t_R _29281_ (.A1(_08068_),
    .A2(net274),
    .B(_10243_),
    .Y(_03260_));
 NOR2x1_ASAP7_75t_R _29282_ (.A(_00763_),
    .B(_10214_),
    .Y(_10244_));
 AO21x1_ASAP7_75t_R _29283_ (.A1(_08110_),
    .A2(_10214_),
    .B(_10244_),
    .Y(_03261_));
 NOR2x1_ASAP7_75t_R _29284_ (.A(_00796_),
    .B(net273),
    .Y(_10245_));
 AO21x1_ASAP7_75t_R _29285_ (.A1(_08151_),
    .A2(net273),
    .B(_10245_),
    .Y(_03262_));
 TAPCELL_ASAP7_75t_R PHY_434 ();
 TAPCELL_ASAP7_75t_R PHY_433 ();
 NOR2x1_ASAP7_75t_R _29288_ (.A(_00829_),
    .B(net273),
    .Y(_10248_));
 AO21x1_ASAP7_75t_R _29289_ (.A1(_08190_),
    .A2(net273),
    .B(_10248_),
    .Y(_03263_));
 NOR2x1_ASAP7_75t_R _29290_ (.A(_00861_),
    .B(_10214_),
    .Y(_10249_));
 AO21x1_ASAP7_75t_R _29291_ (.A1(_08225_),
    .A2(_10214_),
    .B(_10249_),
    .Y(_03264_));
 TAPCELL_ASAP7_75t_R PHY_432 ();
 TAPCELL_ASAP7_75t_R PHY_431 ();
 NOR2x1_ASAP7_75t_R _29294_ (.A(_00894_),
    .B(net273),
    .Y(_10252_));
 AO21x1_ASAP7_75t_R _29295_ (.A1(_08263_),
    .A2(net273),
    .B(_10252_),
    .Y(_03265_));
 NOR2x1_ASAP7_75t_R _29296_ (.A(_00926_),
    .B(_10214_),
    .Y(_10253_));
 AO21x1_ASAP7_75t_R _29297_ (.A1(_08294_),
    .A2(_10214_),
    .B(_10253_),
    .Y(_03266_));
 TAPCELL_ASAP7_75t_R PHY_430 ();
 NOR2x1_ASAP7_75t_R _29299_ (.A(_00959_),
    .B(net273),
    .Y(_10255_));
 AO21x1_ASAP7_75t_R _29300_ (.A1(_08328_),
    .A2(net273),
    .B(_10255_),
    .Y(_03267_));
 NOR2x1_ASAP7_75t_R _29301_ (.A(_00991_),
    .B(_10214_),
    .Y(_10256_));
 AO21x1_ASAP7_75t_R _29302_ (.A1(_08360_),
    .A2(_10214_),
    .B(_10256_),
    .Y(_03268_));
 NOR2x1_ASAP7_75t_R _29303_ (.A(_01025_),
    .B(net274),
    .Y(_10257_));
 AO21x1_ASAP7_75t_R _29304_ (.A1(_08406_),
    .A2(net274),
    .B(_10257_),
    .Y(_03269_));
 NOR2x1_ASAP7_75t_R _29305_ (.A(_01057_),
    .B(_10214_),
    .Y(_10258_));
 AO21x1_ASAP7_75t_R _29306_ (.A1(_08450_),
    .A2(_10214_),
    .B(_10258_),
    .Y(_03270_));
 TAPCELL_ASAP7_75t_R PHY_429 ();
 NOR2x1_ASAP7_75t_R _29308_ (.A(_01090_),
    .B(net273),
    .Y(_10260_));
 AO21x1_ASAP7_75t_R _29309_ (.A1(_08481_),
    .A2(net273),
    .B(_10260_),
    .Y(_03271_));
 NOR2x1_ASAP7_75t_R _29310_ (.A(_01122_),
    .B(net274),
    .Y(_10261_));
 AO21x1_ASAP7_75t_R _29311_ (.A1(_08509_),
    .A2(net274),
    .B(_10261_),
    .Y(_03272_));
 TAPCELL_ASAP7_75t_R PHY_428 ();
 NOR2x1_ASAP7_75t_R _29313_ (.A(_01156_),
    .B(net274),
    .Y(_10263_));
 AO21x1_ASAP7_75t_R _29314_ (.A1(_08537_),
    .A2(net274),
    .B(_10263_),
    .Y(_03273_));
 NOR2x1_ASAP7_75t_R _29315_ (.A(_01188_),
    .B(net274),
    .Y(_10264_));
 AO21x1_ASAP7_75t_R _29316_ (.A1(_08563_),
    .A2(net274),
    .B(_10264_),
    .Y(_03274_));
 NOR2x1_ASAP7_75t_R _29317_ (.A(_01222_),
    .B(net273),
    .Y(_10265_));
 AO21x1_ASAP7_75t_R _29318_ (.A1(net250),
    .A2(net273),
    .B(_10265_),
    .Y(_03275_));
 NOR2x1_ASAP7_75t_R _29319_ (.A(_01254_),
    .B(net274),
    .Y(_10266_));
 AO21x1_ASAP7_75t_R _29320_ (.A1(net2330),
    .A2(net274),
    .B(_10266_),
    .Y(_03276_));
 NAND2x1_ASAP7_75t_R _29321_ (.A(_08648_),
    .B(net274),
    .Y(_10267_));
 OA21x2_ASAP7_75t_R _29322_ (.A1(_05420_),
    .A2(net274),
    .B(_10267_),
    .Y(_03277_));
 INVx1_ASAP7_75t_R _29323_ (.A(_00304_),
    .Y(_10268_));
 OR2x6_ASAP7_75t_R _29324_ (.A(_00187_),
    .B(_00191_),
    .Y(_10269_));
 TAPCELL_ASAP7_75t_R PHY_427 ();
 NOR2x2_ASAP7_75t_R _29326_ (.A(_06985_),
    .B(_10269_),
    .Y(_10271_));
 TAPCELL_ASAP7_75t_R PHY_426 ();
 TAPCELL_ASAP7_75t_R PHY_425 ();
 NAND2x1_ASAP7_75t_R _29329_ (.A(_07248_),
    .B(_10271_),
    .Y(_10274_));
 OA21x2_ASAP7_75t_R _29330_ (.A1(_10268_),
    .A2(_10271_),
    .B(_10274_),
    .Y(_03278_));
 NOR2x1_ASAP7_75t_R _29331_ (.A(_00258_),
    .B(_10271_),
    .Y(_10275_));
 AO21x1_ASAP7_75t_R _29332_ (.A1(_07384_),
    .A2(_10271_),
    .B(_10275_),
    .Y(_03279_));
 NOR2x1_ASAP7_75t_R _29333_ (.A(_00366_),
    .B(net271),
    .Y(_10276_));
 AO21x1_ASAP7_75t_R _29334_ (.A1(_07472_),
    .A2(net271),
    .B(_10276_),
    .Y(_03280_));
 NOR2x1_ASAP7_75t_R _29335_ (.A(_00397_),
    .B(_10271_),
    .Y(_10277_));
 AO21x1_ASAP7_75t_R _29336_ (.A1(_07552_),
    .A2(_10271_),
    .B(_10277_),
    .Y(_03281_));
 NOR2x1_ASAP7_75t_R _29337_ (.A(_00427_),
    .B(net271),
    .Y(_10278_));
 AO21x1_ASAP7_75t_R _29338_ (.A1(_07608_),
    .A2(net271),
    .B(_10278_),
    .Y(_03282_));
 NOR2x1_ASAP7_75t_R _29339_ (.A(_00457_),
    .B(net271),
    .Y(_10279_));
 AO21x1_ASAP7_75t_R _29340_ (.A1(_07663_),
    .A2(net271),
    .B(_10279_),
    .Y(_03283_));
 NOR2x1_ASAP7_75t_R _29341_ (.A(_00487_),
    .B(net271),
    .Y(_10280_));
 AO21x1_ASAP7_75t_R _29342_ (.A1(_07709_),
    .A2(net271),
    .B(_10280_),
    .Y(_03284_));
 TAPCELL_ASAP7_75t_R PHY_424 ();
 NOR2x1_ASAP7_75t_R _29344_ (.A(_00517_),
    .B(net272),
    .Y(_10282_));
 AO21x1_ASAP7_75t_R _29345_ (.A1(net252),
    .A2(net272),
    .B(_10282_),
    .Y(_03285_));
 NOR2x1_ASAP7_75t_R _29346_ (.A(_00547_),
    .B(net272),
    .Y(_10283_));
 AO21x1_ASAP7_75t_R _29347_ (.A1(net257),
    .A2(net272),
    .B(_10283_),
    .Y(_03286_));
 TAPCELL_ASAP7_75t_R PHY_423 ();
 NOR2x1_ASAP7_75t_R _29349_ (.A(_00577_),
    .B(_10271_),
    .Y(_10285_));
 AO21x1_ASAP7_75t_R _29350_ (.A1(net256),
    .A2(_10271_),
    .B(_10285_),
    .Y(_03287_));
 NOR2x1_ASAP7_75t_R _29351_ (.A(_00607_),
    .B(net271),
    .Y(_10286_));
 AO21x1_ASAP7_75t_R _29352_ (.A1(_07903_),
    .A2(net271),
    .B(_10286_),
    .Y(_03288_));
 NOR2x1_ASAP7_75t_R _29353_ (.A(_00637_),
    .B(net271),
    .Y(_10287_));
 AO21x1_ASAP7_75t_R _29354_ (.A1(_07948_),
    .A2(net271),
    .B(_10287_),
    .Y(_03289_));
 NOR2x1_ASAP7_75t_R _29355_ (.A(_00336_),
    .B(net271),
    .Y(_10288_));
 AO21x1_ASAP7_75t_R _29356_ (.A1(_07985_),
    .A2(net271),
    .B(_10288_),
    .Y(_03290_));
 NOR2x1_ASAP7_75t_R _29357_ (.A(_00699_),
    .B(_10271_),
    .Y(_10289_));
 AO21x1_ASAP7_75t_R _29358_ (.A1(_08026_),
    .A2(_10271_),
    .B(_10289_),
    .Y(_03291_));
 NOR2x1_ASAP7_75t_R _29359_ (.A(_00731_),
    .B(net272),
    .Y(_10290_));
 AO21x1_ASAP7_75t_R _29360_ (.A1(_08068_),
    .A2(net272),
    .B(_10290_),
    .Y(_03292_));
 NOR2x1_ASAP7_75t_R _29361_ (.A(_00764_),
    .B(_10271_),
    .Y(_10291_));
 AO21x1_ASAP7_75t_R _29362_ (.A1(_08110_),
    .A2(_10271_),
    .B(_10291_),
    .Y(_03293_));
 NOR2x1_ASAP7_75t_R _29363_ (.A(_00797_),
    .B(net272),
    .Y(_10292_));
 AO21x1_ASAP7_75t_R _29364_ (.A1(_08151_),
    .A2(net272),
    .B(_10292_),
    .Y(_03294_));
 TAPCELL_ASAP7_75t_R PHY_422 ();
 NOR2x1_ASAP7_75t_R _29366_ (.A(_00830_),
    .B(net271),
    .Y(_10294_));
 AO21x1_ASAP7_75t_R _29367_ (.A1(_08190_),
    .A2(net271),
    .B(_10294_),
    .Y(_03295_));
 NOR2x1_ASAP7_75t_R _29368_ (.A(_00862_),
    .B(_10271_),
    .Y(_10295_));
 AO21x1_ASAP7_75t_R _29369_ (.A1(_08225_),
    .A2(_10271_),
    .B(_10295_),
    .Y(_03296_));
 TAPCELL_ASAP7_75t_R PHY_421 ();
 NOR2x1_ASAP7_75t_R _29371_ (.A(_00895_),
    .B(net271),
    .Y(_10297_));
 AO21x1_ASAP7_75t_R _29372_ (.A1(_08263_),
    .A2(net271),
    .B(_10297_),
    .Y(_03297_));
 NOR2x1_ASAP7_75t_R _29373_ (.A(_00927_),
    .B(_10271_),
    .Y(_10298_));
 AO21x1_ASAP7_75t_R _29374_ (.A1(_08294_),
    .A2(_10271_),
    .B(_10298_),
    .Y(_03298_));
 NOR2x1_ASAP7_75t_R _29375_ (.A(_00960_),
    .B(net271),
    .Y(_10299_));
 AO21x1_ASAP7_75t_R _29376_ (.A1(_08328_),
    .A2(net271),
    .B(_10299_),
    .Y(_03299_));
 NOR2x1_ASAP7_75t_R _29377_ (.A(_00992_),
    .B(_10271_),
    .Y(_10300_));
 AO21x1_ASAP7_75t_R _29378_ (.A1(_08360_),
    .A2(_10271_),
    .B(_10300_),
    .Y(_03300_));
 NOR2x1_ASAP7_75t_R _29379_ (.A(_01026_),
    .B(net272),
    .Y(_10301_));
 AO21x1_ASAP7_75t_R _29380_ (.A1(_08406_),
    .A2(net272),
    .B(_10301_),
    .Y(_03301_));
 NOR2x1_ASAP7_75t_R _29381_ (.A(_01058_),
    .B(_10271_),
    .Y(_10302_));
 AO21x1_ASAP7_75t_R _29382_ (.A1(_08450_),
    .A2(_10271_),
    .B(_10302_),
    .Y(_03302_));
 NOR2x1_ASAP7_75t_R _29383_ (.A(_01091_),
    .B(net271),
    .Y(_10303_));
 AO21x1_ASAP7_75t_R _29384_ (.A1(_08481_),
    .A2(net271),
    .B(_10303_),
    .Y(_03303_));
 NOR2x1_ASAP7_75t_R _29385_ (.A(_01123_),
    .B(net272),
    .Y(_10304_));
 AO21x1_ASAP7_75t_R _29386_ (.A1(_08509_),
    .A2(net272),
    .B(_10304_),
    .Y(_03304_));
 NOR2x1_ASAP7_75t_R _29387_ (.A(_01157_),
    .B(net272),
    .Y(_10305_));
 AO21x1_ASAP7_75t_R _29388_ (.A1(_08537_),
    .A2(net272),
    .B(_10305_),
    .Y(_03305_));
 NOR2x1_ASAP7_75t_R _29389_ (.A(_01189_),
    .B(_10271_),
    .Y(_10306_));
 AO21x1_ASAP7_75t_R _29390_ (.A1(_08563_),
    .A2(_10271_),
    .B(_10306_),
    .Y(_03306_));
 NOR2x1_ASAP7_75t_R _29391_ (.A(_01223_),
    .B(net271),
    .Y(_10307_));
 AO21x1_ASAP7_75t_R _29392_ (.A1(net250),
    .A2(net271),
    .B(_10307_),
    .Y(_03307_));
 NOR2x1_ASAP7_75t_R _29393_ (.A(_01255_),
    .B(_10271_),
    .Y(_10308_));
 AO21x1_ASAP7_75t_R _29394_ (.A1(net2198),
    .A2(_10271_),
    .B(_10308_),
    .Y(_03308_));
 NAND2x1_ASAP7_75t_R _29395_ (.A(_08648_),
    .B(net272),
    .Y(_10309_));
 OA21x2_ASAP7_75t_R _29396_ (.A1(_05460_),
    .A2(net272),
    .B(_10309_),
    .Y(_03309_));
 AND2x6_ASAP7_75t_R _29397_ (.A(_09756_),
    .B(_10213_),
    .Y(_10310_));
 TAPCELL_ASAP7_75t_R PHY_420 ();
 TAPCELL_ASAP7_75t_R PHY_419 ();
 TAPCELL_ASAP7_75t_R PHY_418 ();
 NAND2x1_ASAP7_75t_R _29401_ (.A(_07248_),
    .B(_10310_),
    .Y(_10314_));
 OA21x2_ASAP7_75t_R _29402_ (.A1(_13833_),
    .A2(_10310_),
    .B(_10314_),
    .Y(_03310_));
 NOR2x1_ASAP7_75t_R _29403_ (.A(_00259_),
    .B(_10310_),
    .Y(_10315_));
 AO21x1_ASAP7_75t_R _29404_ (.A1(_07384_),
    .A2(_10310_),
    .B(_10315_),
    .Y(_03311_));
 NOR2x1_ASAP7_75t_R _29405_ (.A(_00367_),
    .B(_10310_),
    .Y(_10316_));
 AO21x1_ASAP7_75t_R _29406_ (.A1(_07472_),
    .A2(_10310_),
    .B(_10316_),
    .Y(_03312_));
 NOR2x1_ASAP7_75t_R _29407_ (.A(_00398_),
    .B(_10310_),
    .Y(_10317_));
 AO21x1_ASAP7_75t_R _29408_ (.A1(_07552_),
    .A2(_10310_),
    .B(_10317_),
    .Y(_03313_));
 NOR2x1_ASAP7_75t_R _29409_ (.A(_00428_),
    .B(_10310_),
    .Y(_10318_));
 AO21x1_ASAP7_75t_R _29410_ (.A1(_07608_),
    .A2(_10310_),
    .B(_10318_),
    .Y(_03314_));
 NOR2x1_ASAP7_75t_R _29411_ (.A(_00458_),
    .B(_10310_),
    .Y(_10319_));
 AO21x1_ASAP7_75t_R _29412_ (.A1(_07663_),
    .A2(_10310_),
    .B(_10319_),
    .Y(_03315_));
 NOR2x1_ASAP7_75t_R _29413_ (.A(_00488_),
    .B(_10310_),
    .Y(_10320_));
 AO21x1_ASAP7_75t_R _29414_ (.A1(_07709_),
    .A2(_10310_),
    .B(_10320_),
    .Y(_03316_));
 TAPCELL_ASAP7_75t_R PHY_417 ();
 NOR2x1_ASAP7_75t_R _29416_ (.A(_00518_),
    .B(_10310_),
    .Y(_10322_));
 AO21x1_ASAP7_75t_R _29417_ (.A1(net252),
    .A2(_10310_),
    .B(_10322_),
    .Y(_03317_));
 NOR2x1_ASAP7_75t_R _29418_ (.A(_00548_),
    .B(_10310_),
    .Y(_10323_));
 AO21x1_ASAP7_75t_R _29419_ (.A1(net257),
    .A2(_10310_),
    .B(_10323_),
    .Y(_03318_));
 TAPCELL_ASAP7_75t_R PHY_416 ();
 NOR2x1_ASAP7_75t_R _29421_ (.A(_00578_),
    .B(_10310_),
    .Y(_10325_));
 AO21x1_ASAP7_75t_R _29422_ (.A1(net256),
    .A2(_10310_),
    .B(_10325_),
    .Y(_03319_));
 NOR2x1_ASAP7_75t_R _29423_ (.A(_00608_),
    .B(_10310_),
    .Y(_10326_));
 AO21x1_ASAP7_75t_R _29424_ (.A1(_07903_),
    .A2(_10310_),
    .B(_10326_),
    .Y(_03320_));
 NOR2x1_ASAP7_75t_R _29425_ (.A(_00638_),
    .B(_10310_),
    .Y(_10327_));
 AO21x1_ASAP7_75t_R _29426_ (.A1(_07948_),
    .A2(_10310_),
    .B(_10327_),
    .Y(_03321_));
 NOR2x1_ASAP7_75t_R _29427_ (.A(_00337_),
    .B(_10310_),
    .Y(_10328_));
 AO21x1_ASAP7_75t_R _29428_ (.A1(_07985_),
    .A2(_10310_),
    .B(_10328_),
    .Y(_03322_));
 NOR2x1_ASAP7_75t_R _29429_ (.A(_00700_),
    .B(_10310_),
    .Y(_10329_));
 AO21x1_ASAP7_75t_R _29430_ (.A1(_08026_),
    .A2(_10310_),
    .B(_10329_),
    .Y(_03323_));
 NOR2x1_ASAP7_75t_R _29431_ (.A(_00732_),
    .B(_10310_),
    .Y(_10330_));
 AO21x1_ASAP7_75t_R _29432_ (.A1(_08068_),
    .A2(_10310_),
    .B(_10330_),
    .Y(_03324_));
 NOR2x1_ASAP7_75t_R _29433_ (.A(_00765_),
    .B(_10310_),
    .Y(_10331_));
 AO21x1_ASAP7_75t_R _29434_ (.A1(_08110_),
    .A2(_10310_),
    .B(_10331_),
    .Y(_03325_));
 NOR2x1_ASAP7_75t_R _29435_ (.A(_00798_),
    .B(_10310_),
    .Y(_10332_));
 AO21x1_ASAP7_75t_R _29436_ (.A1(_08151_),
    .A2(_10310_),
    .B(_10332_),
    .Y(_03326_));
 TAPCELL_ASAP7_75t_R PHY_415 ();
 NOR2x1_ASAP7_75t_R _29438_ (.A(_00831_),
    .B(_10310_),
    .Y(_10334_));
 AO21x1_ASAP7_75t_R _29439_ (.A1(_08190_),
    .A2(_10310_),
    .B(_10334_),
    .Y(_03327_));
 NOR2x1_ASAP7_75t_R _29440_ (.A(_00863_),
    .B(_10310_),
    .Y(_10335_));
 AO21x1_ASAP7_75t_R _29441_ (.A1(_08225_),
    .A2(_10310_),
    .B(_10335_),
    .Y(_03328_));
 TAPCELL_ASAP7_75t_R PHY_414 ();
 NOR2x1_ASAP7_75t_R _29443_ (.A(_00896_),
    .B(_10310_),
    .Y(_10337_));
 AO21x1_ASAP7_75t_R _29444_ (.A1(_08263_),
    .A2(_10310_),
    .B(_10337_),
    .Y(_03329_));
 NOR2x1_ASAP7_75t_R _29445_ (.A(_00928_),
    .B(_10310_),
    .Y(_10338_));
 AO21x1_ASAP7_75t_R _29446_ (.A1(_08294_),
    .A2(_10310_),
    .B(_10338_),
    .Y(_03330_));
 NOR2x1_ASAP7_75t_R _29447_ (.A(_00961_),
    .B(_10310_),
    .Y(_10339_));
 AO21x1_ASAP7_75t_R _29448_ (.A1(_08328_),
    .A2(_10310_),
    .B(_10339_),
    .Y(_03331_));
 NOR2x1_ASAP7_75t_R _29449_ (.A(_00993_),
    .B(_10310_),
    .Y(_10340_));
 AO21x1_ASAP7_75t_R _29450_ (.A1(_08360_),
    .A2(_10310_),
    .B(_10340_),
    .Y(_03332_));
 NOR2x1_ASAP7_75t_R _29451_ (.A(_01027_),
    .B(_10310_),
    .Y(_10341_));
 AO21x1_ASAP7_75t_R _29452_ (.A1(_08406_),
    .A2(_10310_),
    .B(_10341_),
    .Y(_03333_));
 NOR2x1_ASAP7_75t_R _29453_ (.A(_01059_),
    .B(_10310_),
    .Y(_10342_));
 AO21x1_ASAP7_75t_R _29454_ (.A1(_08450_),
    .A2(_10310_),
    .B(_10342_),
    .Y(_03334_));
 NOR2x1_ASAP7_75t_R _29455_ (.A(_01092_),
    .B(_10310_),
    .Y(_10343_));
 AO21x1_ASAP7_75t_R _29456_ (.A1(_08481_),
    .A2(_10310_),
    .B(_10343_),
    .Y(_03335_));
 NOR2x1_ASAP7_75t_R _29457_ (.A(_01124_),
    .B(_10310_),
    .Y(_10344_));
 AO21x1_ASAP7_75t_R _29458_ (.A1(_08509_),
    .A2(_10310_),
    .B(_10344_),
    .Y(_03336_));
 NOR2x1_ASAP7_75t_R _29459_ (.A(_01158_),
    .B(_10310_),
    .Y(_10345_));
 AO21x1_ASAP7_75t_R _29460_ (.A1(_08537_),
    .A2(_10310_),
    .B(_10345_),
    .Y(_03337_));
 NOR2x1_ASAP7_75t_R _29461_ (.A(_01190_),
    .B(_10310_),
    .Y(_10346_));
 AO21x1_ASAP7_75t_R _29462_ (.A1(_08563_),
    .A2(_10310_),
    .B(_10346_),
    .Y(_03338_));
 NOR2x1_ASAP7_75t_R _29463_ (.A(_01224_),
    .B(_10310_),
    .Y(_10347_));
 AO21x1_ASAP7_75t_R _29464_ (.A1(net250),
    .A2(_10310_),
    .B(_10347_),
    .Y(_03339_));
 NOR2x1_ASAP7_75t_R _29465_ (.A(_01256_),
    .B(_10310_),
    .Y(_10348_));
 AO21x1_ASAP7_75t_R _29466_ (.A1(net2198),
    .A2(_10310_),
    .B(_10348_),
    .Y(_03340_));
 NAND2x1_ASAP7_75t_R _29467_ (.A(_08648_),
    .B(_10310_),
    .Y(_10349_));
 OA21x2_ASAP7_75t_R _29468_ (.A1(_05469_),
    .A2(_10310_),
    .B(_10349_),
    .Y(_03341_));
 OR2x6_ASAP7_75t_R _29469_ (.A(_09829_),
    .B(_10269_),
    .Y(_10350_));
 TAPCELL_ASAP7_75t_R PHY_413 ();
 NOR2x1_ASAP7_75t_R _29471_ (.A(_07248_),
    .B(_10350_),
    .Y(_10352_));
 AO21x1_ASAP7_75t_R _29472_ (.A1(_13836_),
    .A2(_10350_),
    .B(_10352_),
    .Y(_03342_));
 NOR2x2_ASAP7_75t_R _29473_ (.A(_09829_),
    .B(_10269_),
    .Y(_10353_));
 TAPCELL_ASAP7_75t_R PHY_412 ();
 AND2x2_ASAP7_75t_R _29475_ (.A(_13663_),
    .B(_10350_),
    .Y(_10355_));
 AO21x1_ASAP7_75t_R _29476_ (.A1(_07384_),
    .A2(_10353_),
    .B(_10355_),
    .Y(_03343_));
 AND2x2_ASAP7_75t_R _29477_ (.A(_14146_),
    .B(_10350_),
    .Y(_10356_));
 AO21x1_ASAP7_75t_R _29478_ (.A1(_07472_),
    .A2(_10353_),
    .B(_10356_),
    .Y(_03344_));
 AND2x2_ASAP7_75t_R _29479_ (.A(_14211_),
    .B(_10350_),
    .Y(_10357_));
 AO21x1_ASAP7_75t_R _29480_ (.A1(_07552_),
    .A2(_10353_),
    .B(_10357_),
    .Y(_03345_));
 AND2x2_ASAP7_75t_R _29481_ (.A(_14249_),
    .B(_10350_),
    .Y(_10358_));
 AO21x1_ASAP7_75t_R _29482_ (.A1(_07608_),
    .A2(_10353_),
    .B(_10358_),
    .Y(_03346_));
 AND2x2_ASAP7_75t_R _29483_ (.A(_14337_),
    .B(_10350_),
    .Y(_10359_));
 AO21x1_ASAP7_75t_R _29484_ (.A1(_07663_),
    .A2(_10353_),
    .B(_10359_),
    .Y(_03347_));
 AND2x2_ASAP7_75t_R _29485_ (.A(_14373_),
    .B(_10350_),
    .Y(_10360_));
 AO21x1_ASAP7_75t_R _29486_ (.A1(_07709_),
    .A2(_10353_),
    .B(_10360_),
    .Y(_03348_));
 TAPCELL_ASAP7_75t_R PHY_411 ();
 AND2x2_ASAP7_75t_R _29488_ (.A(_14432_),
    .B(_10350_),
    .Y(_10362_));
 AO21x1_ASAP7_75t_R _29489_ (.A1(net252),
    .A2(_10353_),
    .B(_10362_),
    .Y(_03349_));
 AND2x2_ASAP7_75t_R _29490_ (.A(_14482_),
    .B(_10350_),
    .Y(_10363_));
 AO21x1_ASAP7_75t_R _29491_ (.A1(net257),
    .A2(_10353_),
    .B(_10363_),
    .Y(_03350_));
 AND2x2_ASAP7_75t_R _29492_ (.A(_14555_),
    .B(_10350_),
    .Y(_10364_));
 AO21x1_ASAP7_75t_R _29493_ (.A1(net256),
    .A2(_10353_),
    .B(_10364_),
    .Y(_03351_));
 AND2x2_ASAP7_75t_R _29494_ (.A(_14608_),
    .B(_10350_),
    .Y(_10365_));
 AO21x1_ASAP7_75t_R _29495_ (.A1(_07903_),
    .A2(_10353_),
    .B(_10365_),
    .Y(_03352_));
 TAPCELL_ASAP7_75t_R PHY_410 ();
 AND2x2_ASAP7_75t_R _29497_ (.A(_14663_),
    .B(_10350_),
    .Y(_10367_));
 AO21x1_ASAP7_75t_R _29498_ (.A1(_07948_),
    .A2(_10353_),
    .B(_10367_),
    .Y(_03353_));
 AND2x2_ASAP7_75t_R _29499_ (.A(_14069_),
    .B(_10350_),
    .Y(_10368_));
 AO21x1_ASAP7_75t_R _29500_ (.A1(_07985_),
    .A2(_10353_),
    .B(_10368_),
    .Y(_03354_));
 AND2x2_ASAP7_75t_R _29501_ (.A(_15510_),
    .B(_10350_),
    .Y(_10369_));
 AO21x1_ASAP7_75t_R _29502_ (.A1(_08026_),
    .A2(_10353_),
    .B(_10369_),
    .Y(_03355_));
 AND2x2_ASAP7_75t_R _29503_ (.A(_15683_),
    .B(_10350_),
    .Y(_10370_));
 AO21x1_ASAP7_75t_R _29504_ (.A1(_08068_),
    .A2(_10353_),
    .B(_10370_),
    .Y(_03356_));
 AND2x2_ASAP7_75t_R _29505_ (.A(_15799_),
    .B(_10350_),
    .Y(_10371_));
 AO21x1_ASAP7_75t_R _29506_ (.A1(_08110_),
    .A2(_10353_),
    .B(_10371_),
    .Y(_03357_));
 AND2x2_ASAP7_75t_R _29507_ (.A(_15924_),
    .B(_10350_),
    .Y(_10372_));
 AO21x1_ASAP7_75t_R _29508_ (.A1(_08151_),
    .A2(_10353_),
    .B(_10372_),
    .Y(_03358_));
 TAPCELL_ASAP7_75t_R PHY_409 ();
 AND2x2_ASAP7_75t_R _29510_ (.A(_16038_),
    .B(_10350_),
    .Y(_10374_));
 AO21x1_ASAP7_75t_R _29511_ (.A1(_08190_),
    .A2(_10353_),
    .B(_10374_),
    .Y(_03359_));
 AND2x2_ASAP7_75t_R _29512_ (.A(_16169_),
    .B(_10350_),
    .Y(_10375_));
 AO21x1_ASAP7_75t_R _29513_ (.A1(_08225_),
    .A2(_10353_),
    .B(_10375_),
    .Y(_03360_));
 AND2x2_ASAP7_75t_R _29514_ (.A(_16311_),
    .B(_10350_),
    .Y(_10376_));
 AO21x1_ASAP7_75t_R _29515_ (.A1(_08263_),
    .A2(_10353_),
    .B(_10376_),
    .Y(_03361_));
 AND2x2_ASAP7_75t_R _29516_ (.A(_16415_),
    .B(_10350_),
    .Y(_10377_));
 AO21x1_ASAP7_75t_R _29517_ (.A1(_08294_),
    .A2(_10353_),
    .B(_10377_),
    .Y(_03362_));
 TAPCELL_ASAP7_75t_R PHY_408 ();
 AND2x2_ASAP7_75t_R _29519_ (.A(_16524_),
    .B(_10350_),
    .Y(_10379_));
 AO21x1_ASAP7_75t_R _29520_ (.A1(_08328_),
    .A2(_10353_),
    .B(_10379_),
    .Y(_03363_));
 AND2x2_ASAP7_75t_R _29521_ (.A(_16639_),
    .B(_10350_),
    .Y(_10380_));
 AO21x1_ASAP7_75t_R _29522_ (.A1(_08360_),
    .A2(_10353_),
    .B(_10380_),
    .Y(_03364_));
 AND2x2_ASAP7_75t_R _29523_ (.A(_04536_),
    .B(_10350_),
    .Y(_10381_));
 AO21x1_ASAP7_75t_R _29524_ (.A1(_08406_),
    .A2(_10353_),
    .B(_10381_),
    .Y(_03365_));
 AND2x2_ASAP7_75t_R _29525_ (.A(_04656_),
    .B(_10350_),
    .Y(_10382_));
 AO21x1_ASAP7_75t_R _29526_ (.A1(_08450_),
    .A2(_10353_),
    .B(_10382_),
    .Y(_03366_));
 AND2x2_ASAP7_75t_R _29527_ (.A(_04768_),
    .B(_10350_),
    .Y(_10383_));
 AO21x1_ASAP7_75t_R _29528_ (.A1(_08481_),
    .A2(_10353_),
    .B(_10383_),
    .Y(_03367_));
 AND2x2_ASAP7_75t_R _29529_ (.A(_04861_),
    .B(_10350_),
    .Y(_10384_));
 AO21x1_ASAP7_75t_R _29530_ (.A1(_08509_),
    .A2(_10353_),
    .B(_10384_),
    .Y(_03368_));
 AND2x2_ASAP7_75t_R _29531_ (.A(_04987_),
    .B(_10350_),
    .Y(_10385_));
 AO21x1_ASAP7_75t_R _29532_ (.A1(_08537_),
    .A2(_10353_),
    .B(_10385_),
    .Y(_03369_));
 AND2x2_ASAP7_75t_R _29533_ (.A(_05096_),
    .B(_10350_),
    .Y(_10386_));
 AO21x1_ASAP7_75t_R _29534_ (.A1(_08563_),
    .A2(_10353_),
    .B(_10386_),
    .Y(_03370_));
 AND2x2_ASAP7_75t_R _29535_ (.A(_05204_),
    .B(_10350_),
    .Y(_10387_));
 AO21x1_ASAP7_75t_R _29536_ (.A1(net250),
    .A2(_10353_),
    .B(_10387_),
    .Y(_03371_));
 AND2x2_ASAP7_75t_R _29537_ (.A(_05315_),
    .B(_10350_),
    .Y(_10388_));
 AO21x1_ASAP7_75t_R _29538_ (.A1(net2198),
    .A2(_10353_),
    .B(_10388_),
    .Y(_03372_));
 NOR2x1_ASAP7_75t_R _29539_ (.A(_08648_),
    .B(_10350_),
    .Y(_10389_));
 AO21x1_ASAP7_75t_R _29540_ (.A1(_05417_),
    .A2(_10350_),
    .B(_10389_),
    .Y(_03373_));
 AND4x2_ASAP7_75t_R _29541_ (.A(_00323_),
    .B(_00184_),
    .C(_14293_),
    .D(_09755_),
    .Y(_10390_));
 TAPCELL_ASAP7_75t_R PHY_407 ();
 NAND2x2_ASAP7_75t_R _29543_ (.A(_14834_),
    .B(_10390_),
    .Y(_10392_));
 TAPCELL_ASAP7_75t_R PHY_406 ();
 AND2x6_ASAP7_75t_R _29545_ (.A(_14834_),
    .B(_10390_),
    .Y(_10394_));
 AND2x2_ASAP7_75t_R _29546_ (.A(_07248_),
    .B(_10394_),
    .Y(_10395_));
 AOI21x1_ASAP7_75t_R _29547_ (.A1(_00307_),
    .A2(_10392_),
    .B(_10395_),
    .Y(_03374_));
 TAPCELL_ASAP7_75t_R PHY_405 ();
 AND2x2_ASAP7_75t_R _29549_ (.A(_13740_),
    .B(_10392_),
    .Y(_10397_));
 AO21x1_ASAP7_75t_R _29550_ (.A1(_07384_),
    .A2(_10394_),
    .B(_10397_),
    .Y(_03375_));
 TAPCELL_ASAP7_75t_R PHY_404 ();
 NOR2x1_ASAP7_75t_R _29552_ (.A(_00369_),
    .B(_10394_),
    .Y(_10399_));
 AO21x1_ASAP7_75t_R _29553_ (.A1(_07472_),
    .A2(_10394_),
    .B(_10399_),
    .Y(_03376_));
 NOR2x1_ASAP7_75t_R _29554_ (.A(_00400_),
    .B(_10394_),
    .Y(_10400_));
 AO21x1_ASAP7_75t_R _29555_ (.A1(_07552_),
    .A2(_10394_),
    .B(_10400_),
    .Y(_03377_));
 NOR2x1_ASAP7_75t_R _29556_ (.A(_00430_),
    .B(_10394_),
    .Y(_10401_));
 AO21x1_ASAP7_75t_R _29557_ (.A1(_07608_),
    .A2(_10394_),
    .B(_10401_),
    .Y(_03378_));
 NOR2x1_ASAP7_75t_R _29558_ (.A(_00460_),
    .B(_10394_),
    .Y(_10402_));
 AO21x1_ASAP7_75t_R _29559_ (.A1(_07663_),
    .A2(_10394_),
    .B(_10402_),
    .Y(_03379_));
 NOR2x1_ASAP7_75t_R _29560_ (.A(_00490_),
    .B(_10394_),
    .Y(_10403_));
 AO21x1_ASAP7_75t_R _29561_ (.A1(_07709_),
    .A2(_10394_),
    .B(_10403_),
    .Y(_03380_));
 NOR2x1_ASAP7_75t_R _29562_ (.A(_00520_),
    .B(_10394_),
    .Y(_10404_));
 AO21x1_ASAP7_75t_R _29563_ (.A1(net252),
    .A2(_10394_),
    .B(_10404_),
    .Y(_03381_));
 NOR2x1_ASAP7_75t_R _29564_ (.A(_00550_),
    .B(_10394_),
    .Y(_10405_));
 AO21x1_ASAP7_75t_R _29565_ (.A1(net257),
    .A2(_10394_),
    .B(_10405_),
    .Y(_03382_));
 NOR2x1_ASAP7_75t_R _29566_ (.A(_00580_),
    .B(_10394_),
    .Y(_10406_));
 AO21x1_ASAP7_75t_R _29567_ (.A1(net256),
    .A2(_10394_),
    .B(_10406_),
    .Y(_03383_));
 NOR2x1_ASAP7_75t_R _29568_ (.A(_00610_),
    .B(_10394_),
    .Y(_10407_));
 AO21x1_ASAP7_75t_R _29569_ (.A1(_07903_),
    .A2(_10394_),
    .B(_10407_),
    .Y(_03384_));
 TAPCELL_ASAP7_75t_R PHY_403 ();
 TAPCELL_ASAP7_75t_R PHY_402 ();
 NOR2x1_ASAP7_75t_R _29572_ (.A(_00640_),
    .B(_10394_),
    .Y(_10410_));
 AO21x1_ASAP7_75t_R _29573_ (.A1(_07948_),
    .A2(_10394_),
    .B(_10410_),
    .Y(_03385_));
 TAPCELL_ASAP7_75t_R PHY_401 ();
 NAND2x1_ASAP7_75t_R _29575_ (.A(_00339_),
    .B(_10392_),
    .Y(_10412_));
 OA21x2_ASAP7_75t_R _29576_ (.A1(_07985_),
    .A2(_10392_),
    .B(_10412_),
    .Y(_03386_));
 NOR2x1_ASAP7_75t_R _29577_ (.A(_00702_),
    .B(_10394_),
    .Y(_10413_));
 AO21x1_ASAP7_75t_R _29578_ (.A1(_08026_),
    .A2(_10394_),
    .B(_10413_),
    .Y(_03387_));
 NOR2x1_ASAP7_75t_R _29579_ (.A(_00734_),
    .B(_10394_),
    .Y(_10414_));
 AO21x1_ASAP7_75t_R _29580_ (.A1(_08068_),
    .A2(_10394_),
    .B(_10414_),
    .Y(_03388_));
 NAND2x1_ASAP7_75t_R _29581_ (.A(_00767_),
    .B(_10392_),
    .Y(_10415_));
 OA21x2_ASAP7_75t_R _29582_ (.A1(_08110_),
    .A2(_10392_),
    .B(_10415_),
    .Y(_03389_));
 NOR2x1_ASAP7_75t_R _29583_ (.A(_00800_),
    .B(_10394_),
    .Y(_10416_));
 AO21x1_ASAP7_75t_R _29584_ (.A1(_08151_),
    .A2(_10394_),
    .B(_10416_),
    .Y(_03390_));
 NOR2x1_ASAP7_75t_R _29585_ (.A(_00833_),
    .B(_10394_),
    .Y(_10417_));
 AO21x1_ASAP7_75t_R _29586_ (.A1(_08190_),
    .A2(_10394_),
    .B(_10417_),
    .Y(_03391_));
 NAND2x1_ASAP7_75t_R _29587_ (.A(_00865_),
    .B(_10392_),
    .Y(_10418_));
 OA21x2_ASAP7_75t_R _29588_ (.A1(_08225_),
    .A2(_10392_),
    .B(_10418_),
    .Y(_03392_));
 NOR2x1_ASAP7_75t_R _29589_ (.A(_00898_),
    .B(_10394_),
    .Y(_10419_));
 AO21x1_ASAP7_75t_R _29590_ (.A1(_08263_),
    .A2(_10394_),
    .B(_10419_),
    .Y(_03393_));
 AND2x2_ASAP7_75t_R _29591_ (.A(_16439_),
    .B(_10392_),
    .Y(_10420_));
 AO21x1_ASAP7_75t_R _29592_ (.A1(_08294_),
    .A2(_10394_),
    .B(_10420_),
    .Y(_03394_));
 NOR2x1_ASAP7_75t_R _29593_ (.A(_00963_),
    .B(_10394_),
    .Y(_10421_));
 AO21x1_ASAP7_75t_R _29594_ (.A1(_08328_),
    .A2(_10394_),
    .B(_10421_),
    .Y(_03395_));
 NAND2x1_ASAP7_75t_R _29595_ (.A(_00995_),
    .B(_10392_),
    .Y(_10422_));
 OA21x2_ASAP7_75t_R _29596_ (.A1(_08360_),
    .A2(_10392_),
    .B(_10422_),
    .Y(_03396_));
 NAND2x1_ASAP7_75t_R _29597_ (.A(_01029_),
    .B(_10392_),
    .Y(_10423_));
 OA21x2_ASAP7_75t_R _29598_ (.A1(_08406_),
    .A2(_10392_),
    .B(_10423_),
    .Y(_03397_));
 NAND2x1_ASAP7_75t_R _29599_ (.A(_01061_),
    .B(_10392_),
    .Y(_10424_));
 OA21x2_ASAP7_75t_R _29600_ (.A1(_08450_),
    .A2(_10392_),
    .B(_10424_),
    .Y(_03398_));
 NOR2x1_ASAP7_75t_R _29601_ (.A(_01094_),
    .B(_10394_),
    .Y(_10425_));
 AO21x1_ASAP7_75t_R _29602_ (.A1(_08481_),
    .A2(_10394_),
    .B(_10425_),
    .Y(_03399_));
 NAND2x1_ASAP7_75t_R _29603_ (.A(_01126_),
    .B(_10392_),
    .Y(_10426_));
 OA21x2_ASAP7_75t_R _29604_ (.A1(_08509_),
    .A2(_10392_),
    .B(_10426_),
    .Y(_03400_));
 NOR2x1_ASAP7_75t_R _29605_ (.A(_01160_),
    .B(_10394_),
    .Y(_10427_));
 AO21x1_ASAP7_75t_R _29606_ (.A1(_08537_),
    .A2(_10394_),
    .B(_10427_),
    .Y(_03401_));
 NOR2x1_ASAP7_75t_R _29607_ (.A(_01192_),
    .B(_10394_),
    .Y(_10428_));
 AO21x1_ASAP7_75t_R _29608_ (.A1(_08563_),
    .A2(_10394_),
    .B(_10428_),
    .Y(_03402_));
 NAND2x1_ASAP7_75t_R _29609_ (.A(_01226_),
    .B(_10392_),
    .Y(_10429_));
 OA21x2_ASAP7_75t_R _29610_ (.A1(net250),
    .A2(_10392_),
    .B(_10429_),
    .Y(_03403_));
 NAND2x1_ASAP7_75t_R _29611_ (.A(_01258_),
    .B(_10392_),
    .Y(_10430_));
 OA21x2_ASAP7_75t_R _29612_ (.A1(net2197),
    .A2(_10392_),
    .B(_10430_),
    .Y(_03404_));
 AND2x2_ASAP7_75t_R _29613_ (.A(_08648_),
    .B(_10394_),
    .Y(_10431_));
 AOI21x1_ASAP7_75t_R _29614_ (.A1(_01292_),
    .A2(_10392_),
    .B(_10431_),
    .Y(_03405_));
 OR3x4_ASAP7_75t_R _29615_ (.A(_05658_),
    .B(_00194_),
    .C(_06984_),
    .Y(_10432_));
 TAPCELL_ASAP7_75t_R PHY_400 ();
 NOR2x2_ASAP7_75t_R _29617_ (.A(_06936_),
    .B(_10432_),
    .Y(_10434_));
 TAPCELL_ASAP7_75t_R PHY_399 ();
 OR3x1_ASAP7_75t_R _29619_ (.A(_06936_),
    .B(_07248_),
    .C(_10432_),
    .Y(_10436_));
 OAI21x1_ASAP7_75t_R _29620_ (.A1(_00308_),
    .A2(_10434_),
    .B(_10436_),
    .Y(_03406_));
 TAPCELL_ASAP7_75t_R PHY_398 ();
 NOR2x1_ASAP7_75t_R _29622_ (.A(_00262_),
    .B(net270),
    .Y(_10438_));
 AO21x1_ASAP7_75t_R _29623_ (.A1(_07384_),
    .A2(net270),
    .B(_10438_),
    .Y(_03407_));
 NOR2x1_ASAP7_75t_R _29624_ (.A(_00370_),
    .B(net269),
    .Y(_10439_));
 AO21x1_ASAP7_75t_R _29625_ (.A1(_07472_),
    .A2(net269),
    .B(_10439_),
    .Y(_03408_));
 NOR2x1_ASAP7_75t_R _29626_ (.A(_00401_),
    .B(_10434_),
    .Y(_10440_));
 AO21x1_ASAP7_75t_R _29627_ (.A1(_07552_),
    .A2(_10434_),
    .B(_10440_),
    .Y(_03409_));
 NOR2x1_ASAP7_75t_R _29628_ (.A(_00431_),
    .B(net269),
    .Y(_10441_));
 AO21x1_ASAP7_75t_R _29629_ (.A1(_07608_),
    .A2(net269),
    .B(_10441_),
    .Y(_03410_));
 NOR2x1_ASAP7_75t_R _29630_ (.A(_00461_),
    .B(net269),
    .Y(_10442_));
 AO21x1_ASAP7_75t_R _29631_ (.A1(_07663_),
    .A2(net269),
    .B(_10442_),
    .Y(_03411_));
 NOR2x1_ASAP7_75t_R _29632_ (.A(_00491_),
    .B(net269),
    .Y(_10443_));
 AO21x1_ASAP7_75t_R _29633_ (.A1(_07709_),
    .A2(net269),
    .B(_10443_),
    .Y(_03412_));
 NOR2x1_ASAP7_75t_R _29634_ (.A(_00521_),
    .B(net269),
    .Y(_10444_));
 AO21x1_ASAP7_75t_R _29635_ (.A1(net252),
    .A2(net269),
    .B(_10444_),
    .Y(_03413_));
 NOR2x1_ASAP7_75t_R _29636_ (.A(_00551_),
    .B(net269),
    .Y(_10445_));
 AO21x1_ASAP7_75t_R _29637_ (.A1(net257),
    .A2(net269),
    .B(_10445_),
    .Y(_03414_));
 TAPCELL_ASAP7_75t_R PHY_397 ();
 TAPCELL_ASAP7_75t_R PHY_396 ();
 NOR2x1_ASAP7_75t_R _29640_ (.A(_00581_),
    .B(net270),
    .Y(_10448_));
 AO21x1_ASAP7_75t_R _29641_ (.A1(net256),
    .A2(net270),
    .B(_10448_),
    .Y(_03415_));
 NOR2x1_ASAP7_75t_R _29642_ (.A(_00611_),
    .B(net269),
    .Y(_10449_));
 AO21x1_ASAP7_75t_R _29643_ (.A1(_07903_),
    .A2(net269),
    .B(_10449_),
    .Y(_03416_));
 NOR2x1_ASAP7_75t_R _29644_ (.A(_00641_),
    .B(net269),
    .Y(_10450_));
 AO21x1_ASAP7_75t_R _29645_ (.A1(_07948_),
    .A2(net269),
    .B(_10450_),
    .Y(_03417_));
 NOR2x1_ASAP7_75t_R _29646_ (.A(_00340_),
    .B(net269),
    .Y(_10451_));
 AO21x1_ASAP7_75t_R _29647_ (.A1(_07985_),
    .A2(net269),
    .B(_10451_),
    .Y(_03418_));
 NOR2x1_ASAP7_75t_R _29648_ (.A(_00703_),
    .B(net270),
    .Y(_10452_));
 AO21x1_ASAP7_75t_R _29649_ (.A1(_08026_),
    .A2(net270),
    .B(_10452_),
    .Y(_03419_));
 NOR2x1_ASAP7_75t_R _29650_ (.A(_00735_),
    .B(net270),
    .Y(_10453_));
 AO21x1_ASAP7_75t_R _29651_ (.A1(_08068_),
    .A2(net270),
    .B(_10453_),
    .Y(_03420_));
 NOR2x1_ASAP7_75t_R _29652_ (.A(_00768_),
    .B(_10434_),
    .Y(_10454_));
 AO21x1_ASAP7_75t_R _29653_ (.A1(_08110_),
    .A2(_10434_),
    .B(_10454_),
    .Y(_03421_));
 NOR2x1_ASAP7_75t_R _29654_ (.A(_00801_),
    .B(net269),
    .Y(_10455_));
 AO21x1_ASAP7_75t_R _29655_ (.A1(_08151_),
    .A2(net269),
    .B(_10455_),
    .Y(_03422_));
 NOR2x1_ASAP7_75t_R _29656_ (.A(_00834_),
    .B(net270),
    .Y(_10456_));
 AO21x1_ASAP7_75t_R _29657_ (.A1(_08190_),
    .A2(net270),
    .B(_10456_),
    .Y(_03423_));
 NOR2x1_ASAP7_75t_R _29658_ (.A(_00866_),
    .B(_10434_),
    .Y(_10457_));
 AO21x1_ASAP7_75t_R _29659_ (.A1(_08225_),
    .A2(_10434_),
    .B(_10457_),
    .Y(_03424_));
 TAPCELL_ASAP7_75t_R PHY_395 ();
 TAPCELL_ASAP7_75t_R PHY_394 ();
 NOR2x1_ASAP7_75t_R _29662_ (.A(_00899_),
    .B(net270),
    .Y(_10460_));
 AO21x1_ASAP7_75t_R _29663_ (.A1(_08263_),
    .A2(net270),
    .B(_10460_),
    .Y(_03425_));
 NOR2x1_ASAP7_75t_R _29664_ (.A(_00931_),
    .B(_10434_),
    .Y(_10461_));
 AO21x1_ASAP7_75t_R _29665_ (.A1(_08294_),
    .A2(_10434_),
    .B(_10461_),
    .Y(_03426_));
 NOR2x1_ASAP7_75t_R _29666_ (.A(_00964_),
    .B(net269),
    .Y(_10462_));
 AO21x1_ASAP7_75t_R _29667_ (.A1(_08328_),
    .A2(net269),
    .B(_10462_),
    .Y(_03427_));
 NOR2x1_ASAP7_75t_R _29668_ (.A(_00996_),
    .B(_10434_),
    .Y(_10463_));
 AO21x1_ASAP7_75t_R _29669_ (.A1(_08360_),
    .A2(_10434_),
    .B(_10463_),
    .Y(_03428_));
 NOR2x1_ASAP7_75t_R _29670_ (.A(_01030_),
    .B(net270),
    .Y(_10464_));
 AO21x1_ASAP7_75t_R _29671_ (.A1(_08406_),
    .A2(net270),
    .B(_10464_),
    .Y(_03429_));
 NOR2x1_ASAP7_75t_R _29672_ (.A(_01062_),
    .B(net270),
    .Y(_10465_));
 AO21x1_ASAP7_75t_R _29673_ (.A1(_08450_),
    .A2(net270),
    .B(_10465_),
    .Y(_03430_));
 NOR2x1_ASAP7_75t_R _29674_ (.A(_01095_),
    .B(net269),
    .Y(_10466_));
 AO21x1_ASAP7_75t_R _29675_ (.A1(_08481_),
    .A2(net269),
    .B(_10466_),
    .Y(_03431_));
 NOR2x1_ASAP7_75t_R _29676_ (.A(_01127_),
    .B(net270),
    .Y(_10467_));
 AO21x1_ASAP7_75t_R _29677_ (.A1(_08509_),
    .A2(net270),
    .B(_10467_),
    .Y(_03432_));
 NOR2x1_ASAP7_75t_R _29678_ (.A(_01161_),
    .B(net270),
    .Y(_10468_));
 AO21x1_ASAP7_75t_R _29679_ (.A1(_08537_),
    .A2(net270),
    .B(_10468_),
    .Y(_03433_));
 NOR2x1_ASAP7_75t_R _29680_ (.A(_01193_),
    .B(net269),
    .Y(_10469_));
 AO21x1_ASAP7_75t_R _29681_ (.A1(_08563_),
    .A2(net269),
    .B(_10469_),
    .Y(_03434_));
 NOR2x1_ASAP7_75t_R _29682_ (.A(_01227_),
    .B(net269),
    .Y(_10470_));
 AO21x1_ASAP7_75t_R _29683_ (.A1(net250),
    .A2(net269),
    .B(_10470_),
    .Y(_03435_));
 NOR2x1_ASAP7_75t_R _29684_ (.A(_01259_),
    .B(net270),
    .Y(_10471_));
 AO21x1_ASAP7_75t_R _29685_ (.A1(net2197),
    .A2(net270),
    .B(_10471_),
    .Y(_03436_));
 OR3x1_ASAP7_75t_R _29686_ (.A(_06936_),
    .B(_08648_),
    .C(_10432_),
    .Y(_10472_));
 OAI21x1_ASAP7_75t_R _29687_ (.A1(_01293_),
    .A2(net270),
    .B(_10472_),
    .Y(_03437_));
 AND4x2_ASAP7_75t_R _29688_ (.A(_00323_),
    .B(_05658_),
    .C(_14293_),
    .D(_09755_),
    .Y(_10473_));
 AND2x6_ASAP7_75t_R _29689_ (.A(_14834_),
    .B(_10473_),
    .Y(_10474_));
 TAPCELL_ASAP7_75t_R PHY_393 ();
 TAPCELL_ASAP7_75t_R PHY_392 ();
 TAPCELL_ASAP7_75t_R PHY_391 ();
 NAND2x1_ASAP7_75t_R _29693_ (.A(_07248_),
    .B(_10474_),
    .Y(_10478_));
 OA21x2_ASAP7_75t_R _29694_ (.A1(_13874_),
    .A2(_10474_),
    .B(_10478_),
    .Y(_03438_));
 NOR2x1_ASAP7_75t_R _29695_ (.A(_00263_),
    .B(_10474_),
    .Y(_10479_));
 AO21x1_ASAP7_75t_R _29696_ (.A1(_07384_),
    .A2(_10474_),
    .B(_10479_),
    .Y(_03439_));
 NOR2x1_ASAP7_75t_R _29697_ (.A(_00371_),
    .B(_10474_),
    .Y(_10480_));
 AO21x1_ASAP7_75t_R _29698_ (.A1(_07472_),
    .A2(_10474_),
    .B(_10480_),
    .Y(_03440_));
 NOR2x1_ASAP7_75t_R _29699_ (.A(_00402_),
    .B(_10474_),
    .Y(_10481_));
 AO21x1_ASAP7_75t_R _29700_ (.A1(_07552_),
    .A2(_10474_),
    .B(_10481_),
    .Y(_03441_));
 NOR2x1_ASAP7_75t_R _29701_ (.A(_00432_),
    .B(_10474_),
    .Y(_10482_));
 AO21x1_ASAP7_75t_R _29702_ (.A1(_07608_),
    .A2(_10474_),
    .B(_10482_),
    .Y(_03442_));
 NOR2x1_ASAP7_75t_R _29703_ (.A(_00462_),
    .B(_10474_),
    .Y(_10483_));
 AO21x1_ASAP7_75t_R _29704_ (.A1(_07663_),
    .A2(_10474_),
    .B(_10483_),
    .Y(_03443_));
 NOR2x1_ASAP7_75t_R _29705_ (.A(_00492_),
    .B(_10474_),
    .Y(_10484_));
 AO21x1_ASAP7_75t_R _29706_ (.A1(_07709_),
    .A2(_10474_),
    .B(_10484_),
    .Y(_03444_));
 TAPCELL_ASAP7_75t_R PHY_390 ();
 NOR2x1_ASAP7_75t_R _29708_ (.A(_00522_),
    .B(_10474_),
    .Y(_10486_));
 AO21x1_ASAP7_75t_R _29709_ (.A1(net252),
    .A2(_10474_),
    .B(_10486_),
    .Y(_03445_));
 NOR2x1_ASAP7_75t_R _29710_ (.A(_00552_),
    .B(_10474_),
    .Y(_10487_));
 AO21x1_ASAP7_75t_R _29711_ (.A1(net257),
    .A2(_10474_),
    .B(_10487_),
    .Y(_03446_));
 TAPCELL_ASAP7_75t_R PHY_389 ();
 NOR2x1_ASAP7_75t_R _29713_ (.A(_00582_),
    .B(_10474_),
    .Y(_10489_));
 AO21x1_ASAP7_75t_R _29714_ (.A1(net256),
    .A2(_10474_),
    .B(_10489_),
    .Y(_03447_));
 NOR2x1_ASAP7_75t_R _29715_ (.A(_00612_),
    .B(_10474_),
    .Y(_10490_));
 AO21x1_ASAP7_75t_R _29716_ (.A1(_07903_),
    .A2(_10474_),
    .B(_10490_),
    .Y(_03448_));
 NOR2x1_ASAP7_75t_R _29717_ (.A(_00642_),
    .B(_10474_),
    .Y(_10491_));
 AO21x1_ASAP7_75t_R _29718_ (.A1(_07948_),
    .A2(_10474_),
    .B(_10491_),
    .Y(_03449_));
 NOR2x1_ASAP7_75t_R _29719_ (.A(_00341_),
    .B(_10474_),
    .Y(_10492_));
 AO21x1_ASAP7_75t_R _29720_ (.A1(_07985_),
    .A2(_10474_),
    .B(_10492_),
    .Y(_03450_));
 NOR2x1_ASAP7_75t_R _29721_ (.A(_00704_),
    .B(_10474_),
    .Y(_10493_));
 AO21x1_ASAP7_75t_R _29722_ (.A1(_08026_),
    .A2(_10474_),
    .B(_10493_),
    .Y(_03451_));
 NOR2x1_ASAP7_75t_R _29723_ (.A(_00736_),
    .B(_10474_),
    .Y(_10494_));
 AO21x1_ASAP7_75t_R _29724_ (.A1(_08068_),
    .A2(_10474_),
    .B(_10494_),
    .Y(_03452_));
 NOR2x1_ASAP7_75t_R _29725_ (.A(_00769_),
    .B(_10474_),
    .Y(_10495_));
 AO21x1_ASAP7_75t_R _29726_ (.A1(_08110_),
    .A2(_10474_),
    .B(_10495_),
    .Y(_03453_));
 NOR2x1_ASAP7_75t_R _29727_ (.A(_00802_),
    .B(_10474_),
    .Y(_10496_));
 AO21x1_ASAP7_75t_R _29728_ (.A1(_08151_),
    .A2(_10474_),
    .B(_10496_),
    .Y(_03454_));
 TAPCELL_ASAP7_75t_R PHY_388 ();
 NOR2x1_ASAP7_75t_R _29730_ (.A(_00835_),
    .B(_10474_),
    .Y(_10498_));
 AO21x1_ASAP7_75t_R _29731_ (.A1(_08190_),
    .A2(_10474_),
    .B(_10498_),
    .Y(_03455_));
 NOR2x1_ASAP7_75t_R _29732_ (.A(_00867_),
    .B(_10474_),
    .Y(_10499_));
 AO21x1_ASAP7_75t_R _29733_ (.A1(_08225_),
    .A2(_10474_),
    .B(_10499_),
    .Y(_03456_));
 TAPCELL_ASAP7_75t_R PHY_387 ();
 NOR2x1_ASAP7_75t_R _29735_ (.A(_00900_),
    .B(_10474_),
    .Y(_10501_));
 AO21x1_ASAP7_75t_R _29736_ (.A1(_08263_),
    .A2(_10474_),
    .B(_10501_),
    .Y(_03457_));
 NOR2x1_ASAP7_75t_R _29737_ (.A(_00932_),
    .B(_10474_),
    .Y(_10502_));
 AO21x1_ASAP7_75t_R _29738_ (.A1(_08294_),
    .A2(_10474_),
    .B(_10502_),
    .Y(_03458_));
 NOR2x1_ASAP7_75t_R _29739_ (.A(_00965_),
    .B(_10474_),
    .Y(_10503_));
 AO21x1_ASAP7_75t_R _29740_ (.A1(_08328_),
    .A2(_10474_),
    .B(_10503_),
    .Y(_03459_));
 NOR2x1_ASAP7_75t_R _29741_ (.A(_00997_),
    .B(_10474_),
    .Y(_10504_));
 AO21x1_ASAP7_75t_R _29742_ (.A1(_08360_),
    .A2(_10474_),
    .B(_10504_),
    .Y(_03460_));
 NOR2x1_ASAP7_75t_R _29743_ (.A(_01031_),
    .B(_10474_),
    .Y(_10505_));
 AO21x1_ASAP7_75t_R _29744_ (.A1(_08406_),
    .A2(_10474_),
    .B(_10505_),
    .Y(_03461_));
 NOR2x1_ASAP7_75t_R _29745_ (.A(_01063_),
    .B(_10474_),
    .Y(_10506_));
 AO21x1_ASAP7_75t_R _29746_ (.A1(_08450_),
    .A2(_10474_),
    .B(_10506_),
    .Y(_03462_));
 NOR2x1_ASAP7_75t_R _29747_ (.A(_01096_),
    .B(_10474_),
    .Y(_10507_));
 AO21x1_ASAP7_75t_R _29748_ (.A1(_08481_),
    .A2(_10474_),
    .B(_10507_),
    .Y(_03463_));
 NOR2x1_ASAP7_75t_R _29749_ (.A(_01128_),
    .B(_10474_),
    .Y(_10508_));
 AO21x1_ASAP7_75t_R _29750_ (.A1(_08509_),
    .A2(_10474_),
    .B(_10508_),
    .Y(_03464_));
 NOR2x1_ASAP7_75t_R _29751_ (.A(_01162_),
    .B(_10474_),
    .Y(_10509_));
 AO21x1_ASAP7_75t_R _29752_ (.A1(_08537_),
    .A2(_10474_),
    .B(_10509_),
    .Y(_03465_));
 NOR2x1_ASAP7_75t_R _29753_ (.A(_01194_),
    .B(_10474_),
    .Y(_10510_));
 AO21x1_ASAP7_75t_R _29754_ (.A1(_08563_),
    .A2(_10474_),
    .B(_10510_),
    .Y(_03466_));
 NOR2x1_ASAP7_75t_R _29755_ (.A(_01228_),
    .B(_10474_),
    .Y(_10511_));
 AO21x1_ASAP7_75t_R _29756_ (.A1(net250),
    .A2(_10474_),
    .B(_10511_),
    .Y(_03467_));
 NOR2x1_ASAP7_75t_R _29757_ (.A(_01260_),
    .B(_10474_),
    .Y(_10512_));
 AO21x1_ASAP7_75t_R _29758_ (.A1(net2197),
    .A2(_10474_),
    .B(_10512_),
    .Y(_03468_));
 NAND2x1_ASAP7_75t_R _29759_ (.A(_08648_),
    .B(_10474_),
    .Y(_10513_));
 OA21x2_ASAP7_75t_R _29760_ (.A1(_05408_),
    .A2(_10474_),
    .B(_10513_),
    .Y(_03469_));
 OR3x4_ASAP7_75t_R _29761_ (.A(_00184_),
    .B(_00194_),
    .C(_06984_),
    .Y(_10514_));
 TAPCELL_ASAP7_75t_R PHY_386 ();
 OR2x6_ASAP7_75t_R _29763_ (.A(_06936_),
    .B(_10514_),
    .Y(_10516_));
 TAPCELL_ASAP7_75t_R PHY_385 ();
 NOR2x1_ASAP7_75t_R _29765_ (.A(_07248_),
    .B(_10516_),
    .Y(_10518_));
 AO21x1_ASAP7_75t_R _29766_ (.A1(_13881_),
    .A2(_10516_),
    .B(_10518_),
    .Y(_03470_));
 NOR2x2_ASAP7_75t_R _29767_ (.A(_06936_),
    .B(_10514_),
    .Y(_10519_));
 TAPCELL_ASAP7_75t_R PHY_384 ();
 AND2x2_ASAP7_75t_R _29769_ (.A(_13340_),
    .B(_10516_),
    .Y(_10521_));
 AO21x1_ASAP7_75t_R _29770_ (.A1(_07384_),
    .A2(_10519_),
    .B(_10521_),
    .Y(_03471_));
 AND2x2_ASAP7_75t_R _29771_ (.A(_14870_),
    .B(_10516_),
    .Y(_10522_));
 AO21x1_ASAP7_75t_R _29772_ (.A1(_07472_),
    .A2(_10519_),
    .B(_10522_),
    .Y(_03472_));
 AND2x2_ASAP7_75t_R _29773_ (.A(_14194_),
    .B(_10516_),
    .Y(_10523_));
 AO21x1_ASAP7_75t_R _29774_ (.A1(_07552_),
    .A2(_10519_),
    .B(_10523_),
    .Y(_03473_));
 AND2x2_ASAP7_75t_R _29775_ (.A(_15002_),
    .B(_10516_),
    .Y(_10524_));
 AO21x1_ASAP7_75t_R _29776_ (.A1(_07608_),
    .A2(_10519_),
    .B(_10524_),
    .Y(_03474_));
 AND2x2_ASAP7_75t_R _29777_ (.A(_14301_),
    .B(_10516_),
    .Y(_10525_));
 AO21x1_ASAP7_75t_R _29778_ (.A1(_07663_),
    .A2(_10519_),
    .B(_10525_),
    .Y(_03475_));
 AND2x2_ASAP7_75t_R _29779_ (.A(_15125_),
    .B(_10516_),
    .Y(_10526_));
 AO21x1_ASAP7_75t_R _29780_ (.A1(_07709_),
    .A2(_10519_),
    .B(_10526_),
    .Y(_03476_));
 TAPCELL_ASAP7_75t_R PHY_383 ();
 AND2x2_ASAP7_75t_R _29782_ (.A(_15215_),
    .B(_10516_),
    .Y(_10528_));
 AO21x1_ASAP7_75t_R _29783_ (.A1(net252),
    .A2(_10519_),
    .B(_10528_),
    .Y(_03477_));
 AND2x2_ASAP7_75t_R _29784_ (.A(_14534_),
    .B(_10516_),
    .Y(_10529_));
 AO21x1_ASAP7_75t_R _29785_ (.A1(net257),
    .A2(_10519_),
    .B(_10529_),
    .Y(_03478_));
 AND2x2_ASAP7_75t_R _29786_ (.A(_14582_),
    .B(_10516_),
    .Y(_10530_));
 AO21x1_ASAP7_75t_R _29787_ (.A1(net256),
    .A2(_10519_),
    .B(_10530_),
    .Y(_03479_));
 AND2x2_ASAP7_75t_R _29788_ (.A(_15351_),
    .B(_10516_),
    .Y(_10531_));
 AO21x1_ASAP7_75t_R _29789_ (.A1(_07903_),
    .A2(_10519_),
    .B(_10531_),
    .Y(_03480_));
 TAPCELL_ASAP7_75t_R PHY_382 ();
 AND2x2_ASAP7_75t_R _29791_ (.A(_14729_),
    .B(_10516_),
    .Y(_10533_));
 AO21x1_ASAP7_75t_R _29792_ (.A1(_07948_),
    .A2(_10519_),
    .B(_10533_),
    .Y(_03481_));
 AND2x2_ASAP7_75t_R _29793_ (.A(_14043_),
    .B(_10516_),
    .Y(_10534_));
 AO21x1_ASAP7_75t_R _29794_ (.A1(_07985_),
    .A2(_10519_),
    .B(_10534_),
    .Y(_03482_));
 AND2x2_ASAP7_75t_R _29795_ (.A(_15551_),
    .B(_10516_),
    .Y(_10535_));
 AO21x1_ASAP7_75t_R _29796_ (.A1(_08026_),
    .A2(_10519_),
    .B(_10535_),
    .Y(_03483_));
 AND2x2_ASAP7_75t_R _29797_ (.A(_15699_),
    .B(_10516_),
    .Y(_10536_));
 AO21x1_ASAP7_75t_R _29798_ (.A1(_08068_),
    .A2(_10519_),
    .B(_10536_),
    .Y(_03484_));
 AND2x2_ASAP7_75t_R _29799_ (.A(_15808_),
    .B(_10516_),
    .Y(_10537_));
 AO21x1_ASAP7_75t_R _29800_ (.A1(_08110_),
    .A2(_10519_),
    .B(_10537_),
    .Y(_03485_));
 AND2x2_ASAP7_75t_R _29801_ (.A(_15955_),
    .B(_10516_),
    .Y(_10538_));
 AO21x1_ASAP7_75t_R _29802_ (.A1(_08151_),
    .A2(_10519_),
    .B(_10538_),
    .Y(_03486_));
 TAPCELL_ASAP7_75t_R PHY_381 ();
 AND2x2_ASAP7_75t_R _29804_ (.A(_16061_),
    .B(_10516_),
    .Y(_10540_));
 AO21x1_ASAP7_75t_R _29805_ (.A1(_08190_),
    .A2(_10519_),
    .B(_10540_),
    .Y(_03487_));
 AND2x2_ASAP7_75t_R _29806_ (.A(_16204_),
    .B(_10516_),
    .Y(_10541_));
 AO21x1_ASAP7_75t_R _29807_ (.A1(_08225_),
    .A2(_10519_),
    .B(_10541_),
    .Y(_03488_));
 AND2x2_ASAP7_75t_R _29808_ (.A(_16272_),
    .B(_10516_),
    .Y(_10542_));
 AO21x1_ASAP7_75t_R _29809_ (.A1(_08263_),
    .A2(_10519_),
    .B(_10542_),
    .Y(_03489_));
 AND2x2_ASAP7_75t_R _29810_ (.A(_16442_),
    .B(_10516_),
    .Y(_10543_));
 AO21x1_ASAP7_75t_R _29811_ (.A1(_08294_),
    .A2(_10519_),
    .B(_10543_),
    .Y(_03490_));
 TAPCELL_ASAP7_75t_R PHY_380 ();
 AND2x2_ASAP7_75t_R _29813_ (.A(_16544_),
    .B(_10516_),
    .Y(_10545_));
 AO21x1_ASAP7_75t_R _29814_ (.A1(_08328_),
    .A2(_10519_),
    .B(_10545_),
    .Y(_03491_));
 AND2x2_ASAP7_75t_R _29815_ (.A(_16655_),
    .B(_10516_),
    .Y(_10546_));
 AO21x1_ASAP7_75t_R _29816_ (.A1(_08360_),
    .A2(_10519_),
    .B(_10546_),
    .Y(_03492_));
 AND2x2_ASAP7_75t_R _29817_ (.A(_04567_),
    .B(_10516_),
    .Y(_10547_));
 AO21x1_ASAP7_75t_R _29818_ (.A1(_08406_),
    .A2(_10519_),
    .B(_10547_),
    .Y(_03493_));
 AND2x2_ASAP7_75t_R _29819_ (.A(_04673_),
    .B(_10516_),
    .Y(_10548_));
 AO21x1_ASAP7_75t_R _29820_ (.A1(_08450_),
    .A2(_10519_),
    .B(_10548_),
    .Y(_03494_));
 AND2x2_ASAP7_75t_R _29821_ (.A(_04784_),
    .B(_10516_),
    .Y(_10549_));
 AO21x1_ASAP7_75t_R _29822_ (.A1(_08481_),
    .A2(_10519_),
    .B(_10549_),
    .Y(_03495_));
 AND2x2_ASAP7_75t_R _29823_ (.A(_04885_),
    .B(_10516_),
    .Y(_10550_));
 AO21x1_ASAP7_75t_R _29824_ (.A1(_08509_),
    .A2(_10519_),
    .B(_10550_),
    .Y(_03496_));
 AND2x2_ASAP7_75t_R _29825_ (.A(_05019_),
    .B(_10516_),
    .Y(_10551_));
 AO21x1_ASAP7_75t_R _29826_ (.A1(_08537_),
    .A2(_10519_),
    .B(_10551_),
    .Y(_03497_));
 AND2x2_ASAP7_75t_R _29827_ (.A(_05120_),
    .B(_10516_),
    .Y(_10552_));
 AO21x1_ASAP7_75t_R _29828_ (.A1(_08563_),
    .A2(_10519_),
    .B(_10552_),
    .Y(_03498_));
 AND2x2_ASAP7_75t_R _29829_ (.A(_05228_),
    .B(_10516_),
    .Y(_10553_));
 AO21x1_ASAP7_75t_R _29830_ (.A1(net250),
    .A2(_10519_),
    .B(_10553_),
    .Y(_03499_));
 AND2x2_ASAP7_75t_R _29831_ (.A(_05331_),
    .B(_10516_),
    .Y(_10554_));
 AO21x1_ASAP7_75t_R _29832_ (.A1(net2197),
    .A2(_10519_),
    .B(_10554_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _29833_ (.A(_08648_),
    .B(_10516_),
    .Y(_10555_));
 AO21x1_ASAP7_75t_R _29834_ (.A1(_05405_),
    .A2(_10516_),
    .B(_10555_),
    .Y(_03501_));
 NAND2x2_ASAP7_75t_R _29835_ (.A(_09872_),
    .B(_10390_),
    .Y(_10556_));
 AND2x6_ASAP7_75t_R _29836_ (.A(_09872_),
    .B(_10390_),
    .Y(_10557_));
 TAPCELL_ASAP7_75t_R PHY_379 ();
 AND2x2_ASAP7_75t_R _29838_ (.A(_07248_),
    .B(_10557_),
    .Y(_10559_));
 AOI21x1_ASAP7_75t_R _29839_ (.A1(_00311_),
    .A2(_10556_),
    .B(_10559_),
    .Y(_03502_));
 TAPCELL_ASAP7_75t_R PHY_378 ();
 TAPCELL_ASAP7_75t_R PHY_377 ();
 NOR2x1_ASAP7_75t_R _29842_ (.A(_00265_),
    .B(_10557_),
    .Y(_10562_));
 AO21x1_ASAP7_75t_R _29843_ (.A1(_07384_),
    .A2(_10557_),
    .B(_10562_),
    .Y(_03503_));
 AND2x2_ASAP7_75t_R _29844_ (.A(_14114_),
    .B(_10556_),
    .Y(_10563_));
 AO21x1_ASAP7_75t_R _29845_ (.A1(_07472_),
    .A2(_10557_),
    .B(_10563_),
    .Y(_03504_));
 NOR2x1_ASAP7_75t_R _29846_ (.A(_00404_),
    .B(_10557_),
    .Y(_10564_));
 AO21x1_ASAP7_75t_R _29847_ (.A1(_07552_),
    .A2(_10557_),
    .B(_10564_),
    .Y(_03505_));
 NOR2x1_ASAP7_75t_R _29848_ (.A(_00434_),
    .B(_10557_),
    .Y(_10565_));
 AO21x1_ASAP7_75t_R _29849_ (.A1(_07608_),
    .A2(_10557_),
    .B(_10565_),
    .Y(_03506_));
 NOR2x1_ASAP7_75t_R _29850_ (.A(_00464_),
    .B(_10557_),
    .Y(_10566_));
 AO21x1_ASAP7_75t_R _29851_ (.A1(_07663_),
    .A2(_10557_),
    .B(_10566_),
    .Y(_03507_));
 NOR2x1_ASAP7_75t_R _29852_ (.A(_00494_),
    .B(_10557_),
    .Y(_10567_));
 AO21x1_ASAP7_75t_R _29853_ (.A1(_07709_),
    .A2(_10557_),
    .B(_10567_),
    .Y(_03508_));
 NOR2x1_ASAP7_75t_R _29854_ (.A(_00524_),
    .B(_10557_),
    .Y(_10568_));
 AO21x1_ASAP7_75t_R _29855_ (.A1(net252),
    .A2(_10557_),
    .B(_10568_),
    .Y(_03509_));
 NOR2x1_ASAP7_75t_R _29856_ (.A(_00554_),
    .B(_10557_),
    .Y(_10569_));
 AO21x1_ASAP7_75t_R _29857_ (.A1(net257),
    .A2(_10557_),
    .B(_10569_),
    .Y(_03510_));
 NOR2x1_ASAP7_75t_R _29858_ (.A(_00584_),
    .B(_10557_),
    .Y(_10570_));
 AO21x1_ASAP7_75t_R _29859_ (.A1(net256),
    .A2(_10557_),
    .B(_10570_),
    .Y(_03511_));
 NOR2x1_ASAP7_75t_R _29860_ (.A(_00614_),
    .B(_10557_),
    .Y(_10571_));
 AO21x1_ASAP7_75t_R _29861_ (.A1(_07903_),
    .A2(_10557_),
    .B(_10571_),
    .Y(_03512_));
 TAPCELL_ASAP7_75t_R PHY_376 ();
 AND2x2_ASAP7_75t_R _29863_ (.A(_14695_),
    .B(_10556_),
    .Y(_10573_));
 AO21x1_ASAP7_75t_R _29864_ (.A1(_07948_),
    .A2(_10557_),
    .B(_10573_),
    .Y(_03513_));
 NOR2x1_ASAP7_75t_R _29865_ (.A(_00343_),
    .B(_10557_),
    .Y(_10574_));
 AO21x1_ASAP7_75t_R _29866_ (.A1(_07985_),
    .A2(_10557_),
    .B(_10574_),
    .Y(_03514_));
 TAPCELL_ASAP7_75t_R PHY_375 ();
 NOR2x1_ASAP7_75t_R _29868_ (.A(_00706_),
    .B(_10557_),
    .Y(_10576_));
 AO21x1_ASAP7_75t_R _29869_ (.A1(_08026_),
    .A2(_10557_),
    .B(_10576_),
    .Y(_03515_));
 NOR2x1_ASAP7_75t_R _29870_ (.A(_00738_),
    .B(_10557_),
    .Y(_10577_));
 AO21x1_ASAP7_75t_R _29871_ (.A1(_08068_),
    .A2(_10557_),
    .B(_10577_),
    .Y(_03516_));
 NOR2x1_ASAP7_75t_R _29872_ (.A(_00771_),
    .B(_10557_),
    .Y(_10578_));
 AO21x1_ASAP7_75t_R _29873_ (.A1(_08110_),
    .A2(_10557_),
    .B(_10578_),
    .Y(_03517_));
 NOR2x1_ASAP7_75t_R _29874_ (.A(_00804_),
    .B(_10557_),
    .Y(_10579_));
 AO21x1_ASAP7_75t_R _29875_ (.A1(_08151_),
    .A2(_10557_),
    .B(_10579_),
    .Y(_03518_));
 NOR2x1_ASAP7_75t_R _29876_ (.A(_00837_),
    .B(_10557_),
    .Y(_10580_));
 AO21x1_ASAP7_75t_R _29877_ (.A1(_08190_),
    .A2(_10557_),
    .B(_10580_),
    .Y(_03519_));
 NOR2x1_ASAP7_75t_R _29878_ (.A(_00869_),
    .B(_10557_),
    .Y(_10581_));
 AO21x1_ASAP7_75t_R _29879_ (.A1(_08225_),
    .A2(_10557_),
    .B(_10581_),
    .Y(_03520_));
 NOR2x1_ASAP7_75t_R _29880_ (.A(_00902_),
    .B(_10557_),
    .Y(_10582_));
 AO21x1_ASAP7_75t_R _29881_ (.A1(_08263_),
    .A2(_10557_),
    .B(_10582_),
    .Y(_03521_));
 AND2x2_ASAP7_75t_R _29882_ (.A(_16488_),
    .B(_10556_),
    .Y(_10583_));
 AO21x1_ASAP7_75t_R _29883_ (.A1(_08294_),
    .A2(_10557_),
    .B(_10583_),
    .Y(_03522_));
 TAPCELL_ASAP7_75t_R PHY_374 ();
 NOR2x1_ASAP7_75t_R _29885_ (.A(_00967_),
    .B(_10557_),
    .Y(_10585_));
 AO21x1_ASAP7_75t_R _29886_ (.A1(_08328_),
    .A2(_10557_),
    .B(_10585_),
    .Y(_03523_));
 NOR2x1_ASAP7_75t_R _29887_ (.A(_00999_),
    .B(_10557_),
    .Y(_10586_));
 AO21x1_ASAP7_75t_R _29888_ (.A1(_08360_),
    .A2(_10557_),
    .B(_10586_),
    .Y(_03524_));
 NOR2x1_ASAP7_75t_R _29889_ (.A(_01033_),
    .B(_10557_),
    .Y(_10587_));
 AO21x1_ASAP7_75t_R _29890_ (.A1(_08406_),
    .A2(_10557_),
    .B(_10587_),
    .Y(_03525_));
 NOR2x1_ASAP7_75t_R _29891_ (.A(_01065_),
    .B(_10557_),
    .Y(_10588_));
 AO21x1_ASAP7_75t_R _29892_ (.A1(_08450_),
    .A2(_10557_),
    .B(_10588_),
    .Y(_03526_));
 NOR2x1_ASAP7_75t_R _29893_ (.A(_01098_),
    .B(_10557_),
    .Y(_10589_));
 AO21x1_ASAP7_75t_R _29894_ (.A1(_08481_),
    .A2(_10557_),
    .B(_10589_),
    .Y(_03527_));
 NOR2x1_ASAP7_75t_R _29895_ (.A(_01130_),
    .B(_10557_),
    .Y(_10590_));
 AO21x1_ASAP7_75t_R _29896_ (.A1(_08509_),
    .A2(_10557_),
    .B(_10590_),
    .Y(_03528_));
 NOR2x1_ASAP7_75t_R _29897_ (.A(_01164_),
    .B(_10557_),
    .Y(_10591_));
 AO21x1_ASAP7_75t_R _29898_ (.A1(_08537_),
    .A2(_10557_),
    .B(_10591_),
    .Y(_03529_));
 NOR2x1_ASAP7_75t_R _29899_ (.A(_01196_),
    .B(_10557_),
    .Y(_10592_));
 AO21x1_ASAP7_75t_R _29900_ (.A1(_08563_),
    .A2(_10557_),
    .B(_10592_),
    .Y(_03530_));
 NOR2x1_ASAP7_75t_R _29901_ (.A(_01230_),
    .B(_10557_),
    .Y(_10593_));
 AO21x1_ASAP7_75t_R _29902_ (.A1(net250),
    .A2(_10557_),
    .B(_10593_),
    .Y(_03531_));
 NOR2x1_ASAP7_75t_R _29903_ (.A(_01262_),
    .B(_10557_),
    .Y(_10594_));
 AO21x1_ASAP7_75t_R _29904_ (.A1(net2197),
    .A2(_10557_),
    .B(_10594_),
    .Y(_03532_));
 AND2x2_ASAP7_75t_R _29905_ (.A(_08648_),
    .B(_10557_),
    .Y(_10595_));
 AOI21x1_ASAP7_75t_R _29906_ (.A1(_01296_),
    .A2(_10556_),
    .B(_10595_),
    .Y(_03533_));
 NOR2x2_ASAP7_75t_R _29907_ (.A(_09914_),
    .B(_10432_),
    .Y(_10596_));
 TAPCELL_ASAP7_75t_R PHY_373 ();
 OR3x1_ASAP7_75t_R _29909_ (.A(_07248_),
    .B(_09914_),
    .C(_10432_),
    .Y(_10598_));
 OAI21x1_ASAP7_75t_R _29910_ (.A1(_00312_),
    .A2(_10596_),
    .B(_10598_),
    .Y(_03534_));
 TAPCELL_ASAP7_75t_R PHY_372 ();
 TAPCELL_ASAP7_75t_R PHY_371 ();
 NOR2x1_ASAP7_75t_R _29913_ (.A(_00266_),
    .B(net268),
    .Y(_10601_));
 AO21x1_ASAP7_75t_R _29914_ (.A1(_07384_),
    .A2(net268),
    .B(_10601_),
    .Y(_03535_));
 NOR2x1_ASAP7_75t_R _29915_ (.A(_00374_),
    .B(net268),
    .Y(_10602_));
 AO21x1_ASAP7_75t_R _29916_ (.A1(_07472_),
    .A2(net268),
    .B(_10602_),
    .Y(_03536_));
 NOR2x1_ASAP7_75t_R _29917_ (.A(_00405_),
    .B(_10596_),
    .Y(_10603_));
 AO21x1_ASAP7_75t_R _29918_ (.A1(_07552_),
    .A2(_10596_),
    .B(_10603_),
    .Y(_03537_));
 NOR2x1_ASAP7_75t_R _29919_ (.A(_00435_),
    .B(net268),
    .Y(_10604_));
 AO21x1_ASAP7_75t_R _29920_ (.A1(_07608_),
    .A2(net268),
    .B(_10604_),
    .Y(_03538_));
 TAPCELL_ASAP7_75t_R PHY_370 ();
 NOR2x1_ASAP7_75t_R _29922_ (.A(_00465_),
    .B(net267),
    .Y(_10606_));
 AO21x1_ASAP7_75t_R _29923_ (.A1(_07663_),
    .A2(net267),
    .B(_10606_),
    .Y(_03539_));
 NOR2x1_ASAP7_75t_R _29924_ (.A(_00495_),
    .B(net268),
    .Y(_10607_));
 AO21x1_ASAP7_75t_R _29925_ (.A1(_07709_),
    .A2(net268),
    .B(_10607_),
    .Y(_03540_));
 NOR2x1_ASAP7_75t_R _29926_ (.A(_00525_),
    .B(net268),
    .Y(_10608_));
 AO21x1_ASAP7_75t_R _29927_ (.A1(net252),
    .A2(net268),
    .B(_10608_),
    .Y(_03541_));
 TAPCELL_ASAP7_75t_R PHY_369 ();
 NOR2x1_ASAP7_75t_R _29929_ (.A(_00555_),
    .B(net268),
    .Y(_10610_));
 AO21x1_ASAP7_75t_R _29930_ (.A1(net257),
    .A2(net268),
    .B(_10610_),
    .Y(_03542_));
 TAPCELL_ASAP7_75t_R PHY_368 ();
 TAPCELL_ASAP7_75t_R PHY_367 ();
 NOR2x1_ASAP7_75t_R _29933_ (.A(_00585_),
    .B(_10596_),
    .Y(_10613_));
 AO21x1_ASAP7_75t_R _29934_ (.A1(net256),
    .A2(_10596_),
    .B(_10613_),
    .Y(_03543_));
 NOR2x1_ASAP7_75t_R _29935_ (.A(_00615_),
    .B(net267),
    .Y(_10614_));
 AO21x1_ASAP7_75t_R _29936_ (.A1(_07903_),
    .A2(net267),
    .B(_10614_),
    .Y(_03544_));
 NOR2x1_ASAP7_75t_R _29937_ (.A(_00645_),
    .B(net268),
    .Y(_10615_));
 AO21x1_ASAP7_75t_R _29938_ (.A1(_07948_),
    .A2(net268),
    .B(_10615_),
    .Y(_03545_));
 NOR2x1_ASAP7_75t_R _29939_ (.A(_00344_),
    .B(net267),
    .Y(_10616_));
 AO21x1_ASAP7_75t_R _29940_ (.A1(_07985_),
    .A2(net267),
    .B(_10616_),
    .Y(_03546_));
 TAPCELL_ASAP7_75t_R PHY_366 ();
 NOR2x1_ASAP7_75t_R _29942_ (.A(_00707_),
    .B(_10596_),
    .Y(_10618_));
 AO21x1_ASAP7_75t_R _29943_ (.A1(_08026_),
    .A2(_10596_),
    .B(_10618_),
    .Y(_03547_));
 NOR2x1_ASAP7_75t_R _29944_ (.A(_00739_),
    .B(net267),
    .Y(_10619_));
 AO21x1_ASAP7_75t_R _29945_ (.A1(_08068_),
    .A2(net267),
    .B(_10619_),
    .Y(_03548_));
 TAPCELL_ASAP7_75t_R PHY_365 ();
 NOR2x1_ASAP7_75t_R _29947_ (.A(_00772_),
    .B(_10596_),
    .Y(_10621_));
 AO21x1_ASAP7_75t_R _29948_ (.A1(_08110_),
    .A2(_10596_),
    .B(_10621_),
    .Y(_03549_));
 TAPCELL_ASAP7_75t_R PHY_364 ();
 NOR2x1_ASAP7_75t_R _29950_ (.A(_00805_),
    .B(net268),
    .Y(_10623_));
 AO21x1_ASAP7_75t_R _29951_ (.A1(_08151_),
    .A2(net268),
    .B(_10623_),
    .Y(_03550_));
 NOR2x1_ASAP7_75t_R _29952_ (.A(_00838_),
    .B(net267),
    .Y(_10624_));
 AO21x1_ASAP7_75t_R _29953_ (.A1(_08190_),
    .A2(net267),
    .B(_10624_),
    .Y(_03551_));
 NOR2x1_ASAP7_75t_R _29954_ (.A(_00870_),
    .B(_10596_),
    .Y(_10625_));
 AO21x1_ASAP7_75t_R _29955_ (.A1(_08225_),
    .A2(_10596_),
    .B(_10625_),
    .Y(_03552_));
 TAPCELL_ASAP7_75t_R PHY_363 ();
 TAPCELL_ASAP7_75t_R PHY_362 ();
 NOR2x1_ASAP7_75t_R _29958_ (.A(_00903_),
    .B(net267),
    .Y(_10628_));
 AO21x1_ASAP7_75t_R _29959_ (.A1(_08263_),
    .A2(net267),
    .B(_10628_),
    .Y(_03553_));
 TAPCELL_ASAP7_75t_R PHY_361 ();
 NOR2x1_ASAP7_75t_R _29961_ (.A(_00935_),
    .B(_10596_),
    .Y(_10630_));
 AO21x1_ASAP7_75t_R _29962_ (.A1(_08294_),
    .A2(_10596_),
    .B(_10630_),
    .Y(_03554_));
 NOR2x1_ASAP7_75t_R _29963_ (.A(_00968_),
    .B(net267),
    .Y(_10631_));
 AO21x1_ASAP7_75t_R _29964_ (.A1(_08328_),
    .A2(net267),
    .B(_10631_),
    .Y(_03555_));
 TAPCELL_ASAP7_75t_R PHY_360 ();
 NOR2x1_ASAP7_75t_R _29966_ (.A(_01000_),
    .B(_10596_),
    .Y(_10633_));
 AO21x1_ASAP7_75t_R _29967_ (.A1(_08360_),
    .A2(_10596_),
    .B(_10633_),
    .Y(_03556_));
 NOR2x1_ASAP7_75t_R _29968_ (.A(_01034_),
    .B(net267),
    .Y(_10634_));
 AO21x1_ASAP7_75t_R _29969_ (.A1(_08406_),
    .A2(net267),
    .B(_10634_),
    .Y(_03557_));
 TAPCELL_ASAP7_75t_R PHY_359 ();
 NOR2x1_ASAP7_75t_R _29971_ (.A(_01066_),
    .B(_10596_),
    .Y(_10636_));
 AO21x1_ASAP7_75t_R _29972_ (.A1(_08450_),
    .A2(_10596_),
    .B(_10636_),
    .Y(_03558_));
 NOR2x1_ASAP7_75t_R _29973_ (.A(_01099_),
    .B(net268),
    .Y(_10637_));
 AO21x1_ASAP7_75t_R _29974_ (.A1(_08481_),
    .A2(net268),
    .B(_10637_),
    .Y(_03559_));
 TAPCELL_ASAP7_75t_R PHY_358 ();
 NOR2x1_ASAP7_75t_R _29976_ (.A(_01131_),
    .B(net267),
    .Y(_10639_));
 AO21x1_ASAP7_75t_R _29977_ (.A1(_08509_),
    .A2(net267),
    .B(_10639_),
    .Y(_03560_));
 NOR2x1_ASAP7_75t_R _29978_ (.A(_01165_),
    .B(net267),
    .Y(_10640_));
 AO21x1_ASAP7_75t_R _29979_ (.A1(_08537_),
    .A2(net267),
    .B(_10640_),
    .Y(_03561_));
 TAPCELL_ASAP7_75t_R PHY_357 ();
 NOR2x1_ASAP7_75t_R _29981_ (.A(_01197_),
    .B(net267),
    .Y(_10642_));
 AO21x1_ASAP7_75t_R _29982_ (.A1(_08563_),
    .A2(net267),
    .B(_10642_),
    .Y(_03562_));
 NOR2x1_ASAP7_75t_R _29983_ (.A(_01231_),
    .B(net267),
    .Y(_10643_));
 AO21x1_ASAP7_75t_R _29984_ (.A1(net250),
    .A2(net267),
    .B(_10643_),
    .Y(_03563_));
 TAPCELL_ASAP7_75t_R PHY_356 ();
 NOR2x1_ASAP7_75t_R _29986_ (.A(_01263_),
    .B(_10596_),
    .Y(_10645_));
 AO21x1_ASAP7_75t_R _29987_ (.A1(net2197),
    .A2(_10596_),
    .B(_10645_),
    .Y(_03564_));
 OR3x1_ASAP7_75t_R _29988_ (.A(_08648_),
    .B(_09914_),
    .C(_10432_),
    .Y(_10646_));
 OAI21x1_ASAP7_75t_R _29989_ (.A1(_01297_),
    .A2(_10596_),
    .B(_10646_),
    .Y(_03565_));
 NAND2x2_ASAP7_75t_R _29990_ (.A(_09872_),
    .B(_10473_),
    .Y(_10647_));
 TAPCELL_ASAP7_75t_R PHY_355 ();
 NOR2x1_ASAP7_75t_R _29992_ (.A(_07248_),
    .B(_10647_),
    .Y(_10649_));
 AO21x1_ASAP7_75t_R _29993_ (.A1(_13871_),
    .A2(_10647_),
    .B(_10649_),
    .Y(_03566_));
 AND2x6_ASAP7_75t_R _29994_ (.A(_09872_),
    .B(_10473_),
    .Y(_10650_));
 TAPCELL_ASAP7_75t_R PHY_354 ();
 AND2x2_ASAP7_75t_R _29996_ (.A(_13718_),
    .B(_10647_),
    .Y(_10652_));
 AO21x1_ASAP7_75t_R _29997_ (.A1(_07384_),
    .A2(_10650_),
    .B(_10652_),
    .Y(_03567_));
 TAPCELL_ASAP7_75t_R PHY_353 ();
 AND2x2_ASAP7_75t_R _29999_ (.A(_14864_),
    .B(_10647_),
    .Y(_10654_));
 AO21x1_ASAP7_75t_R _30000_ (.A1(_07472_),
    .A2(_10650_),
    .B(_10654_),
    .Y(_03568_));
 TAPCELL_ASAP7_75t_R PHY_352 ();
 AND2x2_ASAP7_75t_R _30002_ (.A(_14970_),
    .B(_10647_),
    .Y(_10656_));
 AO21x1_ASAP7_75t_R _30003_ (.A1(_07552_),
    .A2(_10650_),
    .B(_10656_),
    .Y(_03569_));
 TAPCELL_ASAP7_75t_R PHY_351 ();
 AND2x2_ASAP7_75t_R _30005_ (.A(_14264_),
    .B(_10647_),
    .Y(_10658_));
 AO21x1_ASAP7_75t_R _30006_ (.A1(_07608_),
    .A2(_10650_),
    .B(_10658_),
    .Y(_03570_));
 AND2x2_ASAP7_75t_R _30007_ (.A(_14309_),
    .B(_10647_),
    .Y(_10659_));
 AO21x1_ASAP7_75t_R _30008_ (.A1(_07663_),
    .A2(_10650_),
    .B(_10659_),
    .Y(_03571_));
 TAPCELL_ASAP7_75t_R PHY_350 ();
 AND2x2_ASAP7_75t_R _30010_ (.A(_14395_),
    .B(_10647_),
    .Y(_10661_));
 AO21x1_ASAP7_75t_R _30011_ (.A1(_07709_),
    .A2(_10650_),
    .B(_10661_),
    .Y(_03572_));
 TAPCELL_ASAP7_75t_R PHY_349 ();
 TAPCELL_ASAP7_75t_R PHY_348 ();
 AND2x2_ASAP7_75t_R _30014_ (.A(_14456_),
    .B(_10647_),
    .Y(_10664_));
 AO21x1_ASAP7_75t_R _30015_ (.A1(net252),
    .A2(_10650_),
    .B(_10664_),
    .Y(_03573_));
 AND2x2_ASAP7_75t_R _30016_ (.A(_14524_),
    .B(_10647_),
    .Y(_10665_));
 AO21x1_ASAP7_75t_R _30017_ (.A1(net257),
    .A2(_10650_),
    .B(_10665_),
    .Y(_03574_));
 TAPCELL_ASAP7_75t_R PHY_347 ();
 AND2x2_ASAP7_75t_R _30019_ (.A(_14579_),
    .B(_10647_),
    .Y(_10667_));
 AO21x1_ASAP7_75t_R _30020_ (.A1(net256),
    .A2(_10650_),
    .B(_10667_),
    .Y(_03575_));
 TAPCELL_ASAP7_75t_R PHY_346 ();
 AND2x2_ASAP7_75t_R _30022_ (.A(_14629_),
    .B(_10647_),
    .Y(_10669_));
 AO21x1_ASAP7_75t_R _30023_ (.A1(_07903_),
    .A2(_10650_),
    .B(_10669_),
    .Y(_03576_));
 TAPCELL_ASAP7_75t_R PHY_345 ();
 TAPCELL_ASAP7_75t_R PHY_344 ();
 AND2x2_ASAP7_75t_R _30026_ (.A(_14716_),
    .B(_10647_),
    .Y(_10672_));
 AO21x1_ASAP7_75t_R _30027_ (.A1(_07948_),
    .A2(_10650_),
    .B(_10672_),
    .Y(_03577_));
 AND3x1_ASAP7_75t_R _30028_ (.A(_07961_),
    .B(_07984_),
    .C(_10650_),
    .Y(_10673_));
 AO21x1_ASAP7_75t_R _30029_ (.A1(_14027_),
    .A2(_10647_),
    .B(_10673_),
    .Y(_03578_));
 AND2x2_ASAP7_75t_R _30030_ (.A(_15567_),
    .B(_10647_),
    .Y(_10674_));
 AO21x1_ASAP7_75t_R _30031_ (.A1(_08026_),
    .A2(_10650_),
    .B(_10674_),
    .Y(_03579_));
 TAPCELL_ASAP7_75t_R PHY_343 ();
 AND2x2_ASAP7_75t_R _30033_ (.A(_15695_),
    .B(_10647_),
    .Y(_10676_));
 AO21x1_ASAP7_75t_R _30034_ (.A1(_08068_),
    .A2(_10650_),
    .B(_10676_),
    .Y(_03580_));
 AND2x2_ASAP7_75t_R _30035_ (.A(_15818_),
    .B(_10647_),
    .Y(_10677_));
 AO21x1_ASAP7_75t_R _30036_ (.A1(_08110_),
    .A2(_10650_),
    .B(_10677_),
    .Y(_03581_));
 AND2x2_ASAP7_75t_R _30037_ (.A(_15939_),
    .B(_10647_),
    .Y(_10678_));
 AO21x1_ASAP7_75t_R _30038_ (.A1(_08151_),
    .A2(_10650_),
    .B(_10678_),
    .Y(_03582_));
 TAPCELL_ASAP7_75t_R PHY_342 ();
 AND2x2_ASAP7_75t_R _30040_ (.A(_16057_),
    .B(_10647_),
    .Y(_10680_));
 AO21x1_ASAP7_75t_R _30041_ (.A1(_08190_),
    .A2(_10650_),
    .B(_10680_),
    .Y(_03583_));
 TAPCELL_ASAP7_75t_R PHY_341 ();
 TAPCELL_ASAP7_75t_R PHY_340 ();
 AND2x2_ASAP7_75t_R _30044_ (.A(_16181_),
    .B(_10647_),
    .Y(_10683_));
 AO21x1_ASAP7_75t_R _30045_ (.A1(_08225_),
    .A2(_10650_),
    .B(_10683_),
    .Y(_03584_));
 TAPCELL_ASAP7_75t_R PHY_339 ();
 AND2x2_ASAP7_75t_R _30047_ (.A(_16268_),
    .B(_10647_),
    .Y(_10685_));
 AO21x1_ASAP7_75t_R _30048_ (.A1(_08263_),
    .A2(_10650_),
    .B(_10685_),
    .Y(_03585_));
 AND2x2_ASAP7_75t_R _30049_ (.A(_16450_),
    .B(_10647_),
    .Y(_10686_));
 AO21x1_ASAP7_75t_R _30050_ (.A1(_08294_),
    .A2(_10650_),
    .B(_10686_),
    .Y(_03586_));
 TAPCELL_ASAP7_75t_R PHY_338 ();
 AND2x2_ASAP7_75t_R _30052_ (.A(_16555_),
    .B(_10647_),
    .Y(_10688_));
 AO21x1_ASAP7_75t_R _30053_ (.A1(_08328_),
    .A2(_10650_),
    .B(_10688_),
    .Y(_03587_));
 TAPCELL_ASAP7_75t_R PHY_337 ();
 AND2x2_ASAP7_75t_R _30055_ (.A(_16651_),
    .B(_10647_),
    .Y(_10690_));
 AO21x1_ASAP7_75t_R _30056_ (.A1(_08360_),
    .A2(_10650_),
    .B(_10690_),
    .Y(_03588_));
 TAPCELL_ASAP7_75t_R PHY_336 ();
 AND2x2_ASAP7_75t_R _30058_ (.A(_04548_),
    .B(_10647_),
    .Y(_10692_));
 AO21x1_ASAP7_75t_R _30059_ (.A1(_08406_),
    .A2(_10650_),
    .B(_10692_),
    .Y(_03589_));
 AND2x2_ASAP7_75t_R _30060_ (.A(_04669_),
    .B(_10647_),
    .Y(_10693_));
 AO21x1_ASAP7_75t_R _30061_ (.A1(_08450_),
    .A2(_10650_),
    .B(_10693_),
    .Y(_03590_));
 TAPCELL_ASAP7_75t_R PHY_335 ();
 AND2x2_ASAP7_75t_R _30063_ (.A(_04780_),
    .B(_10647_),
    .Y(_10695_));
 AO21x1_ASAP7_75t_R _30064_ (.A1(_08481_),
    .A2(_10650_),
    .B(_10695_),
    .Y(_03591_));
 AND2x2_ASAP7_75t_R _30065_ (.A(_04895_),
    .B(_10647_),
    .Y(_10696_));
 AO21x1_ASAP7_75t_R _30066_ (.A1(_08509_),
    .A2(_10650_),
    .B(_10696_),
    .Y(_03592_));
 TAPCELL_ASAP7_75t_R PHY_334 ();
 AND2x2_ASAP7_75t_R _30068_ (.A(_04999_),
    .B(_10647_),
    .Y(_10698_));
 AO21x1_ASAP7_75t_R _30069_ (.A1(_08537_),
    .A2(_10650_),
    .B(_10698_),
    .Y(_03593_));
 AND2x2_ASAP7_75t_R _30070_ (.A(_05108_),
    .B(_10647_),
    .Y(_10699_));
 AO21x1_ASAP7_75t_R _30071_ (.A1(_08563_),
    .A2(_10650_),
    .B(_10699_),
    .Y(_03594_));
 TAPCELL_ASAP7_75t_R PHY_333 ();
 AND2x2_ASAP7_75t_R _30073_ (.A(_05238_),
    .B(_10647_),
    .Y(_10701_));
 AO21x1_ASAP7_75t_R _30074_ (.A1(net250),
    .A2(_10650_),
    .B(_10701_),
    .Y(_03595_));
 AND2x2_ASAP7_75t_R _30075_ (.A(_05327_),
    .B(_10647_),
    .Y(_10702_));
 AO21x1_ASAP7_75t_R _30076_ (.A1(net2197),
    .A2(_10650_),
    .B(_10702_),
    .Y(_03596_));
 AND2x2_ASAP7_75t_R _30077_ (.A(_08648_),
    .B(_10650_),
    .Y(_10703_));
 AOI21x1_ASAP7_75t_R _30078_ (.A1(_01298_),
    .A2(_10647_),
    .B(_10703_),
    .Y(_03597_));
 OR2x6_ASAP7_75t_R _30079_ (.A(_09914_),
    .B(_10514_),
    .Y(_10704_));
 TAPCELL_ASAP7_75t_R PHY_332 ();
 NOR2x1_ASAP7_75t_R _30081_ (.A(_07248_),
    .B(_10704_),
    .Y(_10706_));
 AO21x1_ASAP7_75t_R _30082_ (.A1(_13878_),
    .A2(_10704_),
    .B(_10706_),
    .Y(_03598_));
 NOR2x2_ASAP7_75t_R _30083_ (.A(_09914_),
    .B(_10514_),
    .Y(_10707_));
 TAPCELL_ASAP7_75t_R PHY_331 ();
 AND2x2_ASAP7_75t_R _30085_ (.A(_13348_),
    .B(_10704_),
    .Y(_10709_));
 AO21x1_ASAP7_75t_R _30086_ (.A1(_07384_),
    .A2(_10707_),
    .B(_10709_),
    .Y(_03599_));
 AND2x2_ASAP7_75t_R _30087_ (.A(_14118_),
    .B(_10704_),
    .Y(_10710_));
 AO21x1_ASAP7_75t_R _30088_ (.A1(_07472_),
    .A2(_10707_),
    .B(_10710_),
    .Y(_03600_));
 AND2x2_ASAP7_75t_R _30089_ (.A(_14200_),
    .B(_10704_),
    .Y(_10711_));
 AO21x1_ASAP7_75t_R _30090_ (.A1(_07552_),
    .A2(_10707_),
    .B(_10711_),
    .Y(_03601_));
 AND2x2_ASAP7_75t_R _30091_ (.A(_14995_),
    .B(_10704_),
    .Y(_10712_));
 AO21x1_ASAP7_75t_R _30092_ (.A1(_07608_),
    .A2(_10707_),
    .B(_10712_),
    .Y(_03602_));
 AND2x2_ASAP7_75t_R _30093_ (.A(_14305_),
    .B(_10704_),
    .Y(_10713_));
 AO21x1_ASAP7_75t_R _30094_ (.A1(_07663_),
    .A2(_10707_),
    .B(_10713_),
    .Y(_03603_));
 AND2x2_ASAP7_75t_R _30095_ (.A(_14398_),
    .B(_10704_),
    .Y(_10714_));
 AO21x1_ASAP7_75t_R _30096_ (.A1(_07709_),
    .A2(_10707_),
    .B(_10714_),
    .Y(_03604_));
 AND2x2_ASAP7_75t_R _30097_ (.A(_14453_),
    .B(_10704_),
    .Y(_10715_));
 AO21x1_ASAP7_75t_R _30098_ (.A1(net252),
    .A2(_10707_),
    .B(_10715_),
    .Y(_03605_));
 TAPCELL_ASAP7_75t_R PHY_330 ();
 AND2x2_ASAP7_75t_R _30100_ (.A(_14531_),
    .B(_10704_),
    .Y(_10717_));
 AO21x1_ASAP7_75t_R _30101_ (.A1(net257),
    .A2(_10707_),
    .B(_10717_),
    .Y(_03606_));
 AND2x2_ASAP7_75t_R _30102_ (.A(_14573_),
    .B(_10704_),
    .Y(_10718_));
 AO21x1_ASAP7_75t_R _30103_ (.A1(net256),
    .A2(_10707_),
    .B(_10718_),
    .Y(_03607_));
 AND2x2_ASAP7_75t_R _30104_ (.A(_14626_),
    .B(_10704_),
    .Y(_10719_));
 AO21x1_ASAP7_75t_R _30105_ (.A1(_07903_),
    .A2(_10707_),
    .B(_10719_),
    .Y(_03608_));
 TAPCELL_ASAP7_75t_R PHY_329 ();
 AND2x2_ASAP7_75t_R _30107_ (.A(_14726_),
    .B(_10704_),
    .Y(_10721_));
 AO21x1_ASAP7_75t_R _30108_ (.A1(_07948_),
    .A2(_10707_),
    .B(_10721_),
    .Y(_03609_));
 AND2x2_ASAP7_75t_R _30109_ (.A(_14040_),
    .B(_10704_),
    .Y(_10722_));
 AO21x1_ASAP7_75t_R _30110_ (.A1(_07985_),
    .A2(_10707_),
    .B(_10722_),
    .Y(_03610_));
 AND2x2_ASAP7_75t_R _30111_ (.A(_15564_),
    .B(_10704_),
    .Y(_10723_));
 AO21x1_ASAP7_75t_R _30112_ (.A1(_08026_),
    .A2(_10707_),
    .B(_10723_),
    .Y(_03611_));
 AND2x2_ASAP7_75t_R _30113_ (.A(_15692_),
    .B(_10704_),
    .Y(_10724_));
 AO21x1_ASAP7_75t_R _30114_ (.A1(_08068_),
    .A2(_10707_),
    .B(_10724_),
    .Y(_03612_));
 AND2x2_ASAP7_75t_R _30115_ (.A(_15815_),
    .B(_10704_),
    .Y(_10725_));
 AO21x1_ASAP7_75t_R _30116_ (.A1(_08110_),
    .A2(_10707_),
    .B(_10725_),
    .Y(_03613_));
 AND2x2_ASAP7_75t_R _30117_ (.A(_15936_),
    .B(_10704_),
    .Y(_10726_));
 AO21x1_ASAP7_75t_R _30118_ (.A1(_08151_),
    .A2(_10707_),
    .B(_10726_),
    .Y(_03614_));
 AND2x2_ASAP7_75t_R _30119_ (.A(_16053_),
    .B(_10704_),
    .Y(_10727_));
 AO21x1_ASAP7_75t_R _30120_ (.A1(_08190_),
    .A2(_10707_),
    .B(_10727_),
    .Y(_03615_));
 TAPCELL_ASAP7_75t_R PHY_328 ();
 AND2x2_ASAP7_75t_R _30122_ (.A(_16178_),
    .B(_10704_),
    .Y(_10729_));
 AO21x1_ASAP7_75t_R _30123_ (.A1(_08225_),
    .A2(_10707_),
    .B(_10729_),
    .Y(_03616_));
 AND2x2_ASAP7_75t_R _30124_ (.A(_16265_),
    .B(_10704_),
    .Y(_10730_));
 AO21x1_ASAP7_75t_R _30125_ (.A1(_08263_),
    .A2(_10707_),
    .B(_10730_),
    .Y(_03617_));
 AND2x2_ASAP7_75t_R _30126_ (.A(_16447_),
    .B(_10704_),
    .Y(_10731_));
 AO21x1_ASAP7_75t_R _30127_ (.A1(_08294_),
    .A2(_10707_),
    .B(_10731_),
    .Y(_03618_));
 TAPCELL_ASAP7_75t_R PHY_327 ();
 AND2x2_ASAP7_75t_R _30129_ (.A(_16552_),
    .B(_10704_),
    .Y(_10733_));
 AO21x1_ASAP7_75t_R _30130_ (.A1(_08328_),
    .A2(_10707_),
    .B(_10733_),
    .Y(_03619_));
 AND2x2_ASAP7_75t_R _30131_ (.A(_16648_),
    .B(_10704_),
    .Y(_10734_));
 AO21x1_ASAP7_75t_R _30132_ (.A1(_08360_),
    .A2(_10707_),
    .B(_10734_),
    .Y(_03620_));
 AND2x2_ASAP7_75t_R _30133_ (.A(_04545_),
    .B(_10704_),
    .Y(_10735_));
 AO21x1_ASAP7_75t_R _30134_ (.A1(_08406_),
    .A2(_10707_),
    .B(_10735_),
    .Y(_03621_));
 AND2x2_ASAP7_75t_R _30135_ (.A(_04666_),
    .B(_10704_),
    .Y(_10736_));
 AO21x1_ASAP7_75t_R _30136_ (.A1(_08450_),
    .A2(_10707_),
    .B(_10736_),
    .Y(_03622_));
 AND2x2_ASAP7_75t_R _30137_ (.A(_04777_),
    .B(_10704_),
    .Y(_10737_));
 AO21x1_ASAP7_75t_R _30138_ (.A1(_08481_),
    .A2(_10707_),
    .B(_10737_),
    .Y(_03623_));
 AND2x2_ASAP7_75t_R _30139_ (.A(_04892_),
    .B(_10704_),
    .Y(_10738_));
 AO21x1_ASAP7_75t_R _30140_ (.A1(_08509_),
    .A2(_10707_),
    .B(_10738_),
    .Y(_03624_));
 AND2x2_ASAP7_75t_R _30141_ (.A(_04996_),
    .B(_10704_),
    .Y(_10739_));
 AO21x1_ASAP7_75t_R _30142_ (.A1(_08537_),
    .A2(_10707_),
    .B(_10739_),
    .Y(_03625_));
 AND2x2_ASAP7_75t_R _30143_ (.A(_05105_),
    .B(_10704_),
    .Y(_10740_));
 AO21x1_ASAP7_75t_R _30144_ (.A1(_08563_),
    .A2(_10707_),
    .B(_10740_),
    .Y(_03626_));
 AND2x2_ASAP7_75t_R _30145_ (.A(_05235_),
    .B(_10704_),
    .Y(_10741_));
 AO21x1_ASAP7_75t_R _30146_ (.A1(net250),
    .A2(_10707_),
    .B(_10741_),
    .Y(_03627_));
 AND2x2_ASAP7_75t_R _30147_ (.A(_05324_),
    .B(_10704_),
    .Y(_10742_));
 AO21x1_ASAP7_75t_R _30148_ (.A1(net2197),
    .A2(_10707_),
    .B(_10742_),
    .Y(_03628_));
 AND2x2_ASAP7_75t_R _30149_ (.A(_08648_),
    .B(_10707_),
    .Y(_10743_));
 AOI21x1_ASAP7_75t_R _30150_ (.A1(_01299_),
    .A2(_10704_),
    .B(_10743_),
    .Y(_03629_));
 NAND2x2_ASAP7_75t_R _30151_ (.A(_10036_),
    .B(_10390_),
    .Y(_10744_));
 TAPCELL_ASAP7_75t_R PHY_326 ();
 AND2x6_ASAP7_75t_R _30153_ (.A(_10036_),
    .B(_10390_),
    .Y(_10746_));
 TAPCELL_ASAP7_75t_R PHY_325 ();
 AND2x2_ASAP7_75t_R _30155_ (.A(_07248_),
    .B(_10746_),
    .Y(_10748_));
 AOI21x1_ASAP7_75t_R _30156_ (.A1(_00315_),
    .A2(_10744_),
    .B(_10748_),
    .Y(_03630_));
 TAPCELL_ASAP7_75t_R PHY_324 ();
 TAPCELL_ASAP7_75t_R PHY_323 ();
 NOR2x1_ASAP7_75t_R _30159_ (.A(_00269_),
    .B(_10746_),
    .Y(_10751_));
 AO21x1_ASAP7_75t_R _30160_ (.A1(_07384_),
    .A2(_10746_),
    .B(_10751_),
    .Y(_03631_));
 TAPCELL_ASAP7_75t_R PHY_322 ();
 AND2x2_ASAP7_75t_R _30162_ (.A(_14908_),
    .B(_10744_),
    .Y(_10753_));
 AO21x1_ASAP7_75t_R _30163_ (.A1(_07472_),
    .A2(_10746_),
    .B(_10753_),
    .Y(_03632_));
 NOR2x1_ASAP7_75t_R _30164_ (.A(_00408_),
    .B(_10746_),
    .Y(_10754_));
 AO21x1_ASAP7_75t_R _30165_ (.A1(_07552_),
    .A2(_10746_),
    .B(_10754_),
    .Y(_03633_));
 NOR2x1_ASAP7_75t_R _30166_ (.A(_00438_),
    .B(_10746_),
    .Y(_10755_));
 AO21x1_ASAP7_75t_R _30167_ (.A1(_07608_),
    .A2(_10746_),
    .B(_10755_),
    .Y(_03634_));
 TAPCELL_ASAP7_75t_R PHY_321 ();
 NAND2x1_ASAP7_75t_R _30169_ (.A(_00468_),
    .B(_10744_),
    .Y(_10757_));
 OA21x2_ASAP7_75t_R _30170_ (.A1(_07663_),
    .A2(_10744_),
    .B(_10757_),
    .Y(_03635_));
 NOR2x1_ASAP7_75t_R _30171_ (.A(_00498_),
    .B(_10746_),
    .Y(_10758_));
 AO21x1_ASAP7_75t_R _30172_ (.A1(_07709_),
    .A2(_10746_),
    .B(_10758_),
    .Y(_03636_));
 NOR2x1_ASAP7_75t_R _30173_ (.A(_00528_),
    .B(_10746_),
    .Y(_10759_));
 AO21x1_ASAP7_75t_R _30174_ (.A1(net252),
    .A2(_10746_),
    .B(_10759_),
    .Y(_03637_));
 NAND2x1_ASAP7_75t_R _30175_ (.A(_00558_),
    .B(_10744_),
    .Y(_10760_));
 OA21x2_ASAP7_75t_R _30176_ (.A1(net257),
    .A2(_10744_),
    .B(_10760_),
    .Y(_03638_));
 NOR2x1_ASAP7_75t_R _30177_ (.A(_00588_),
    .B(_10746_),
    .Y(_10761_));
 AO21x1_ASAP7_75t_R _30178_ (.A1(_07866_),
    .A2(_10746_),
    .B(_10761_),
    .Y(_03639_));
 AND2x2_ASAP7_75t_R _30179_ (.A(_15383_),
    .B(_10744_),
    .Y(_10762_));
 AO21x1_ASAP7_75t_R _30180_ (.A1(_07903_),
    .A2(_10746_),
    .B(_10762_),
    .Y(_03640_));
 NOR2x1_ASAP7_75t_R _30181_ (.A(_00648_),
    .B(_10746_),
    .Y(_10763_));
 AO21x1_ASAP7_75t_R _30182_ (.A1(_07948_),
    .A2(_10746_),
    .B(_10763_),
    .Y(_03641_));
 NAND2x1_ASAP7_75t_R _30183_ (.A(_00347_),
    .B(_10744_),
    .Y(_10764_));
 OA21x2_ASAP7_75t_R _30184_ (.A1(_07985_),
    .A2(_10744_),
    .B(_10764_),
    .Y(_03642_));
 NAND2x1_ASAP7_75t_R _30185_ (.A(_00710_),
    .B(_10744_),
    .Y(_10765_));
 OA21x2_ASAP7_75t_R _30186_ (.A1(net251),
    .A2(_10744_),
    .B(_10765_),
    .Y(_03643_));
 AND2x2_ASAP7_75t_R _30187_ (.A(_15760_),
    .B(_10744_),
    .Y(_10766_));
 AO21x1_ASAP7_75t_R _30188_ (.A1(_08068_),
    .A2(_10746_),
    .B(_10766_),
    .Y(_03644_));
 NAND2x1_ASAP7_75t_R _30189_ (.A(_00775_),
    .B(_10744_),
    .Y(_10767_));
 OA21x2_ASAP7_75t_R _30190_ (.A1(_08110_),
    .A2(_10744_),
    .B(_10767_),
    .Y(_03645_));
 NAND2x1_ASAP7_75t_R _30191_ (.A(_00808_),
    .B(_10744_),
    .Y(_10768_));
 OA21x2_ASAP7_75t_R _30192_ (.A1(_08151_),
    .A2(_10744_),
    .B(_10768_),
    .Y(_03646_));
 AND2x2_ASAP7_75t_R _30193_ (.A(_16125_),
    .B(_10744_),
    .Y(_10769_));
 AO21x1_ASAP7_75t_R _30194_ (.A1(_08190_),
    .A2(_10746_),
    .B(_10769_),
    .Y(_03647_));
 AND2x2_ASAP7_75t_R _30195_ (.A(_16195_),
    .B(_10744_),
    .Y(_10770_));
 AO21x1_ASAP7_75t_R _30196_ (.A1(_08225_),
    .A2(_10746_),
    .B(_10770_),
    .Y(_03648_));
 AND2x2_ASAP7_75t_R _30197_ (.A(_16366_),
    .B(_10744_),
    .Y(_10771_));
 AO21x1_ASAP7_75t_R _30198_ (.A1(_08263_),
    .A2(_10746_),
    .B(_10771_),
    .Y(_03649_));
 NAND2x1_ASAP7_75t_R _30199_ (.A(_00938_),
    .B(_10744_),
    .Y(_10772_));
 OA21x2_ASAP7_75t_R _30200_ (.A1(_08294_),
    .A2(_10744_),
    .B(_10772_),
    .Y(_03650_));
 NOR2x1_ASAP7_75t_R _30201_ (.A(_00971_),
    .B(_10746_),
    .Y(_10773_));
 AO21x1_ASAP7_75t_R _30202_ (.A1(_08328_),
    .A2(_10746_),
    .B(_10773_),
    .Y(_03651_));
 NAND2x1_ASAP7_75t_R _30203_ (.A(_01003_),
    .B(_10744_),
    .Y(_10774_));
 OA21x2_ASAP7_75t_R _30204_ (.A1(_08360_),
    .A2(_10744_),
    .B(_10774_),
    .Y(_03652_));
 NOR2x1_ASAP7_75t_R _30205_ (.A(_01037_),
    .B(_10746_),
    .Y(_10775_));
 AO21x1_ASAP7_75t_R _30206_ (.A1(_08406_),
    .A2(_10746_),
    .B(_10775_),
    .Y(_03653_));
 NAND2x1_ASAP7_75t_R _30207_ (.A(_01069_),
    .B(_10744_),
    .Y(_10776_));
 OA21x2_ASAP7_75t_R _30208_ (.A1(_08450_),
    .A2(_10744_),
    .B(_10776_),
    .Y(_03654_));
 NOR2x1_ASAP7_75t_R _30209_ (.A(_01102_),
    .B(_10746_),
    .Y(_10777_));
 AO21x1_ASAP7_75t_R _30210_ (.A1(_08481_),
    .A2(_10746_),
    .B(_10777_),
    .Y(_03655_));
 NAND2x1_ASAP7_75t_R _30211_ (.A(_01134_),
    .B(_10744_),
    .Y(_10778_));
 OA21x2_ASAP7_75t_R _30212_ (.A1(_08509_),
    .A2(_10744_),
    .B(_10778_),
    .Y(_03656_));
 AND2x2_ASAP7_75t_R _30213_ (.A(_05011_),
    .B(_10744_),
    .Y(_10779_));
 AO21x1_ASAP7_75t_R _30214_ (.A1(_08537_),
    .A2(_10746_),
    .B(_10779_),
    .Y(_03657_));
 NAND2x1_ASAP7_75t_R _30215_ (.A(_01200_),
    .B(_10744_),
    .Y(_10780_));
 OA21x2_ASAP7_75t_R _30216_ (.A1(_08563_),
    .A2(_10744_),
    .B(_10780_),
    .Y(_03658_));
 AND2x2_ASAP7_75t_R _30217_ (.A(_05213_),
    .B(_10744_),
    .Y(_10781_));
 AO21x1_ASAP7_75t_R _30218_ (.A1(net250),
    .A2(_10746_),
    .B(_10781_),
    .Y(_03659_));
 NAND2x1_ASAP7_75t_R _30219_ (.A(_01266_),
    .B(_10744_),
    .Y(_10782_));
 OA21x2_ASAP7_75t_R _30220_ (.A1(net2197),
    .A2(_10744_),
    .B(_10782_),
    .Y(_03660_));
 AND2x2_ASAP7_75t_R _30221_ (.A(_08648_),
    .B(_10746_),
    .Y(_10783_));
 AOI21x1_ASAP7_75t_R _30222_ (.A1(_01300_),
    .A2(_10744_),
    .B(_10783_),
    .Y(_03661_));
 NOR2x2_ASAP7_75t_R _30223_ (.A(_10077_),
    .B(_10432_),
    .Y(_10784_));
 TAPCELL_ASAP7_75t_R PHY_320 ();
 TAPCELL_ASAP7_75t_R PHY_319 ();
 NAND2x1_ASAP7_75t_R _30226_ (.A(_07248_),
    .B(_10784_),
    .Y(_10787_));
 OA21x2_ASAP7_75t_R _30227_ (.A1(_13974_),
    .A2(_10784_),
    .B(_10787_),
    .Y(_03662_));
 NOR2x1_ASAP7_75t_R _30228_ (.A(_00270_),
    .B(net266),
    .Y(_10788_));
 AO21x1_ASAP7_75t_R _30229_ (.A1(_07384_),
    .A2(net266),
    .B(_10788_),
    .Y(_03663_));
 NOR2x1_ASAP7_75t_R _30230_ (.A(_00378_),
    .B(net265),
    .Y(_10789_));
 AO21x1_ASAP7_75t_R _30231_ (.A1(_07472_),
    .A2(net265),
    .B(_10789_),
    .Y(_03664_));
 NOR2x1_ASAP7_75t_R _30232_ (.A(_00409_),
    .B(_10784_),
    .Y(_10790_));
 AO21x1_ASAP7_75t_R _30233_ (.A1(_07552_),
    .A2(_10784_),
    .B(_10790_),
    .Y(_03665_));
 NOR2x1_ASAP7_75t_R _30234_ (.A(_00439_),
    .B(net265),
    .Y(_10791_));
 AO21x1_ASAP7_75t_R _30235_ (.A1(_07608_),
    .A2(net265),
    .B(_10791_),
    .Y(_03666_));
 NOR2x1_ASAP7_75t_R _30236_ (.A(_00469_),
    .B(net265),
    .Y(_10792_));
 AO21x1_ASAP7_75t_R _30237_ (.A1(_07663_),
    .A2(net265),
    .B(_10792_),
    .Y(_03667_));
 NOR2x1_ASAP7_75t_R _30238_ (.A(_00499_),
    .B(net265),
    .Y(_10793_));
 AO21x1_ASAP7_75t_R _30239_ (.A1(_07709_),
    .A2(net265),
    .B(_10793_),
    .Y(_03668_));
 NOR2x1_ASAP7_75t_R _30240_ (.A(_00529_),
    .B(net265),
    .Y(_10794_));
 AO21x1_ASAP7_75t_R _30241_ (.A1(net252),
    .A2(net265),
    .B(_10794_),
    .Y(_03669_));
 TAPCELL_ASAP7_75t_R PHY_318 ();
 NOR2x1_ASAP7_75t_R _30243_ (.A(_00559_),
    .B(net266),
    .Y(_10796_));
 AO21x1_ASAP7_75t_R _30244_ (.A1(_07825_),
    .A2(net266),
    .B(_10796_),
    .Y(_03670_));
 TAPCELL_ASAP7_75t_R PHY_317 ();
 NOR2x1_ASAP7_75t_R _30246_ (.A(_00589_),
    .B(net266),
    .Y(_10798_));
 AO21x1_ASAP7_75t_R _30247_ (.A1(_07866_),
    .A2(net266),
    .B(_10798_),
    .Y(_03671_));
 NOR2x1_ASAP7_75t_R _30248_ (.A(_00619_),
    .B(net265),
    .Y(_10799_));
 AO21x1_ASAP7_75t_R _30249_ (.A1(_07903_),
    .A2(net265),
    .B(_10799_),
    .Y(_03672_));
 NOR2x1_ASAP7_75t_R _30250_ (.A(_00649_),
    .B(net265),
    .Y(_10800_));
 AO21x1_ASAP7_75t_R _30251_ (.A1(_07948_),
    .A2(net265),
    .B(_10800_),
    .Y(_03673_));
 NOR2x1_ASAP7_75t_R _30252_ (.A(_00348_),
    .B(net265),
    .Y(_10801_));
 AO21x1_ASAP7_75t_R _30253_ (.A1(_07985_),
    .A2(net265),
    .B(_10801_),
    .Y(_03674_));
 NOR2x1_ASAP7_75t_R _30254_ (.A(_00711_),
    .B(net266),
    .Y(_10802_));
 AO21x1_ASAP7_75t_R _30255_ (.A1(net251),
    .A2(net266),
    .B(_10802_),
    .Y(_03675_));
 NOR2x1_ASAP7_75t_R _30256_ (.A(_00743_),
    .B(net265),
    .Y(_10803_));
 AO21x1_ASAP7_75t_R _30257_ (.A1(_08068_),
    .A2(net265),
    .B(_10803_),
    .Y(_03676_));
 NOR2x1_ASAP7_75t_R _30258_ (.A(_00776_),
    .B(_10784_),
    .Y(_10804_));
 AO21x1_ASAP7_75t_R _30259_ (.A1(_08110_),
    .A2(_10784_),
    .B(_10804_),
    .Y(_03677_));
 NOR2x1_ASAP7_75t_R _30260_ (.A(_00809_),
    .B(net265),
    .Y(_10805_));
 AO21x1_ASAP7_75t_R _30261_ (.A1(_08151_),
    .A2(net265),
    .B(_10805_),
    .Y(_03678_));
 NOR2x1_ASAP7_75t_R _30262_ (.A(_00842_),
    .B(net265),
    .Y(_10806_));
 AO21x1_ASAP7_75t_R _30263_ (.A1(_08190_),
    .A2(net265),
    .B(_10806_),
    .Y(_03679_));
 TAPCELL_ASAP7_75t_R PHY_316 ();
 NOR2x1_ASAP7_75t_R _30265_ (.A(_00874_),
    .B(_10784_),
    .Y(_10808_));
 AO21x1_ASAP7_75t_R _30266_ (.A1(_08225_),
    .A2(_10784_),
    .B(_10808_),
    .Y(_03680_));
 TAPCELL_ASAP7_75t_R PHY_315 ();
 NOR2x1_ASAP7_75t_R _30268_ (.A(_00907_),
    .B(net265),
    .Y(_10810_));
 AO21x1_ASAP7_75t_R _30269_ (.A1(_08263_),
    .A2(net265),
    .B(_10810_),
    .Y(_03681_));
 NOR2x1_ASAP7_75t_R _30270_ (.A(_00939_),
    .B(_10784_),
    .Y(_10811_));
 AO21x1_ASAP7_75t_R _30271_ (.A1(_08294_),
    .A2(_10784_),
    .B(_10811_),
    .Y(_03682_));
 NOR2x1_ASAP7_75t_R _30272_ (.A(_00972_),
    .B(net265),
    .Y(_10812_));
 AO21x1_ASAP7_75t_R _30273_ (.A1(_08328_),
    .A2(net265),
    .B(_10812_),
    .Y(_03683_));
 NOR2x1_ASAP7_75t_R _30274_ (.A(_01004_),
    .B(_10784_),
    .Y(_10813_));
 AO21x1_ASAP7_75t_R _30275_ (.A1(_08360_),
    .A2(_10784_),
    .B(_10813_),
    .Y(_03684_));
 NOR2x1_ASAP7_75t_R _30276_ (.A(_01038_),
    .B(net266),
    .Y(_10814_));
 AO21x1_ASAP7_75t_R _30277_ (.A1(_08406_),
    .A2(net266),
    .B(_10814_),
    .Y(_03685_));
 NOR2x1_ASAP7_75t_R _30278_ (.A(_01070_),
    .B(_10784_),
    .Y(_10815_));
 AO21x1_ASAP7_75t_R _30279_ (.A1(_08450_),
    .A2(_10784_),
    .B(_10815_),
    .Y(_03686_));
 NOR2x1_ASAP7_75t_R _30280_ (.A(_01103_),
    .B(net265),
    .Y(_10816_));
 AO21x1_ASAP7_75t_R _30281_ (.A1(_08481_),
    .A2(net265),
    .B(_10816_),
    .Y(_03687_));
 NOR2x1_ASAP7_75t_R _30282_ (.A(_01135_),
    .B(net266),
    .Y(_10817_));
 AO21x1_ASAP7_75t_R _30283_ (.A1(_08509_),
    .A2(net266),
    .B(_10817_),
    .Y(_03688_));
 NOR2x1_ASAP7_75t_R _30284_ (.A(_01169_),
    .B(net266),
    .Y(_10818_));
 AO21x1_ASAP7_75t_R _30285_ (.A1(_08537_),
    .A2(net266),
    .B(_10818_),
    .Y(_03689_));
 NOR2x1_ASAP7_75t_R _30286_ (.A(_01201_),
    .B(net266),
    .Y(_10819_));
 AO21x1_ASAP7_75t_R _30287_ (.A1(_08563_),
    .A2(net266),
    .B(_10819_),
    .Y(_03690_));
 NOR2x1_ASAP7_75t_R _30288_ (.A(_01235_),
    .B(net265),
    .Y(_10820_));
 AO21x1_ASAP7_75t_R _30289_ (.A1(net250),
    .A2(net265),
    .B(_10820_),
    .Y(_03691_));
 NOR2x1_ASAP7_75t_R _30290_ (.A(_01267_),
    .B(net266),
    .Y(_10821_));
 AO21x1_ASAP7_75t_R _30291_ (.A1(net2197),
    .A2(net266),
    .B(_10821_),
    .Y(_03692_));
 OR3x1_ASAP7_75t_R _30292_ (.A(_08648_),
    .B(_10077_),
    .C(_10432_),
    .Y(_10822_));
 OAI21x1_ASAP7_75t_R _30293_ (.A1(_01301_),
    .A2(net266),
    .B(_10822_),
    .Y(_03693_));
 NAND2x2_ASAP7_75t_R _30294_ (.A(_10036_),
    .B(_10473_),
    .Y(_10823_));
 TAPCELL_ASAP7_75t_R PHY_314 ();
 NOR2x1_ASAP7_75t_R _30296_ (.A(_07248_),
    .B(_10823_),
    .Y(_10825_));
 AO21x1_ASAP7_75t_R _30297_ (.A1(_13859_),
    .A2(_10823_),
    .B(_10825_),
    .Y(_03694_));
 NAND2x1_ASAP7_75t_R _30298_ (.A(_00271_),
    .B(_10823_),
    .Y(_10826_));
 OA21x2_ASAP7_75t_R _30299_ (.A1(_07384_),
    .A2(_10823_),
    .B(_10826_),
    .Y(_03695_));
 AND2x6_ASAP7_75t_R _30300_ (.A(_10036_),
    .B(_10473_),
    .Y(_10827_));
 TAPCELL_ASAP7_75t_R PHY_313 ();
 TAPCELL_ASAP7_75t_R PHY_312 ();
 NOR2x1_ASAP7_75t_R _30303_ (.A(_00379_),
    .B(_10827_),
    .Y(_10830_));
 AO21x1_ASAP7_75t_R _30304_ (.A1(_07472_),
    .A2(_10827_),
    .B(_10830_),
    .Y(_03696_));
 AND2x2_ASAP7_75t_R _30305_ (.A(_14956_),
    .B(_10823_),
    .Y(_10831_));
 AO21x1_ASAP7_75t_R _30306_ (.A1(_07552_),
    .A2(_10827_),
    .B(_10831_),
    .Y(_03697_));
 AND2x2_ASAP7_75t_R _30307_ (.A(_14280_),
    .B(_10823_),
    .Y(_10832_));
 AO21x1_ASAP7_75t_R _30308_ (.A1(_07608_),
    .A2(_10827_),
    .B(_10832_),
    .Y(_03698_));
 AND2x2_ASAP7_75t_R _30309_ (.A(_14322_),
    .B(_10823_),
    .Y(_10833_));
 AO21x1_ASAP7_75t_R _30310_ (.A1(_07663_),
    .A2(_10827_),
    .B(_10833_),
    .Y(_03699_));
 TAPCELL_ASAP7_75t_R PHY_311 ();
 TAPCELL_ASAP7_75t_R PHY_310 ();
 AND2x2_ASAP7_75t_R _30313_ (.A(_14415_),
    .B(_10823_),
    .Y(_10836_));
 AO21x1_ASAP7_75t_R _30314_ (.A1(_07709_),
    .A2(_10827_),
    .B(_10836_),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _30315_ (.A(_00530_),
    .B(_10827_),
    .Y(_10837_));
 AO21x1_ASAP7_75t_R _30316_ (.A1(net252),
    .A2(_10827_),
    .B(_10837_),
    .Y(_03701_));
 AND2x2_ASAP7_75t_R _30317_ (.A(_14513_),
    .B(_10823_),
    .Y(_10838_));
 AO21x1_ASAP7_75t_R _30318_ (.A1(net257),
    .A2(_10827_),
    .B(_10838_),
    .Y(_03702_));
 AND2x2_ASAP7_75t_R _30319_ (.A(_14588_),
    .B(_10823_),
    .Y(_10839_));
 AO21x1_ASAP7_75t_R _30320_ (.A1(_07866_),
    .A2(_10827_),
    .B(_10839_),
    .Y(_03703_));
 NOR2x1_ASAP7_75t_R _30321_ (.A(_00620_),
    .B(_10827_),
    .Y(_10840_));
 AO21x1_ASAP7_75t_R _30322_ (.A1(_07903_),
    .A2(_10827_),
    .B(_10840_),
    .Y(_03704_));
 AND2x2_ASAP7_75t_R _30323_ (.A(_14678_),
    .B(_10823_),
    .Y(_10841_));
 AO21x1_ASAP7_75t_R _30324_ (.A1(_07948_),
    .A2(_10827_),
    .B(_10841_),
    .Y(_03705_));
 AND3x1_ASAP7_75t_R _30325_ (.A(_07961_),
    .B(_07984_),
    .C(_10827_),
    .Y(_10842_));
 AO21x1_ASAP7_75t_R _30326_ (.A1(_14093_),
    .A2(_10823_),
    .B(_10842_),
    .Y(_03706_));
 TAPCELL_ASAP7_75t_R PHY_309 ();
 AND2x2_ASAP7_75t_R _30328_ (.A(_15573_),
    .B(_10823_),
    .Y(_10844_));
 AO21x1_ASAP7_75t_R _30329_ (.A1(net251),
    .A2(_10827_),
    .B(_10844_),
    .Y(_03707_));
 AND2x2_ASAP7_75t_R _30330_ (.A(_15707_),
    .B(_10823_),
    .Y(_10845_));
 AO21x1_ASAP7_75t_R _30331_ (.A1(_08068_),
    .A2(_10827_),
    .B(_10845_),
    .Y(_03708_));
 AND2x2_ASAP7_75t_R _30332_ (.A(_15833_),
    .B(_10823_),
    .Y(_10846_));
 AO21x1_ASAP7_75t_R _30333_ (.A1(_08110_),
    .A2(_10827_),
    .B(_10846_),
    .Y(_03709_));
 AND2x2_ASAP7_75t_R _30334_ (.A(_15966_),
    .B(_10823_),
    .Y(_10847_));
 AO21x1_ASAP7_75t_R _30335_ (.A1(_08151_),
    .A2(_10827_),
    .B(_10847_),
    .Y(_03710_));
 AND2x2_ASAP7_75t_R _30336_ (.A(_16070_),
    .B(_10823_),
    .Y(_10848_));
 AO21x1_ASAP7_75t_R _30337_ (.A1(_08190_),
    .A2(_10827_),
    .B(_10848_),
    .Y(_03711_));
 NOR2x1_ASAP7_75t_R _30338_ (.A(_00875_),
    .B(_10827_),
    .Y(_10849_));
 AO21x1_ASAP7_75t_R _30339_ (.A1(_08225_),
    .A2(_10827_),
    .B(_10849_),
    .Y(_03712_));
 AND2x2_ASAP7_75t_R _30340_ (.A(_16280_),
    .B(_10823_),
    .Y(_10850_));
 AO21x1_ASAP7_75t_R _30341_ (.A1(_08263_),
    .A2(_10827_),
    .B(_10850_),
    .Y(_03713_));
 AND2x2_ASAP7_75t_R _30342_ (.A(_16434_),
    .B(_10823_),
    .Y(_10851_));
 AO21x1_ASAP7_75t_R _30343_ (.A1(_08294_),
    .A2(_10827_),
    .B(_10851_),
    .Y(_03714_));
 AND2x2_ASAP7_75t_R _30344_ (.A(_16540_),
    .B(_10823_),
    .Y(_10852_));
 AO21x1_ASAP7_75t_R _30345_ (.A1(_08328_),
    .A2(_10827_),
    .B(_10852_),
    .Y(_03715_));
 AND2x2_ASAP7_75t_R _30346_ (.A(_16673_),
    .B(_10823_),
    .Y(_10853_));
 AO21x1_ASAP7_75t_R _30347_ (.A1(_08360_),
    .A2(_10827_),
    .B(_10853_),
    .Y(_03716_));
 AND2x2_ASAP7_75t_R _30348_ (.A(_04563_),
    .B(_10823_),
    .Y(_10854_));
 AO21x1_ASAP7_75t_R _30349_ (.A1(_08406_),
    .A2(_10827_),
    .B(_10854_),
    .Y(_03717_));
 AND2x2_ASAP7_75t_R _30350_ (.A(_04691_),
    .B(_10823_),
    .Y(_10855_));
 AO21x1_ASAP7_75t_R _30351_ (.A1(_08450_),
    .A2(_10827_),
    .B(_10855_),
    .Y(_03718_));
 AND2x2_ASAP7_75t_R _30352_ (.A(_04795_),
    .B(_10823_),
    .Y(_10856_));
 AO21x1_ASAP7_75t_R _30353_ (.A1(_08481_),
    .A2(_10827_),
    .B(_10856_),
    .Y(_03719_));
 AND2x2_ASAP7_75t_R _30354_ (.A(_04903_),
    .B(_10823_),
    .Y(_10857_));
 AO21x1_ASAP7_75t_R _30355_ (.A1(_08509_),
    .A2(_10827_),
    .B(_10857_),
    .Y(_03720_));
 NOR2x1_ASAP7_75t_R _30356_ (.A(_01170_),
    .B(_10827_),
    .Y(_10858_));
 AO21x1_ASAP7_75t_R _30357_ (.A1(_08537_),
    .A2(_10827_),
    .B(_10858_),
    .Y(_03721_));
 AND2x2_ASAP7_75t_R _30358_ (.A(_05130_),
    .B(_10823_),
    .Y(_10859_));
 AO21x1_ASAP7_75t_R _30359_ (.A1(_08563_),
    .A2(_10827_),
    .B(_10859_),
    .Y(_03722_));
 NOR2x1_ASAP7_75t_R _30360_ (.A(_01236_),
    .B(_10827_),
    .Y(_10860_));
 AO21x1_ASAP7_75t_R _30361_ (.A1(net250),
    .A2(_10827_),
    .B(_10860_),
    .Y(_03723_));
 AND2x2_ASAP7_75t_R _30362_ (.A(_05342_),
    .B(_10823_),
    .Y(_10861_));
 AO21x1_ASAP7_75t_R _30363_ (.A1(net2197),
    .A2(_10827_),
    .B(_10861_),
    .Y(_03724_));
 NOR2x1_ASAP7_75t_R _30364_ (.A(_08648_),
    .B(_10823_),
    .Y(_10862_));
 AO21x1_ASAP7_75t_R _30365_ (.A1(_05501_),
    .A2(_10823_),
    .B(_10862_),
    .Y(_03725_));
 OR2x6_ASAP7_75t_R _30366_ (.A(_10077_),
    .B(_10514_),
    .Y(_10863_));
 TAPCELL_ASAP7_75t_R PHY_308 ();
 NOR2x1_ASAP7_75t_R _30368_ (.A(_07248_),
    .B(_10863_),
    .Y(_10865_));
 AO21x1_ASAP7_75t_R _30369_ (.A1(_13867_),
    .A2(_10863_),
    .B(_10865_),
    .Y(_03726_));
 NOR2x2_ASAP7_75t_R _30370_ (.A(_10077_),
    .B(_10514_),
    .Y(_10866_));
 TAPCELL_ASAP7_75t_R PHY_307 ();
 AND2x2_ASAP7_75t_R _30372_ (.A(_13758_),
    .B(_10863_),
    .Y(_10868_));
 AO21x1_ASAP7_75t_R _30373_ (.A1(_07384_),
    .A2(_10866_),
    .B(_10868_),
    .Y(_03727_));
 AND2x2_ASAP7_75t_R _30374_ (.A(_14127_),
    .B(_10863_),
    .Y(_10869_));
 AO21x1_ASAP7_75t_R _30375_ (.A1(_07472_),
    .A2(_10866_),
    .B(_10869_),
    .Y(_03728_));
 AND2x2_ASAP7_75t_R _30376_ (.A(_14952_),
    .B(_10863_),
    .Y(_10870_));
 AO21x1_ASAP7_75t_R _30377_ (.A1(_07552_),
    .A2(_10866_),
    .B(_10870_),
    .Y(_03729_));
 AND2x2_ASAP7_75t_R _30378_ (.A(_15038_),
    .B(_10863_),
    .Y(_10871_));
 AO21x1_ASAP7_75t_R _30379_ (.A1(_07608_),
    .A2(_10866_),
    .B(_10871_),
    .Y(_03730_));
 AND2x2_ASAP7_75t_R _30380_ (.A(_14316_),
    .B(_10863_),
    .Y(_10872_));
 AO21x1_ASAP7_75t_R _30381_ (.A1(_07663_),
    .A2(_10866_),
    .B(_10872_),
    .Y(_03731_));
 AND2x2_ASAP7_75t_R _30382_ (.A(_14412_),
    .B(_10863_),
    .Y(_10873_));
 AO21x1_ASAP7_75t_R _30383_ (.A1(_07709_),
    .A2(_10866_),
    .B(_10873_),
    .Y(_03732_));
 NOR2x1_ASAP7_75t_R _30384_ (.A(_00531_),
    .B(_10866_),
    .Y(_10874_));
 AO21x1_ASAP7_75t_R _30385_ (.A1(net252),
    .A2(_10866_),
    .B(_10874_),
    .Y(_03733_));
 TAPCELL_ASAP7_75t_R PHY_306 ();
 AND2x2_ASAP7_75t_R _30387_ (.A(_14520_),
    .B(_10863_),
    .Y(_10876_));
 AO21x1_ASAP7_75t_R _30388_ (.A1(_07825_),
    .A2(_10866_),
    .B(_10876_),
    .Y(_03734_));
 AND2x2_ASAP7_75t_R _30389_ (.A(_15317_),
    .B(_10863_),
    .Y(_10877_));
 AO21x1_ASAP7_75t_R _30390_ (.A1(net256),
    .A2(_10866_),
    .B(_10877_),
    .Y(_03735_));
 AND2x2_ASAP7_75t_R _30391_ (.A(_15389_),
    .B(_10863_),
    .Y(_10878_));
 AO21x1_ASAP7_75t_R _30392_ (.A1(_07903_),
    .A2(_10866_),
    .B(_10878_),
    .Y(_03736_));
 TAPCELL_ASAP7_75t_R PHY_305 ();
 NOR2x1_ASAP7_75t_R _30394_ (.A(_00651_),
    .B(_10866_),
    .Y(_10880_));
 AO21x1_ASAP7_75t_R _30395_ (.A1(_07948_),
    .A2(_10866_),
    .B(_10880_),
    .Y(_03737_));
 AND2x2_ASAP7_75t_R _30396_ (.A(_14082_),
    .B(_10863_),
    .Y(_10881_));
 AO21x1_ASAP7_75t_R _30397_ (.A1(_07985_),
    .A2(_10866_),
    .B(_10881_),
    .Y(_03738_));
 AND2x2_ASAP7_75t_R _30398_ (.A(_15577_),
    .B(_10863_),
    .Y(_10882_));
 AO21x1_ASAP7_75t_R _30399_ (.A1(net251),
    .A2(_10866_),
    .B(_10882_),
    .Y(_03739_));
 AND2x2_ASAP7_75t_R _30400_ (.A(_15710_),
    .B(_10863_),
    .Y(_10883_));
 AO21x1_ASAP7_75t_R _30401_ (.A1(_08068_),
    .A2(_10866_),
    .B(_10883_),
    .Y(_03740_));
 AND2x2_ASAP7_75t_R _30402_ (.A(_15830_),
    .B(_10863_),
    .Y(_10884_));
 AO21x1_ASAP7_75t_R _30403_ (.A1(_08110_),
    .A2(_10866_),
    .B(_10884_),
    .Y(_03741_));
 AND2x2_ASAP7_75t_R _30404_ (.A(_15963_),
    .B(_10863_),
    .Y(_10885_));
 AO21x1_ASAP7_75t_R _30405_ (.A1(_08151_),
    .A2(_10866_),
    .B(_10885_),
    .Y(_03742_));
 AND2x2_ASAP7_75t_R _30406_ (.A(_16073_),
    .B(_10863_),
    .Y(_10886_));
 AO21x1_ASAP7_75t_R _30407_ (.A1(_08190_),
    .A2(_10866_),
    .B(_10886_),
    .Y(_03743_));
 AND2x2_ASAP7_75t_R _30408_ (.A(_16200_),
    .B(_10863_),
    .Y(_10887_));
 AO21x1_ASAP7_75t_R _30409_ (.A1(_08225_),
    .A2(_10866_),
    .B(_10887_),
    .Y(_03744_));
 TAPCELL_ASAP7_75t_R PHY_304 ();
 AND2x2_ASAP7_75t_R _30411_ (.A(_16283_),
    .B(_10863_),
    .Y(_10889_));
 AO21x1_ASAP7_75t_R _30412_ (.A1(_08263_),
    .A2(_10866_),
    .B(_10889_),
    .Y(_03745_));
 AND2x2_ASAP7_75t_R _30413_ (.A(_16431_),
    .B(_10863_),
    .Y(_10890_));
 AO21x1_ASAP7_75t_R _30414_ (.A1(_08294_),
    .A2(_10866_),
    .B(_10890_),
    .Y(_03746_));
 TAPCELL_ASAP7_75t_R PHY_303 ();
 AND2x2_ASAP7_75t_R _30416_ (.A(_16537_),
    .B(_10863_),
    .Y(_10892_));
 AO21x1_ASAP7_75t_R _30417_ (.A1(_08328_),
    .A2(_10866_),
    .B(_10892_),
    .Y(_03747_));
 AND2x2_ASAP7_75t_R _30418_ (.A(_16670_),
    .B(_10863_),
    .Y(_10893_));
 AO21x1_ASAP7_75t_R _30419_ (.A1(_08360_),
    .A2(_10866_),
    .B(_10893_),
    .Y(_03748_));
 AND2x2_ASAP7_75t_R _30420_ (.A(_04560_),
    .B(_10863_),
    .Y(_10894_));
 AO21x1_ASAP7_75t_R _30421_ (.A1(_08406_),
    .A2(_10866_),
    .B(_10894_),
    .Y(_03749_));
 AND2x2_ASAP7_75t_R _30422_ (.A(_04688_),
    .B(_10863_),
    .Y(_10895_));
 AO21x1_ASAP7_75t_R _30423_ (.A1(_08450_),
    .A2(_10866_),
    .B(_10895_),
    .Y(_03750_));
 AND2x2_ASAP7_75t_R _30424_ (.A(_04792_),
    .B(_10863_),
    .Y(_10896_));
 AO21x1_ASAP7_75t_R _30425_ (.A1(_08481_),
    .A2(_10866_),
    .B(_10896_),
    .Y(_03751_));
 AND2x2_ASAP7_75t_R _30426_ (.A(_04900_),
    .B(_10863_),
    .Y(_10897_));
 AO21x1_ASAP7_75t_R _30427_ (.A1(_08509_),
    .A2(_10866_),
    .B(_10897_),
    .Y(_03752_));
 AND2x2_ASAP7_75t_R _30428_ (.A(_05014_),
    .B(_10863_),
    .Y(_10898_));
 AO21x1_ASAP7_75t_R _30429_ (.A1(_08537_),
    .A2(_10866_),
    .B(_10898_),
    .Y(_03753_));
 AND2x2_ASAP7_75t_R _30430_ (.A(_05127_),
    .B(_10863_),
    .Y(_10899_));
 AO21x1_ASAP7_75t_R _30431_ (.A1(_08563_),
    .A2(_10866_),
    .B(_10899_),
    .Y(_03754_));
 AND2x2_ASAP7_75t_R _30432_ (.A(_05216_),
    .B(_10863_),
    .Y(_10900_));
 AO21x1_ASAP7_75t_R _30433_ (.A1(net250),
    .A2(_10866_),
    .B(_10900_),
    .Y(_03755_));
 AND2x2_ASAP7_75t_R _30434_ (.A(_05339_),
    .B(_10863_),
    .Y(_10901_));
 AO21x1_ASAP7_75t_R _30435_ (.A1(net2197),
    .A2(_10866_),
    .B(_10901_),
    .Y(_03756_));
 NOR2x1_ASAP7_75t_R _30436_ (.A(_08648_),
    .B(_10863_),
    .Y(_10902_));
 AO21x1_ASAP7_75t_R _30437_ (.A1(_05498_),
    .A2(_10863_),
    .B(_10902_),
    .Y(_03757_));
 INVx1_ASAP7_75t_R _30438_ (.A(_00319_),
    .Y(_10903_));
 AND2x6_ASAP7_75t_R _30439_ (.A(_10213_),
    .B(_10390_),
    .Y(_10904_));
 TAPCELL_ASAP7_75t_R PHY_302 ();
 TAPCELL_ASAP7_75t_R PHY_301 ();
 TAPCELL_ASAP7_75t_R PHY_300 ();
 NAND2x1_ASAP7_75t_R _30443_ (.A(_07248_),
    .B(_10904_),
    .Y(_10908_));
 OA21x2_ASAP7_75t_R _30444_ (.A1(_10903_),
    .A2(_10904_),
    .B(_10908_),
    .Y(_03758_));
 NOR2x1_ASAP7_75t_R _30445_ (.A(_00273_),
    .B(_10904_),
    .Y(_10909_));
 AO21x1_ASAP7_75t_R _30446_ (.A1(_07384_),
    .A2(_10904_),
    .B(_10909_),
    .Y(_03759_));
 NOR2x1_ASAP7_75t_R _30447_ (.A(_00381_),
    .B(_10904_),
    .Y(_10910_));
 AO21x1_ASAP7_75t_R _30448_ (.A1(_07472_),
    .A2(_10904_),
    .B(_10910_),
    .Y(_03760_));
 NOR2x1_ASAP7_75t_R _30449_ (.A(_00412_),
    .B(_10904_),
    .Y(_10911_));
 AO21x1_ASAP7_75t_R _30450_ (.A1(_07552_),
    .A2(_10904_),
    .B(_10911_),
    .Y(_03761_));
 NOR2x1_ASAP7_75t_R _30451_ (.A(_00442_),
    .B(_10904_),
    .Y(_10912_));
 AO21x1_ASAP7_75t_R _30452_ (.A1(_07608_),
    .A2(_10904_),
    .B(_10912_),
    .Y(_03762_));
 NOR2x1_ASAP7_75t_R _30453_ (.A(_00472_),
    .B(_10904_),
    .Y(_10913_));
 AO21x1_ASAP7_75t_R _30454_ (.A1(_07663_),
    .A2(_10904_),
    .B(_10913_),
    .Y(_03763_));
 NOR2x1_ASAP7_75t_R _30455_ (.A(_00502_),
    .B(_10904_),
    .Y(_10914_));
 AO21x1_ASAP7_75t_R _30456_ (.A1(_07709_),
    .A2(_10904_),
    .B(_10914_),
    .Y(_03764_));
 TAPCELL_ASAP7_75t_R PHY_299 ();
 NOR2x1_ASAP7_75t_R _30458_ (.A(_00532_),
    .B(_10904_),
    .Y(_10916_));
 AO21x1_ASAP7_75t_R _30459_ (.A1(_07760_),
    .A2(_10904_),
    .B(_10916_),
    .Y(_03765_));
 NOR2x1_ASAP7_75t_R _30460_ (.A(_00562_),
    .B(_10904_),
    .Y(_10917_));
 AO21x1_ASAP7_75t_R _30461_ (.A1(net257),
    .A2(_10904_),
    .B(_10917_),
    .Y(_03766_));
 TAPCELL_ASAP7_75t_R PHY_298 ();
 NOR2x1_ASAP7_75t_R _30463_ (.A(_00592_),
    .B(_10904_),
    .Y(_10919_));
 AO21x1_ASAP7_75t_R _30464_ (.A1(net256),
    .A2(_10904_),
    .B(_10919_),
    .Y(_03767_));
 NOR2x1_ASAP7_75t_R _30465_ (.A(_00622_),
    .B(_10904_),
    .Y(_10920_));
 AO21x1_ASAP7_75t_R _30466_ (.A1(_07903_),
    .A2(_10904_),
    .B(_10920_),
    .Y(_03768_));
 NOR2x1_ASAP7_75t_R _30467_ (.A(_00652_),
    .B(_10904_),
    .Y(_10921_));
 AO21x1_ASAP7_75t_R _30468_ (.A1(_07948_),
    .A2(_10904_),
    .B(_10921_),
    .Y(_03769_));
 NOR2x1_ASAP7_75t_R _30469_ (.A(_00351_),
    .B(_10904_),
    .Y(_10922_));
 AO21x1_ASAP7_75t_R _30470_ (.A1(_07985_),
    .A2(_10904_),
    .B(_10922_),
    .Y(_03770_));
 NOR2x1_ASAP7_75t_R _30471_ (.A(_00714_),
    .B(_10904_),
    .Y(_10923_));
 AO21x1_ASAP7_75t_R _30472_ (.A1(net251),
    .A2(_10904_),
    .B(_10923_),
    .Y(_03771_));
 NOR2x1_ASAP7_75t_R _30473_ (.A(_00746_),
    .B(_10904_),
    .Y(_10924_));
 AO21x1_ASAP7_75t_R _30474_ (.A1(_08068_),
    .A2(_10904_),
    .B(_10924_),
    .Y(_03772_));
 NOR2x1_ASAP7_75t_R _30475_ (.A(_00779_),
    .B(_10904_),
    .Y(_10925_));
 AO21x1_ASAP7_75t_R _30476_ (.A1(_08110_),
    .A2(_10904_),
    .B(_10925_),
    .Y(_03773_));
 NOR2x1_ASAP7_75t_R _30477_ (.A(_00812_),
    .B(_10904_),
    .Y(_10926_));
 AO21x1_ASAP7_75t_R _30478_ (.A1(_08151_),
    .A2(_10904_),
    .B(_10926_),
    .Y(_03774_));
 TAPCELL_ASAP7_75t_R PHY_297 ();
 NOR2x1_ASAP7_75t_R _30480_ (.A(_00845_),
    .B(_10904_),
    .Y(_10928_));
 AO21x1_ASAP7_75t_R _30481_ (.A1(_08190_),
    .A2(_10904_),
    .B(_10928_),
    .Y(_03775_));
 NOR2x1_ASAP7_75t_R _30482_ (.A(_00877_),
    .B(_10904_),
    .Y(_10929_));
 AO21x1_ASAP7_75t_R _30483_ (.A1(_08225_),
    .A2(_10904_),
    .B(_10929_),
    .Y(_03776_));
 TAPCELL_ASAP7_75t_R PHY_296 ();
 NOR2x1_ASAP7_75t_R _30485_ (.A(_00910_),
    .B(_10904_),
    .Y(_10931_));
 AO21x1_ASAP7_75t_R _30486_ (.A1(_08263_),
    .A2(_10904_),
    .B(_10931_),
    .Y(_03777_));
 NOR2x1_ASAP7_75t_R _30487_ (.A(_00942_),
    .B(_10904_),
    .Y(_10932_));
 AO21x1_ASAP7_75t_R _30488_ (.A1(_08294_),
    .A2(_10904_),
    .B(_10932_),
    .Y(_03778_));
 NOR2x1_ASAP7_75t_R _30489_ (.A(_00975_),
    .B(_10904_),
    .Y(_10933_));
 AO21x1_ASAP7_75t_R _30490_ (.A1(_08328_),
    .A2(_10904_),
    .B(_10933_),
    .Y(_03779_));
 NOR2x1_ASAP7_75t_R _30491_ (.A(_01007_),
    .B(_10904_),
    .Y(_10934_));
 AO21x1_ASAP7_75t_R _30492_ (.A1(_08360_),
    .A2(_10904_),
    .B(_10934_),
    .Y(_03780_));
 NOR2x1_ASAP7_75t_R _30493_ (.A(_01041_),
    .B(_10904_),
    .Y(_10935_));
 AO21x1_ASAP7_75t_R _30494_ (.A1(_08406_),
    .A2(_10904_),
    .B(_10935_),
    .Y(_03781_));
 NOR2x1_ASAP7_75t_R _30495_ (.A(_01073_),
    .B(_10904_),
    .Y(_10936_));
 AO21x1_ASAP7_75t_R _30496_ (.A1(_08450_),
    .A2(_10904_),
    .B(_10936_),
    .Y(_03782_));
 NOR2x1_ASAP7_75t_R _30497_ (.A(_01106_),
    .B(_10904_),
    .Y(_10937_));
 AO21x1_ASAP7_75t_R _30498_ (.A1(_08481_),
    .A2(_10904_),
    .B(_10937_),
    .Y(_03783_));
 NOR2x1_ASAP7_75t_R _30499_ (.A(_01138_),
    .B(_10904_),
    .Y(_10938_));
 AO21x1_ASAP7_75t_R _30500_ (.A1(_08509_),
    .A2(_10904_),
    .B(_10938_),
    .Y(_03784_));
 NOR2x1_ASAP7_75t_R _30501_ (.A(_01172_),
    .B(_10904_),
    .Y(_10939_));
 AO21x1_ASAP7_75t_R _30502_ (.A1(_08537_),
    .A2(_10904_),
    .B(_10939_),
    .Y(_03785_));
 NOR2x1_ASAP7_75t_R _30503_ (.A(_01204_),
    .B(_10904_),
    .Y(_10940_));
 AO21x1_ASAP7_75t_R _30504_ (.A1(_08563_),
    .A2(_10904_),
    .B(_10940_),
    .Y(_03786_));
 NOR2x1_ASAP7_75t_R _30505_ (.A(_01238_),
    .B(_10904_),
    .Y(_10941_));
 AO21x1_ASAP7_75t_R _30506_ (.A1(net250),
    .A2(_10904_),
    .B(_10941_),
    .Y(_03787_));
 NOR2x1_ASAP7_75t_R _30507_ (.A(_01270_),
    .B(_10904_),
    .Y(_10942_));
 AO21x1_ASAP7_75t_R _30508_ (.A1(net2197),
    .A2(_10904_),
    .B(_10942_),
    .Y(_03788_));
 INVx1_ASAP7_75t_R _30509_ (.A(_01304_),
    .Y(_10943_));
 NAND2x1_ASAP7_75t_R _30510_ (.A(_08648_),
    .B(_10904_),
    .Y(_10944_));
 OA21x2_ASAP7_75t_R _30511_ (.A1(_10943_),
    .A2(_10904_),
    .B(_10944_),
    .Y(_03789_));
 INVx1_ASAP7_75t_R _30512_ (.A(_00320_),
    .Y(_10945_));
 NOR2x2_ASAP7_75t_R _30513_ (.A(_10269_),
    .B(_10432_),
    .Y(_10946_));
 TAPCELL_ASAP7_75t_R PHY_295 ();
 TAPCELL_ASAP7_75t_R PHY_294 ();
 NAND2x1_ASAP7_75t_R _30516_ (.A(_07248_),
    .B(_10946_),
    .Y(_10949_));
 OA21x2_ASAP7_75t_R _30517_ (.A1(_10945_),
    .A2(_10946_),
    .B(_10949_),
    .Y(_03790_));
 NOR2x1_ASAP7_75t_R _30518_ (.A(_00274_),
    .B(net264),
    .Y(_10950_));
 AO21x1_ASAP7_75t_R _30519_ (.A1(_07384_),
    .A2(net264),
    .B(_10950_),
    .Y(_03791_));
 NOR2x1_ASAP7_75t_R _30520_ (.A(_00382_),
    .B(net264),
    .Y(_10951_));
 AO21x1_ASAP7_75t_R _30521_ (.A1(_07472_),
    .A2(net264),
    .B(_10951_),
    .Y(_03792_));
 NOR2x1_ASAP7_75t_R _30522_ (.A(_00413_),
    .B(_10946_),
    .Y(_10952_));
 AO21x1_ASAP7_75t_R _30523_ (.A1(_07552_),
    .A2(_10946_),
    .B(_10952_),
    .Y(_03793_));
 NOR2x1_ASAP7_75t_R _30524_ (.A(_00443_),
    .B(net264),
    .Y(_10953_));
 AO21x1_ASAP7_75t_R _30525_ (.A1(_07608_),
    .A2(net264),
    .B(_10953_),
    .Y(_03794_));
 NOR2x1_ASAP7_75t_R _30526_ (.A(_00473_),
    .B(net263),
    .Y(_10954_));
 AO21x1_ASAP7_75t_R _30527_ (.A1(_07663_),
    .A2(net263),
    .B(_10954_),
    .Y(_03795_));
 NOR2x1_ASAP7_75t_R _30528_ (.A(_00503_),
    .B(net264),
    .Y(_10955_));
 AO21x1_ASAP7_75t_R _30529_ (.A1(_07709_),
    .A2(net264),
    .B(_10955_),
    .Y(_03796_));
 NOR2x1_ASAP7_75t_R _30530_ (.A(_00533_),
    .B(net264),
    .Y(_10956_));
 AO21x1_ASAP7_75t_R _30531_ (.A1(net252),
    .A2(net264),
    .B(_10956_),
    .Y(_03797_));
 TAPCELL_ASAP7_75t_R PHY_293 ();
 NOR2x1_ASAP7_75t_R _30533_ (.A(_00563_),
    .B(net263),
    .Y(_10958_));
 AO21x1_ASAP7_75t_R _30534_ (.A1(net257),
    .A2(net263),
    .B(_10958_),
    .Y(_03798_));
 TAPCELL_ASAP7_75t_R PHY_292 ();
 NOR2x1_ASAP7_75t_R _30536_ (.A(_00593_),
    .B(net264),
    .Y(_10960_));
 AO21x1_ASAP7_75t_R _30537_ (.A1(net256),
    .A2(net264),
    .B(_10960_),
    .Y(_03799_));
 NOR2x1_ASAP7_75t_R _30538_ (.A(_00623_),
    .B(net263),
    .Y(_10961_));
 AO21x1_ASAP7_75t_R _30539_ (.A1(_07903_),
    .A2(net263),
    .B(_10961_),
    .Y(_03800_));
 NOR2x1_ASAP7_75t_R _30540_ (.A(_00653_),
    .B(net264),
    .Y(_10962_));
 AO21x1_ASAP7_75t_R _30541_ (.A1(_07948_),
    .A2(net264),
    .B(_10962_),
    .Y(_03801_));
 NOR2x1_ASAP7_75t_R _30542_ (.A(_00352_),
    .B(net263),
    .Y(_10963_));
 AO21x1_ASAP7_75t_R _30543_ (.A1(_07985_),
    .A2(net263),
    .B(_10963_),
    .Y(_03802_));
 NOR2x1_ASAP7_75t_R _30544_ (.A(_00715_),
    .B(net263),
    .Y(_10964_));
 AO21x1_ASAP7_75t_R _30545_ (.A1(net251),
    .A2(net263),
    .B(_10964_),
    .Y(_03803_));
 NOR2x1_ASAP7_75t_R _30546_ (.A(_00747_),
    .B(net263),
    .Y(_10965_));
 AO21x1_ASAP7_75t_R _30547_ (.A1(_08068_),
    .A2(net263),
    .B(_10965_),
    .Y(_03804_));
 NOR2x1_ASAP7_75t_R _30548_ (.A(_00780_),
    .B(_10946_),
    .Y(_10966_));
 AO21x1_ASAP7_75t_R _30549_ (.A1(_08110_),
    .A2(_10946_),
    .B(_10966_),
    .Y(_03805_));
 NOR2x1_ASAP7_75t_R _30550_ (.A(_00813_),
    .B(net263),
    .Y(_10967_));
 AO21x1_ASAP7_75t_R _30551_ (.A1(_08151_),
    .A2(net263),
    .B(_10967_),
    .Y(_03806_));
 NOR2x1_ASAP7_75t_R _30552_ (.A(_00846_),
    .B(net263),
    .Y(_10968_));
 AO21x1_ASAP7_75t_R _30553_ (.A1(_08190_),
    .A2(net263),
    .B(_10968_),
    .Y(_03807_));
 TAPCELL_ASAP7_75t_R PHY_291 ();
 NOR2x1_ASAP7_75t_R _30555_ (.A(_00878_),
    .B(net264),
    .Y(_10970_));
 AO21x1_ASAP7_75t_R _30556_ (.A1(_08225_),
    .A2(net264),
    .B(_10970_),
    .Y(_03808_));
 TAPCELL_ASAP7_75t_R PHY_290 ();
 NOR2x1_ASAP7_75t_R _30558_ (.A(_00911_),
    .B(net263),
    .Y(_10972_));
 AO21x1_ASAP7_75t_R _30559_ (.A1(_08263_),
    .A2(net263),
    .B(_10972_),
    .Y(_03809_));
 NOR2x1_ASAP7_75t_R _30560_ (.A(_00943_),
    .B(_10946_),
    .Y(_10973_));
 AO21x1_ASAP7_75t_R _30561_ (.A1(_08294_),
    .A2(_10946_),
    .B(_10973_),
    .Y(_03810_));
 NOR2x1_ASAP7_75t_R _30562_ (.A(_00976_),
    .B(net263),
    .Y(_10974_));
 AO21x1_ASAP7_75t_R _30563_ (.A1(_08328_),
    .A2(net263),
    .B(_10974_),
    .Y(_03811_));
 NOR2x1_ASAP7_75t_R _30564_ (.A(_01008_),
    .B(_10946_),
    .Y(_10975_));
 AO21x1_ASAP7_75t_R _30565_ (.A1(_08360_),
    .A2(_10946_),
    .B(_10975_),
    .Y(_03812_));
 NOR2x1_ASAP7_75t_R _30566_ (.A(_01042_),
    .B(net263),
    .Y(_10976_));
 AO21x1_ASAP7_75t_R _30567_ (.A1(_08406_),
    .A2(net263),
    .B(_10976_),
    .Y(_03813_));
 NOR2x1_ASAP7_75t_R _30568_ (.A(_01074_),
    .B(_10946_),
    .Y(_10977_));
 AO21x1_ASAP7_75t_R _30569_ (.A1(_08450_),
    .A2(_10946_),
    .B(_10977_),
    .Y(_03814_));
 NOR2x1_ASAP7_75t_R _30570_ (.A(_01107_),
    .B(net263),
    .Y(_10978_));
 AO21x1_ASAP7_75t_R _30571_ (.A1(_08481_),
    .A2(net263),
    .B(_10978_),
    .Y(_03815_));
 NOR2x1_ASAP7_75t_R _30572_ (.A(_01139_),
    .B(net263),
    .Y(_10979_));
 AO21x1_ASAP7_75t_R _30573_ (.A1(_08509_),
    .A2(net263),
    .B(_10979_),
    .Y(_03816_));
 NOR2x1_ASAP7_75t_R _30574_ (.A(_01173_),
    .B(net263),
    .Y(_10980_));
 AO21x1_ASAP7_75t_R _30575_ (.A1(_08537_),
    .A2(net263),
    .B(_10980_),
    .Y(_03817_));
 NOR2x1_ASAP7_75t_R _30576_ (.A(_01205_),
    .B(net264),
    .Y(_10981_));
 AO21x1_ASAP7_75t_R _30577_ (.A1(_08563_),
    .A2(net264),
    .B(_10981_),
    .Y(_03818_));
 NOR2x1_ASAP7_75t_R _30578_ (.A(_01239_),
    .B(net263),
    .Y(_10982_));
 AO21x1_ASAP7_75t_R _30579_ (.A1(net250),
    .A2(net263),
    .B(_10982_),
    .Y(_03819_));
 NOR2x1_ASAP7_75t_R _30580_ (.A(_01271_),
    .B(net264),
    .Y(_10983_));
 AO21x1_ASAP7_75t_R _30581_ (.A1(net2329),
    .A2(net264),
    .B(_10983_),
    .Y(_03820_));
 OR3x1_ASAP7_75t_R _30582_ (.A(_08648_),
    .B(_10269_),
    .C(_10432_),
    .Y(_10984_));
 OAI21x1_ASAP7_75t_R _30583_ (.A1(_01305_),
    .A2(net264),
    .B(_10984_),
    .Y(_03821_));
 AND2x6_ASAP7_75t_R _30584_ (.A(_10213_),
    .B(_10473_),
    .Y(_10985_));
 TAPCELL_ASAP7_75t_R PHY_289 ();
 TAPCELL_ASAP7_75t_R PHY_288 ();
 TAPCELL_ASAP7_75t_R PHY_287 ();
 NAND2x1_ASAP7_75t_R _30588_ (.A(_07248_),
    .B(_10985_),
    .Y(_10989_));
 OA21x2_ASAP7_75t_R _30589_ (.A1(_13856_),
    .A2(_10985_),
    .B(_10989_),
    .Y(_03822_));
 NOR2x1_ASAP7_75t_R _30590_ (.A(_00275_),
    .B(_10985_),
    .Y(_10990_));
 AO21x1_ASAP7_75t_R _30591_ (.A1(_07384_),
    .A2(_10985_),
    .B(_10990_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _30592_ (.A(_00383_),
    .B(_10985_),
    .Y(_10991_));
 AO21x1_ASAP7_75t_R _30593_ (.A1(_07472_),
    .A2(_10985_),
    .B(_10991_),
    .Y(_03824_));
 NOR2x1_ASAP7_75t_R _30594_ (.A(_00414_),
    .B(_10985_),
    .Y(_10992_));
 AO21x1_ASAP7_75t_R _30595_ (.A1(_07552_),
    .A2(_10985_),
    .B(_10992_),
    .Y(_03825_));
 NOR2x1_ASAP7_75t_R _30596_ (.A(_00444_),
    .B(_10985_),
    .Y(_10993_));
 AO21x1_ASAP7_75t_R _30597_ (.A1(_07608_),
    .A2(_10985_),
    .B(_10993_),
    .Y(_03826_));
 NOR2x1_ASAP7_75t_R _30598_ (.A(_00474_),
    .B(_10985_),
    .Y(_10994_));
 AO21x1_ASAP7_75t_R _30599_ (.A1(_07663_),
    .A2(_10985_),
    .B(_10994_),
    .Y(_03827_));
 NOR2x1_ASAP7_75t_R _30600_ (.A(_00504_),
    .B(_10985_),
    .Y(_10995_));
 AO21x1_ASAP7_75t_R _30601_ (.A1(_07709_),
    .A2(_10985_),
    .B(_10995_),
    .Y(_03828_));
 TAPCELL_ASAP7_75t_R PHY_286 ();
 NOR2x1_ASAP7_75t_R _30603_ (.A(_00534_),
    .B(_10985_),
    .Y(_10997_));
 AO21x1_ASAP7_75t_R _30604_ (.A1(_07760_),
    .A2(_10985_),
    .B(_10997_),
    .Y(_03829_));
 NOR2x1_ASAP7_75t_R _30605_ (.A(_00564_),
    .B(_10985_),
    .Y(_10998_));
 AO21x1_ASAP7_75t_R _30606_ (.A1(net257),
    .A2(_10985_),
    .B(_10998_),
    .Y(_03830_));
 TAPCELL_ASAP7_75t_R PHY_285 ();
 NOR2x1_ASAP7_75t_R _30608_ (.A(_00594_),
    .B(_10985_),
    .Y(_11000_));
 AO21x1_ASAP7_75t_R _30609_ (.A1(net256),
    .A2(_10985_),
    .B(_11000_),
    .Y(_03831_));
 NOR2x1_ASAP7_75t_R _30610_ (.A(_00624_),
    .B(_10985_),
    .Y(_11001_));
 AO21x1_ASAP7_75t_R _30611_ (.A1(_07903_),
    .A2(_10985_),
    .B(_11001_),
    .Y(_03832_));
 NOR2x1_ASAP7_75t_R _30612_ (.A(_00654_),
    .B(_10985_),
    .Y(_11002_));
 AO21x1_ASAP7_75t_R _30613_ (.A1(_07948_),
    .A2(_10985_),
    .B(_11002_),
    .Y(_03833_));
 NOR2x1_ASAP7_75t_R _30614_ (.A(_00353_),
    .B(_10985_),
    .Y(_11003_));
 AO21x1_ASAP7_75t_R _30615_ (.A1(_07985_),
    .A2(_10985_),
    .B(_11003_),
    .Y(_03834_));
 NOR2x1_ASAP7_75t_R _30616_ (.A(_00716_),
    .B(_10985_),
    .Y(_11004_));
 AO21x1_ASAP7_75t_R _30617_ (.A1(_08026_),
    .A2(_10985_),
    .B(_11004_),
    .Y(_03835_));
 NOR2x1_ASAP7_75t_R _30618_ (.A(_00748_),
    .B(_10985_),
    .Y(_11005_));
 AO21x1_ASAP7_75t_R _30619_ (.A1(_08068_),
    .A2(_10985_),
    .B(_11005_),
    .Y(_03836_));
 NOR2x1_ASAP7_75t_R _30620_ (.A(_00781_),
    .B(_10985_),
    .Y(_11006_));
 AO21x1_ASAP7_75t_R _30621_ (.A1(_08110_),
    .A2(_10985_),
    .B(_11006_),
    .Y(_03837_));
 NOR2x1_ASAP7_75t_R _30622_ (.A(_00814_),
    .B(_10985_),
    .Y(_11007_));
 AO21x1_ASAP7_75t_R _30623_ (.A1(_08151_),
    .A2(_10985_),
    .B(_11007_),
    .Y(_03838_));
 TAPCELL_ASAP7_75t_R PHY_284 ();
 NOR2x1_ASAP7_75t_R _30625_ (.A(_00847_),
    .B(_10985_),
    .Y(_11009_));
 AO21x1_ASAP7_75t_R _30626_ (.A1(_08190_),
    .A2(_10985_),
    .B(_11009_),
    .Y(_03839_));
 NOR2x1_ASAP7_75t_R _30627_ (.A(_00879_),
    .B(_10985_),
    .Y(_11010_));
 AO21x1_ASAP7_75t_R _30628_ (.A1(_08225_),
    .A2(_10985_),
    .B(_11010_),
    .Y(_03840_));
 TAPCELL_ASAP7_75t_R PHY_283 ();
 NOR2x1_ASAP7_75t_R _30630_ (.A(_00912_),
    .B(_10985_),
    .Y(_11012_));
 AO21x1_ASAP7_75t_R _30631_ (.A1(_08263_),
    .A2(_10985_),
    .B(_11012_),
    .Y(_03841_));
 NOR2x1_ASAP7_75t_R _30632_ (.A(_00944_),
    .B(_10985_),
    .Y(_11013_));
 AO21x1_ASAP7_75t_R _30633_ (.A1(_08294_),
    .A2(_10985_),
    .B(_11013_),
    .Y(_03842_));
 NOR2x1_ASAP7_75t_R _30634_ (.A(_00977_),
    .B(_10985_),
    .Y(_11014_));
 AO21x1_ASAP7_75t_R _30635_ (.A1(_08328_),
    .A2(_10985_),
    .B(_11014_),
    .Y(_03843_));
 NOR2x1_ASAP7_75t_R _30636_ (.A(_01009_),
    .B(_10985_),
    .Y(_11015_));
 AO21x1_ASAP7_75t_R _30637_ (.A1(_08360_),
    .A2(_10985_),
    .B(_11015_),
    .Y(_03844_));
 NOR2x1_ASAP7_75t_R _30638_ (.A(_01043_),
    .B(_10985_),
    .Y(_11016_));
 AO21x1_ASAP7_75t_R _30639_ (.A1(_08406_),
    .A2(_10985_),
    .B(_11016_),
    .Y(_03845_));
 NOR2x1_ASAP7_75t_R _30640_ (.A(_01075_),
    .B(_10985_),
    .Y(_11017_));
 AO21x1_ASAP7_75t_R _30641_ (.A1(_08450_),
    .A2(_10985_),
    .B(_11017_),
    .Y(_03846_));
 NOR2x1_ASAP7_75t_R _30642_ (.A(_01108_),
    .B(_10985_),
    .Y(_11018_));
 AO21x1_ASAP7_75t_R _30643_ (.A1(_08481_),
    .A2(_10985_),
    .B(_11018_),
    .Y(_03847_));
 NOR2x1_ASAP7_75t_R _30644_ (.A(_01140_),
    .B(_10985_),
    .Y(_11019_));
 AO21x1_ASAP7_75t_R _30645_ (.A1(_08509_),
    .A2(_10985_),
    .B(_11019_),
    .Y(_03848_));
 NOR2x1_ASAP7_75t_R _30646_ (.A(_01174_),
    .B(_10985_),
    .Y(_11020_));
 AO21x1_ASAP7_75t_R _30647_ (.A1(_08537_),
    .A2(_10985_),
    .B(_11020_),
    .Y(_03849_));
 NOR2x1_ASAP7_75t_R _30648_ (.A(_01206_),
    .B(_10985_),
    .Y(_11021_));
 AO21x1_ASAP7_75t_R _30649_ (.A1(_08563_),
    .A2(_10985_),
    .B(_11021_),
    .Y(_03850_));
 NOR2x1_ASAP7_75t_R _30650_ (.A(_01240_),
    .B(_10985_),
    .Y(_11022_));
 AO21x1_ASAP7_75t_R _30651_ (.A1(net250),
    .A2(_10985_),
    .B(_11022_),
    .Y(_03851_));
 NOR2x1_ASAP7_75t_R _30652_ (.A(_01272_),
    .B(_10985_),
    .Y(_11023_));
 AO21x1_ASAP7_75t_R _30653_ (.A1(net2197),
    .A2(_10985_),
    .B(_11023_),
    .Y(_03852_));
 NAND2x1_ASAP7_75t_R _30654_ (.A(_08648_),
    .B(_10985_),
    .Y(_11024_));
 OA21x2_ASAP7_75t_R _30655_ (.A1(_05444_),
    .A2(_10985_),
    .B(_11024_),
    .Y(_03853_));
 OR2x6_ASAP7_75t_R _30656_ (.A(_10269_),
    .B(_10514_),
    .Y(_11025_));
 TAPCELL_ASAP7_75t_R PHY_282 ();
 NOR2x1_ASAP7_75t_R _30658_ (.A(_07248_),
    .B(_11025_),
    .Y(_11027_));
 AO21x1_ASAP7_75t_R _30659_ (.A1(_13864_),
    .A2(_11025_),
    .B(_11027_),
    .Y(_03854_));
 NOR2x2_ASAP7_75t_R _30660_ (.A(_10269_),
    .B(_10514_),
    .Y(_11028_));
 TAPCELL_ASAP7_75t_R PHY_281 ();
 AND2x2_ASAP7_75t_R _30662_ (.A(_13426_),
    .B(_11025_),
    .Y(_11030_));
 AO21x1_ASAP7_75t_R _30663_ (.A1(_07384_),
    .A2(_11028_),
    .B(_11030_),
    .Y(_03855_));
 AND2x2_ASAP7_75t_R _30664_ (.A(_14135_),
    .B(_11025_),
    .Y(_11031_));
 AO21x1_ASAP7_75t_R _30665_ (.A1(_07472_),
    .A2(_11028_),
    .B(_11031_),
    .Y(_03856_));
 AND2x2_ASAP7_75t_R _30666_ (.A(_14960_),
    .B(_11025_),
    .Y(_11032_));
 AO21x1_ASAP7_75t_R _30667_ (.A1(_07552_),
    .A2(_11028_),
    .B(_11032_),
    .Y(_03857_));
 AND2x2_ASAP7_75t_R _30668_ (.A(_14286_),
    .B(_11025_),
    .Y(_11033_));
 AO21x1_ASAP7_75t_R _30669_ (.A1(_07608_),
    .A2(_11028_),
    .B(_11033_),
    .Y(_03858_));
 AND2x2_ASAP7_75t_R _30670_ (.A(_14319_),
    .B(_11025_),
    .Y(_11034_));
 AO21x1_ASAP7_75t_R _30671_ (.A1(_07663_),
    .A2(_11028_),
    .B(_11034_),
    .Y(_03859_));
 AND2x2_ASAP7_75t_R _30672_ (.A(_15135_),
    .B(_11025_),
    .Y(_11035_));
 AO21x1_ASAP7_75t_R _30673_ (.A1(_07709_),
    .A2(_11028_),
    .B(_11035_),
    .Y(_03860_));
 TAPCELL_ASAP7_75t_R PHY_280 ();
 AND2x2_ASAP7_75t_R _30675_ (.A(_14471_),
    .B(_11025_),
    .Y(_11037_));
 AO21x1_ASAP7_75t_R _30676_ (.A1(net252),
    .A2(_11028_),
    .B(_11037_),
    .Y(_03861_));
 AND2x2_ASAP7_75t_R _30677_ (.A(_14517_),
    .B(_11025_),
    .Y(_11038_));
 AO21x1_ASAP7_75t_R _30678_ (.A1(net257),
    .A2(_11028_),
    .B(_11038_),
    .Y(_03862_));
 AND2x2_ASAP7_75t_R _30679_ (.A(_15323_),
    .B(_11025_),
    .Y(_11039_));
 AO21x1_ASAP7_75t_R _30680_ (.A1(net256),
    .A2(_11028_),
    .B(_11039_),
    .Y(_03863_));
 AND2x2_ASAP7_75t_R _30681_ (.A(_14641_),
    .B(_11025_),
    .Y(_11040_));
 AO21x1_ASAP7_75t_R _30682_ (.A1(_07903_),
    .A2(_11028_),
    .B(_11040_),
    .Y(_03864_));
 TAPCELL_ASAP7_75t_R PHY_279 ();
 AND2x2_ASAP7_75t_R _30684_ (.A(_14768_),
    .B(_11025_),
    .Y(_11042_));
 AO21x1_ASAP7_75t_R _30685_ (.A1(_07948_),
    .A2(_11028_),
    .B(_11042_),
    .Y(_03865_));
 AND2x2_ASAP7_75t_R _30686_ (.A(_14078_),
    .B(_11025_),
    .Y(_11043_));
 AO21x1_ASAP7_75t_R _30687_ (.A1(_07985_),
    .A2(_11028_),
    .B(_11043_),
    .Y(_03866_));
 AND2x2_ASAP7_75t_R _30688_ (.A(_15581_),
    .B(_11025_),
    .Y(_11044_));
 AO21x1_ASAP7_75t_R _30689_ (.A1(net251),
    .A2(_11028_),
    .B(_11044_),
    .Y(_03867_));
 AND2x2_ASAP7_75t_R _30690_ (.A(_15714_),
    .B(_11025_),
    .Y(_11045_));
 AO21x1_ASAP7_75t_R _30691_ (.A1(_08068_),
    .A2(_11028_),
    .B(_11045_),
    .Y(_03868_));
 AND2x2_ASAP7_75t_R _30692_ (.A(_15823_),
    .B(_11025_),
    .Y(_11046_));
 AO21x1_ASAP7_75t_R _30693_ (.A1(_08110_),
    .A2(_11028_),
    .B(_11046_),
    .Y(_03869_));
 AND2x2_ASAP7_75t_R _30694_ (.A(_15943_),
    .B(_11025_),
    .Y(_11047_));
 AO21x1_ASAP7_75t_R _30695_ (.A1(_08151_),
    .A2(_11028_),
    .B(_11047_),
    .Y(_03870_));
 TAPCELL_ASAP7_75t_R PHY_278 ();
 AND2x2_ASAP7_75t_R _30697_ (.A(_16077_),
    .B(_11025_),
    .Y(_11049_));
 AO21x1_ASAP7_75t_R _30698_ (.A1(_08190_),
    .A2(_11028_),
    .B(_11049_),
    .Y(_03871_));
 AND2x2_ASAP7_75t_R _30699_ (.A(_16185_),
    .B(_11025_),
    .Y(_11050_));
 AO21x1_ASAP7_75t_R _30700_ (.A1(_08225_),
    .A2(_11028_),
    .B(_11050_),
    .Y(_03872_));
 AND2x2_ASAP7_75t_R _30701_ (.A(_16287_),
    .B(_11025_),
    .Y(_11051_));
 AO21x1_ASAP7_75t_R _30702_ (.A1(_08263_),
    .A2(_11028_),
    .B(_11051_),
    .Y(_03873_));
 AND2x2_ASAP7_75t_R _30703_ (.A(_16424_),
    .B(_11025_),
    .Y(_11052_));
 AO21x1_ASAP7_75t_R _30704_ (.A1(_08294_),
    .A2(_11028_),
    .B(_11052_),
    .Y(_03874_));
 TAPCELL_ASAP7_75t_R PHY_277 ();
 AND2x2_ASAP7_75t_R _30706_ (.A(_16559_),
    .B(_11025_),
    .Y(_11054_));
 AO21x1_ASAP7_75t_R _30707_ (.A1(_08328_),
    .A2(_11028_),
    .B(_11054_),
    .Y(_03875_));
 AND2x2_ASAP7_75t_R _30708_ (.A(_16663_),
    .B(_11025_),
    .Y(_11055_));
 AO21x1_ASAP7_75t_R _30709_ (.A1(_08360_),
    .A2(_11028_),
    .B(_11055_),
    .Y(_03876_));
 AND2x2_ASAP7_75t_R _30710_ (.A(_04552_),
    .B(_11025_),
    .Y(_11056_));
 AO21x1_ASAP7_75t_R _30711_ (.A1(_08406_),
    .A2(_11028_),
    .B(_11056_),
    .Y(_03877_));
 AND2x2_ASAP7_75t_R _30712_ (.A(_04681_),
    .B(_11025_),
    .Y(_11057_));
 AO21x1_ASAP7_75t_R _30713_ (.A1(_08450_),
    .A2(_11028_),
    .B(_11057_),
    .Y(_03878_));
 AND2x2_ASAP7_75t_R _30714_ (.A(_04799_),
    .B(_11025_),
    .Y(_11058_));
 AO21x1_ASAP7_75t_R _30715_ (.A1(_08481_),
    .A2(_11028_),
    .B(_11058_),
    .Y(_03879_));
 AND2x2_ASAP7_75t_R _30716_ (.A(_04907_),
    .B(_11025_),
    .Y(_11059_));
 AO21x1_ASAP7_75t_R _30717_ (.A1(_08509_),
    .A2(_11028_),
    .B(_11059_),
    .Y(_03880_));
 AND2x2_ASAP7_75t_R _30718_ (.A(_05003_),
    .B(_11025_),
    .Y(_11060_));
 AO21x1_ASAP7_75t_R _30719_ (.A1(_08537_),
    .A2(_11028_),
    .B(_11060_),
    .Y(_03881_));
 AND2x2_ASAP7_75t_R _30720_ (.A(_05112_),
    .B(_11025_),
    .Y(_11061_));
 AO21x1_ASAP7_75t_R _30721_ (.A1(_08563_),
    .A2(_11028_),
    .B(_11061_),
    .Y(_03882_));
 AND2x2_ASAP7_75t_R _30722_ (.A(_05220_),
    .B(_11025_),
    .Y(_11062_));
 AO21x1_ASAP7_75t_R _30723_ (.A1(net250),
    .A2(_11028_),
    .B(_11062_),
    .Y(_03883_));
 AND2x2_ASAP7_75t_R _30724_ (.A(_05346_),
    .B(_11025_),
    .Y(_11063_));
 AO21x1_ASAP7_75t_R _30725_ (.A1(net2198),
    .A2(_11028_),
    .B(_11063_),
    .Y(_03884_));
 NOR2x1_ASAP7_75t_R _30726_ (.A(_08648_),
    .B(_11025_),
    .Y(_11064_));
 AO21x1_ASAP7_75t_R _30727_ (.A1(_05441_),
    .A2(_11025_),
    .B(_11064_),
    .Y(_03885_));
 OR4x1_ASAP7_75t_R _30728_ (.A(_01872_),
    .B(_05547_),
    .C(_05769_),
    .D(_08653_),
    .Y(_11065_));
 NAND2x1_ASAP7_75t_R _30729_ (.A(_01519_),
    .B(_11065_),
    .Y(_11066_));
 OA21x2_ASAP7_75t_R _30730_ (.A1(_06627_),
    .A2(_11065_),
    .B(_11066_),
    .Y(_03886_));
 AND2x2_ASAP7_75t_R _30731_ (.A(_13999_),
    .B(_14713_),
    .Y(_11067_));
 AO21x1_ASAP7_75t_R _30732_ (.A1(_02289_),
    .A2(_18326_),
    .B(_11067_),
    .Y(_11068_));
 AO22x2_ASAP7_75t_R _30733_ (.A1(_18326_),
    .A2(_07032_),
    .B1(_11068_),
    .B2(_02286_),
    .Y(_11069_));
 TAPCELL_ASAP7_75t_R PHY_276 ();
 AND4x1_ASAP7_75t_R _30735_ (.A(_14297_),
    .B(_05643_),
    .C(net310),
    .D(_05596_),
    .Y(_11071_));
 AND3x1_ASAP7_75t_R _30736_ (.A(_05586_),
    .B(_11071_),
    .C(_06945_),
    .Y(_11072_));
 OR5x1_ASAP7_75t_R _30737_ (.A(_13595_),
    .B(_01740_),
    .C(_01741_),
    .D(_13497_),
    .E(_05563_),
    .Y(_11073_));
 AO21x2_ASAP7_75t_R _30738_ (.A1(_13520_),
    .A2(_14542_),
    .B(_11073_),
    .Y(_11074_));
 NOR2x1_ASAP7_75t_R _30739_ (.A(_14709_),
    .B(_11074_),
    .Y(_11075_));
 NAND3x2_ASAP7_75t_R _30740_ (.B(_13894_),
    .C(_06954_),
    .Y(_11076_),
    .A(_13523_));
 AO32x2_ASAP7_75t_R _30741_ (.A1(_05613_),
    .A2(_11075_),
    .A3(_11076_),
    .B1(_11071_),
    .B2(_05656_),
    .Y(_11077_));
 AND2x2_ASAP7_75t_R _30742_ (.A(_14296_),
    .B(_06973_),
    .Y(_11078_));
 AND3x1_ASAP7_75t_R _30743_ (.A(_05663_),
    .B(_05679_),
    .C(_11078_),
    .Y(_11079_));
 AND3x1_ASAP7_75t_R _30744_ (.A(_05601_),
    .B(_06942_),
    .C(_06943_),
    .Y(_11080_));
 AOI211x1_ASAP7_75t_R _30745_ (.A1(_05594_),
    .A2(_14424_),
    .B(_05598_),
    .C(_11074_),
    .Y(_11081_));
 AND2x2_ASAP7_75t_R _30746_ (.A(_14296_),
    .B(_11081_),
    .Y(_11082_));
 OA211x2_ASAP7_75t_R _30747_ (.A1(_14359_),
    .A2(_05693_),
    .B(_06955_),
    .C(_11082_),
    .Y(_11083_));
 OR4x1_ASAP7_75t_R _30748_ (.A(_11077_),
    .B(_11079_),
    .C(_11080_),
    .D(_11083_),
    .Y(_11084_));
 NOR2x1_ASAP7_75t_R _30749_ (.A(_05598_),
    .B(_11074_),
    .Y(_11085_));
 AND3x4_ASAP7_75t_R _30750_ (.A(_05627_),
    .B(_05630_),
    .C(_11085_),
    .Y(_11086_));
 AND4x2_ASAP7_75t_R _30751_ (.A(_14710_),
    .B(_05568_),
    .C(_05584_),
    .D(_05586_),
    .Y(_11087_));
 AND3x1_ASAP7_75t_R _30752_ (.A(_05724_),
    .B(_06968_),
    .C(_11087_),
    .Y(_11088_));
 AO21x1_ASAP7_75t_R _30753_ (.A1(_06968_),
    .A2(_11086_),
    .B(_11088_),
    .Y(_11089_));
 OR2x2_ASAP7_75t_R _30754_ (.A(_05667_),
    .B(_06962_),
    .Y(_11090_));
 AO33x2_ASAP7_75t_R _30755_ (.A1(_14358_),
    .A2(_11081_),
    .A3(_11090_),
    .B1(_06971_),
    .B2(_06972_),
    .B3(_11085_),
    .Y(_11091_));
 OR2x2_ASAP7_75t_R _30756_ (.A(_05693_),
    .B(_06959_),
    .Y(_11092_));
 OA21x2_ASAP7_75t_R _30757_ (.A1(_14297_),
    .A2(_11076_),
    .B(_14359_),
    .Y(_11093_));
 AO33x2_ASAP7_75t_R _30758_ (.A1(_11081_),
    .A2(_11092_),
    .A3(_06960_),
    .B1(_11093_),
    .B2(_05568_),
    .B3(_11075_),
    .Y(_11094_));
 OR4x1_ASAP7_75t_R _30759_ (.A(_11084_),
    .B(_11089_),
    .C(_11091_),
    .D(_11094_),
    .Y(_11095_));
 OA21x2_ASAP7_75t_R _30760_ (.A1(_11072_),
    .A2(_11095_),
    .B(_09443_),
    .Y(_11096_));
 TAPCELL_ASAP7_75t_R PHY_275 ();
 AND3x4_ASAP7_75t_R _30762_ (.A(_05568_),
    .B(_05616_),
    .C(_05627_),
    .Y(_11098_));
 NOR2x2_ASAP7_75t_R _30763_ (.A(_07359_),
    .B(_11098_),
    .Y(_11099_));
 INVx2_ASAP7_75t_R _30764_ (.A(_11099_),
    .Y(_11100_));
 AND3x4_ASAP7_75t_R _30765_ (.A(_05693_),
    .B(_11096_),
    .C(_11100_),
    .Y(_11101_));
 TAPCELL_ASAP7_75t_R PHY_274 ();
 INVx1_ASAP7_75t_R _30767_ (.A(_00661_),
    .Y(_11103_));
 AND3x1_ASAP7_75t_R _30768_ (.A(_05693_),
    .B(_09443_),
    .C(_11098_),
    .Y(_11104_));
 AND3x2_ASAP7_75t_R _30769_ (.A(_05693_),
    .B(_07359_),
    .C(_09443_),
    .Y(_11105_));
 INVx2_ASAP7_75t_R _30770_ (.A(_11105_),
    .Y(_11106_));
 OA21x2_ASAP7_75t_R _30771_ (.A1(_11103_),
    .A2(_11104_),
    .B(_11106_),
    .Y(_11107_));
 TAPCELL_ASAP7_75t_R PHY_273 ();
 TAPCELL_ASAP7_75t_R PHY_272 ();
 AO21x1_ASAP7_75t_R _30774_ (.A1(net3517),
    .A2(_11101_),
    .B(_11107_),
    .Y(_11110_));
 NOR2x2_ASAP7_75t_R _30775_ (.A(_05698_),
    .B(_11098_),
    .Y(_11111_));
 AND3x1_ASAP7_75t_R _30776_ (.A(net302),
    .B(_05602_),
    .C(_07790_),
    .Y(_11112_));
 AND2x2_ASAP7_75t_R _30777_ (.A(_11092_),
    .B(_07450_),
    .Y(_11113_));
 AO32x1_ASAP7_75t_R _30778_ (.A1(_06968_),
    .A2(_05627_),
    .A3(_05630_),
    .B1(_06971_),
    .B2(_06972_),
    .Y(_11114_));
 AO32x1_ASAP7_75t_R _30779_ (.A1(_14358_),
    .A2(_05602_),
    .A3(_11090_),
    .B1(_11114_),
    .B2(_05601_),
    .Y(_11115_));
 OR4x1_ASAP7_75t_R _30780_ (.A(_05591_),
    .B(_11113_),
    .C(_11115_),
    .D(_11079_),
    .Y(_11116_));
 OR4x1_ASAP7_75t_R _30781_ (.A(_07438_),
    .B(_07441_),
    .C(_07443_),
    .D(_11080_),
    .Y(_11117_));
 OR3x2_ASAP7_75t_R _30782_ (.A(_11112_),
    .B(_11116_),
    .C(_11117_),
    .Y(_11118_));
 NAND2x2_ASAP7_75t_R _30783_ (.A(_09443_),
    .B(_11118_),
    .Y(_11119_));
 OR3x4_ASAP7_75t_R _30784_ (.A(_06992_),
    .B(_11111_),
    .C(_11119_),
    .Y(_11120_));
 TAPCELL_ASAP7_75t_R PHY_271 ();
 NAND3x2_ASAP7_75t_R _30786_ (.B(_09443_),
    .C(_11098_),
    .Y(_11122_),
    .A(_05693_));
 AO21x2_ASAP7_75t_R _30787_ (.A1(_00661_),
    .A2(_11122_),
    .B(_11105_),
    .Y(_11123_));
 TAPCELL_ASAP7_75t_R PHY_270 ();
 OA211x2_ASAP7_75t_R _30789_ (.A1(net3517),
    .A2(_11120_),
    .B(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .C(_11123_),
    .Y(_11125_));
 AOI21x1_ASAP7_75t_R _30790_ (.A1(_00659_),
    .A2(_11110_),
    .B(_11125_),
    .Y(_03887_));
 AND3x1_ASAP7_75t_R _30791_ (.A(_05627_),
    .B(_05630_),
    .C(_06941_),
    .Y(_11126_));
 AND3x1_ASAP7_75t_R _30792_ (.A(_05724_),
    .B(_14424_),
    .C(_05585_),
    .Y(_11127_));
 AND4x1_ASAP7_75t_R _30793_ (.A(_14710_),
    .B(_05568_),
    .C(_05584_),
    .D(_11127_),
    .Y(_11128_));
 OA21x2_ASAP7_75t_R _30794_ (.A1(_11126_),
    .A2(_11128_),
    .B(_06968_),
    .Y(_11129_));
 AND5x2_ASAP7_75t_R _30795_ (.A(_13531_),
    .B(_14424_),
    .C(_14709_),
    .D(_05570_),
    .E(_05572_),
    .Y(_11130_));
 AND3x1_ASAP7_75t_R _30796_ (.A(_13523_),
    .B(_06954_),
    .C(_09439_),
    .Y(_11131_));
 AO32x1_ASAP7_75t_R _30797_ (.A1(_14358_),
    .A2(_11090_),
    .A3(_11130_),
    .B1(_11131_),
    .B2(_05588_),
    .Y(_11132_));
 AND4x1_ASAP7_75t_R _30798_ (.A(_14297_),
    .B(_14359_),
    .C(_05570_),
    .D(_05596_),
    .Y(_11133_));
 AO33x2_ASAP7_75t_R _30799_ (.A1(_14296_),
    .A2(_07790_),
    .A3(_11130_),
    .B1(_11133_),
    .B2(_06945_),
    .B3(_05586_),
    .Y(_11134_));
 OR4x1_ASAP7_75t_R _30800_ (.A(_09438_),
    .B(_11129_),
    .C(_11132_),
    .D(_11134_),
    .Y(_11135_));
 AND2x2_ASAP7_75t_R _30801_ (.A(_06960_),
    .B(_11130_),
    .Y(_11136_));
 AO32x1_ASAP7_75t_R _30802_ (.A1(_05616_),
    .A2(_11076_),
    .A3(_06949_),
    .B1(_11133_),
    .B2(_05656_),
    .Y(_11137_));
 OA211x2_ASAP7_75t_R _30803_ (.A1(_14297_),
    .A2(_11076_),
    .B(_08426_),
    .C(_14359_),
    .Y(_11138_));
 OR3x1_ASAP7_75t_R _30804_ (.A(_06944_),
    .B(_11137_),
    .C(_11138_),
    .Y(_11139_));
 AO21x1_ASAP7_75t_R _30805_ (.A1(_11092_),
    .A2(_11136_),
    .B(_11139_),
    .Y(_11140_));
 OA21x2_ASAP7_75t_R _30806_ (.A1(_11135_),
    .A2(_11140_),
    .B(_09443_),
    .Y(_11141_));
 TAPCELL_ASAP7_75t_R PHY_269 ();
 INVx1_ASAP7_75t_R _30808_ (.A(_11141_),
    .Y(_11143_));
 OR3x4_ASAP7_75t_R _30809_ (.A(_06992_),
    .B(_11143_),
    .C(_11099_),
    .Y(_11144_));
 TAPCELL_ASAP7_75t_R PHY_268 ();
 TAPCELL_ASAP7_75t_R PHY_267 ();
 INVx1_ASAP7_75t_R _30812_ (.A(_11096_),
    .Y(_11147_));
 OR3x4_ASAP7_75t_R _30813_ (.A(_06992_),
    .B(_11147_),
    .C(_11099_),
    .Y(_11148_));
 TAPCELL_ASAP7_75t_R PHY_266 ();
 NAND2x1_ASAP7_75t_R _30815_ (.A(_02456_),
    .B(_11148_),
    .Y(_11150_));
 TAPCELL_ASAP7_75t_R PHY_265 ();
 OA211x2_ASAP7_75t_R _30817_ (.A1(net3647),
    .A2(_11144_),
    .B(_11150_),
    .C(_11123_),
    .Y(_11152_));
 AO21x1_ASAP7_75t_R _30818_ (.A1(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .A2(_11107_),
    .B(_11152_),
    .Y(_03888_));
 TAPCELL_ASAP7_75t_R PHY_264 ();
 TAPCELL_ASAP7_75t_R PHY_263 ();
 OR2x6_ASAP7_75t_R _30821_ (.A(_05657_),
    .B(_07359_),
    .Y(_11155_));
 AND3x4_ASAP7_75t_R _30822_ (.A(_05693_),
    .B(_11141_),
    .C(_11155_),
    .Y(_11156_));
 TAPCELL_ASAP7_75t_R PHY_262 ();
 TAPCELL_ASAP7_75t_R PHY_261 ();
 AOI21x1_ASAP7_75t_R _30825_ (.A1(_18336_),
    .A2(net3525),
    .B(_09471_),
    .Y(_11159_));
 AND2x2_ASAP7_75t_R _30826_ (.A(_11159_),
    .B(_11101_),
    .Y(_11160_));
 INVx1_ASAP7_75t_R _30827_ (.A(_11160_),
    .Y(_11161_));
 OA211x2_ASAP7_75t_R _30828_ (.A1(_02458_),
    .A2(_11156_),
    .B(_11161_),
    .C(_11123_),
    .Y(_11162_));
 AOI21x1_ASAP7_75t_R _30829_ (.A1(_01517_),
    .A2(_11107_),
    .B(_11162_),
    .Y(_03889_));
 TAPCELL_ASAP7_75t_R PHY_260 ();
 TAPCELL_ASAP7_75t_R PHY_259 ();
 NOR2x1_ASAP7_75t_R _30832_ (.A(_01516_),
    .B(_02457_),
    .Y(_11165_));
 NOR2x1_ASAP7_75t_R _30833_ (.A(net3544),
    .B(_11148_),
    .Y(_11166_));
 AO21x1_ASAP7_75t_R _30834_ (.A1(_11144_),
    .A2(_11165_),
    .B(_11166_),
    .Y(_11167_));
 TAPCELL_ASAP7_75t_R PHY_258 ();
 AO21x1_ASAP7_75t_R _30836_ (.A1(_02457_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11169_));
 AOI22x1_ASAP7_75t_R _30837_ (.A1(_11123_),
    .A2(_11167_),
    .B1(_11169_),
    .B2(_01516_),
    .Y(_03890_));
 TAPCELL_ASAP7_75t_R PHY_257 ();
 NOR2x1_ASAP7_75t_R _30839_ (.A(_02460_),
    .B(_11156_),
    .Y(_11171_));
 NOR2x1_ASAP7_75t_R _30840_ (.A(net3378),
    .B(_11148_),
    .Y(_11172_));
 OR3x1_ASAP7_75t_R _30841_ (.A(_11107_),
    .B(_11171_),
    .C(_11172_),
    .Y(_11173_));
 OA21x2_ASAP7_75t_R _30842_ (.A1(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .A2(_11123_),
    .B(_11173_),
    .Y(_03891_));
 NOR2x1_ASAP7_75t_R _30843_ (.A(_01514_),
    .B(_02459_),
    .Y(_11174_));
 NOR2x1_ASAP7_75t_R _30844_ (.A(net3632),
    .B(_11120_),
    .Y(_11175_));
 AO21x1_ASAP7_75t_R _30845_ (.A1(_11144_),
    .A2(_11174_),
    .B(_11175_),
    .Y(_11176_));
 AO21x1_ASAP7_75t_R _30846_ (.A1(_02459_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11177_));
 AOI22x1_ASAP7_75t_R _30847_ (.A1(_11123_),
    .A2(_11176_),
    .B1(_11177_),
    .B2(_01514_),
    .Y(_03892_));
 NAND2x1_ASAP7_75t_R _30848_ (.A(_09504_),
    .B(_11156_),
    .Y(_11178_));
 OA211x2_ASAP7_75t_R _30849_ (.A1(_02462_),
    .A2(_11156_),
    .B(_11178_),
    .C(_11123_),
    .Y(_11179_));
 AOI21x1_ASAP7_75t_R _30850_ (.A1(_01513_),
    .A2(_11107_),
    .B(_11179_),
    .Y(_03893_));
 TAPCELL_ASAP7_75t_R PHY_256 ();
 NOR2x1_ASAP7_75t_R _30852_ (.A(_01512_),
    .B(_02461_),
    .Y(_11181_));
 INVx2_ASAP7_75t_R _30853_ (.A(net3615),
    .Y(_11182_));
 AND2x2_ASAP7_75t_R _30854_ (.A(_11182_),
    .B(_11101_),
    .Y(_11183_));
 AO21x1_ASAP7_75t_R _30855_ (.A1(_11120_),
    .A2(_11181_),
    .B(_11183_),
    .Y(_11184_));
 AO21x1_ASAP7_75t_R _30856_ (.A1(_02461_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11185_));
 AOI22x1_ASAP7_75t_R _30857_ (.A1(_11123_),
    .A2(_11184_),
    .B1(_11185_),
    .B2(_01512_),
    .Y(_03894_));
 NAND2x1_ASAP7_75t_R _30858_ (.A(_09518_),
    .B(_11101_),
    .Y(_11186_));
 OA211x2_ASAP7_75t_R _30859_ (.A1(_02464_),
    .A2(_11156_),
    .B(_11186_),
    .C(_11123_),
    .Y(_11187_));
 AOI21x1_ASAP7_75t_R _30860_ (.A1(_01511_),
    .A2(_11107_),
    .B(_11187_),
    .Y(_03895_));
 NOR2x1_ASAP7_75t_R _30861_ (.A(_01510_),
    .B(_02463_),
    .Y(_11188_));
 NOR2x1_ASAP7_75t_R _30862_ (.A(_09524_),
    .B(_11120_),
    .Y(_11189_));
 AO21x1_ASAP7_75t_R _30863_ (.A1(_11144_),
    .A2(_11188_),
    .B(_11189_),
    .Y(_11190_));
 AO21x1_ASAP7_75t_R _30864_ (.A1(_02463_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11191_));
 AOI22x1_ASAP7_75t_R _30865_ (.A1(_11123_),
    .A2(_11190_),
    .B1(_11191_),
    .B2(_01510_),
    .Y(_03896_));
 NAND2x1_ASAP7_75t_R _30866_ (.A(_09531_),
    .B(_11156_),
    .Y(_11192_));
 OA211x2_ASAP7_75t_R _30867_ (.A1(_02466_),
    .A2(_11156_),
    .B(_11192_),
    .C(_11123_),
    .Y(_11193_));
 AOI21x1_ASAP7_75t_R _30868_ (.A1(_01509_),
    .A2(_11107_),
    .B(_11193_),
    .Y(_03897_));
 NOR2x1_ASAP7_75t_R _30869_ (.A(_01508_),
    .B(_02465_),
    .Y(_11194_));
 NOR2x1_ASAP7_75t_R _30870_ (.A(_09538_),
    .B(_11148_),
    .Y(_11195_));
 AO21x1_ASAP7_75t_R _30871_ (.A1(_11144_),
    .A2(_11194_),
    .B(_11195_),
    .Y(_11196_));
 AO21x1_ASAP7_75t_R _30872_ (.A1(_02465_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11197_));
 AOI22x1_ASAP7_75t_R _30873_ (.A1(_11123_),
    .A2(_11196_),
    .B1(_11197_),
    .B2(_01508_),
    .Y(_03898_));
 AND3x4_ASAP7_75t_R _30874_ (.A(_05693_),
    .B(_11141_),
    .C(_11100_),
    .Y(_11198_));
 TAPCELL_ASAP7_75t_R PHY_255 ();
 NAND2x1_ASAP7_75t_R _30876_ (.A(_09548_),
    .B(_11101_),
    .Y(_11200_));
 OA211x2_ASAP7_75t_R _30877_ (.A1(_02468_),
    .A2(_11198_),
    .B(_11200_),
    .C(_11123_),
    .Y(_11201_));
 AOI21x1_ASAP7_75t_R _30878_ (.A1(_01507_),
    .A2(_11107_),
    .B(_11201_),
    .Y(_03899_));
 NOR2x1_ASAP7_75t_R _30879_ (.A(_01506_),
    .B(_02467_),
    .Y(_11202_));
 NOR2x1_ASAP7_75t_R _30880_ (.A(_09556_),
    .B(_11148_),
    .Y(_11203_));
 AO21x1_ASAP7_75t_R _30881_ (.A1(_11120_),
    .A2(_11202_),
    .B(_11203_),
    .Y(_11204_));
 AO21x1_ASAP7_75t_R _30882_ (.A1(_02467_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11205_));
 AOI22x1_ASAP7_75t_R _30883_ (.A1(_11123_),
    .A2(_11204_),
    .B1(_11205_),
    .B2(_01506_),
    .Y(_03900_));
 NAND2x1_ASAP7_75t_R _30884_ (.A(net3541),
    .B(_11156_),
    .Y(_11206_));
 OA211x2_ASAP7_75t_R _30885_ (.A1(_02470_),
    .A2(_11156_),
    .B(_11206_),
    .C(_11123_),
    .Y(_11207_));
 AOI21x1_ASAP7_75t_R _30886_ (.A1(_01505_),
    .A2(_11107_),
    .B(_11207_),
    .Y(_03901_));
 NOR2x1_ASAP7_75t_R _30887_ (.A(_01504_),
    .B(_02469_),
    .Y(_11208_));
 NOR2x1_ASAP7_75t_R _30888_ (.A(_09575_),
    .B(_11148_),
    .Y(_11209_));
 AO21x1_ASAP7_75t_R _30889_ (.A1(_11120_),
    .A2(_11208_),
    .B(_11209_),
    .Y(_11210_));
 AO21x1_ASAP7_75t_R _30890_ (.A1(_02469_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11211_));
 AOI22x1_ASAP7_75t_R _30891_ (.A1(_11123_),
    .A2(_11210_),
    .B1(_11211_),
    .B2(_01504_),
    .Y(_03902_));
 NOR2x1_ASAP7_75t_R _30892_ (.A(_02472_),
    .B(_11156_),
    .Y(_11212_));
 AND2x2_ASAP7_75t_R _30893_ (.A(net3622),
    .B(_11156_),
    .Y(_11213_));
 OR3x1_ASAP7_75t_R _30894_ (.A(_11107_),
    .B(_11212_),
    .C(_11213_),
    .Y(_11214_));
 OA21x2_ASAP7_75t_R _30895_ (.A1(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .A2(_11123_),
    .B(_11214_),
    .Y(_03903_));
 AND3x1_ASAP7_75t_R _30896_ (.A(_05693_),
    .B(_05698_),
    .C(_09443_),
    .Y(_11215_));
 INVx1_ASAP7_75t_R _30897_ (.A(_11215_),
    .Y(_11216_));
 AO21x1_ASAP7_75t_R _30898_ (.A1(_02471_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11217_));
 NAND2x1_ASAP7_75t_R _30899_ (.A(_01502_),
    .B(_11217_),
    .Y(_11218_));
 OR4x1_ASAP7_75t_R _30900_ (.A(_01502_),
    .B(_02471_),
    .C(_11107_),
    .D(_11156_),
    .Y(_11219_));
 OA211x2_ASAP7_75t_R _30901_ (.A1(net3660),
    .A2(_11216_),
    .B(_11218_),
    .C(_11219_),
    .Y(_03904_));
 OR2x2_ASAP7_75t_R _30902_ (.A(net3571),
    .B(_11144_),
    .Y(_11220_));
 OA211x2_ASAP7_75t_R _30903_ (.A1(_02474_),
    .A2(_11198_),
    .B(_11220_),
    .C(_11123_),
    .Y(_11221_));
 AOI21x1_ASAP7_75t_R _30904_ (.A1(_01501_),
    .A2(_11107_),
    .B(_11221_),
    .Y(_03905_));
 NOR2x1_ASAP7_75t_R _30905_ (.A(_01500_),
    .B(_02473_),
    .Y(_11222_));
 NOR2x1_ASAP7_75t_R _30906_ (.A(net3711),
    .B(_11148_),
    .Y(_11223_));
 AO21x1_ASAP7_75t_R _30907_ (.A1(_11144_),
    .A2(_11222_),
    .B(_11223_),
    .Y(_11224_));
 AO21x1_ASAP7_75t_R _30908_ (.A1(_02473_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11225_));
 AOI22x1_ASAP7_75t_R _30909_ (.A1(_11123_),
    .A2(_11224_),
    .B1(_11225_),
    .B2(_01500_),
    .Y(_03906_));
 OR2x2_ASAP7_75t_R _30910_ (.A(_09615_),
    .B(_11148_),
    .Y(_11226_));
 OA211x2_ASAP7_75t_R _30911_ (.A1(_02476_),
    .A2(_11198_),
    .B(_11226_),
    .C(_11123_),
    .Y(_11227_));
 AOI21x1_ASAP7_75t_R _30912_ (.A1(_01499_),
    .A2(_11107_),
    .B(_11227_),
    .Y(_03907_));
 AO21x1_ASAP7_75t_R _30913_ (.A1(_02475_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11228_));
 NAND2x1_ASAP7_75t_R _30914_ (.A(_01498_),
    .B(_11228_),
    .Y(_11229_));
 OR4x1_ASAP7_75t_R _30915_ (.A(_01498_),
    .B(_02475_),
    .C(_11107_),
    .D(_11198_),
    .Y(_11230_));
 OA211x2_ASAP7_75t_R _30916_ (.A1(_09623_),
    .A2(_11106_),
    .B(_11229_),
    .C(_11230_),
    .Y(_03908_));
 NAND2x1_ASAP7_75t_R _30917_ (.A(_09631_),
    .B(_11198_),
    .Y(_11231_));
 OA211x2_ASAP7_75t_R _30918_ (.A1(_02478_),
    .A2(_11198_),
    .B(_11231_),
    .C(_11123_),
    .Y(_11232_));
 AOI21x1_ASAP7_75t_R _30919_ (.A1(_01497_),
    .A2(_11107_),
    .B(_11232_),
    .Y(_03909_));
 NOR2x1_ASAP7_75t_R _30920_ (.A(_01496_),
    .B(_02477_),
    .Y(_11233_));
 AND2x2_ASAP7_75t_R _30921_ (.A(net3599),
    .B(_11101_),
    .Y(_11234_));
 AO21x1_ASAP7_75t_R _30922_ (.A1(_11120_),
    .A2(_11233_),
    .B(_11234_),
    .Y(_11235_));
 AO21x1_ASAP7_75t_R _30923_ (.A1(_02477_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11236_));
 AOI22x1_ASAP7_75t_R _30924_ (.A1(_11123_),
    .A2(_11235_),
    .B1(_11236_),
    .B2(_01496_),
    .Y(_03910_));
 OR2x2_ASAP7_75t_R _30925_ (.A(net3531),
    .B(_09646_),
    .Y(_11237_));
 OR2x2_ASAP7_75t_R _30926_ (.A(_02480_),
    .B(_11156_),
    .Y(_11238_));
 OA211x2_ASAP7_75t_R _30927_ (.A1(_11237_),
    .A2(_11120_),
    .B(_11238_),
    .C(_11123_),
    .Y(_11239_));
 AOI21x1_ASAP7_75t_R _30928_ (.A1(_01495_),
    .A2(_11107_),
    .B(_11239_),
    .Y(_03911_));
 NOR2x1_ASAP7_75t_R _30929_ (.A(_01494_),
    .B(_02479_),
    .Y(_11240_));
 NOR2x1_ASAP7_75t_R _30930_ (.A(net3643),
    .B(_11148_),
    .Y(_11241_));
 AO21x1_ASAP7_75t_R _30931_ (.A1(_11144_),
    .A2(_11240_),
    .B(_11241_),
    .Y(_11242_));
 AO21x1_ASAP7_75t_R _30932_ (.A1(_02479_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11243_));
 AOI22x1_ASAP7_75t_R _30933_ (.A1(_11123_),
    .A2(_11242_),
    .B1(_11243_),
    .B2(_01494_),
    .Y(_03912_));
 NAND2x1_ASAP7_75t_R _30934_ (.A(_09662_),
    .B(_11156_),
    .Y(_11244_));
 OA211x2_ASAP7_75t_R _30935_ (.A1(_02482_),
    .A2(_11156_),
    .B(_11244_),
    .C(_11123_),
    .Y(_11245_));
 AOI21x1_ASAP7_75t_R _30936_ (.A1(_01493_),
    .A2(_11107_),
    .B(_11245_),
    .Y(_03913_));
 NOR2x1_ASAP7_75t_R _30937_ (.A(_01492_),
    .B(_02481_),
    .Y(_11246_));
 NOR2x1_ASAP7_75t_R _30938_ (.A(net3594),
    .B(_11148_),
    .Y(_11247_));
 AO21x1_ASAP7_75t_R _30939_ (.A1(_11120_),
    .A2(_11246_),
    .B(_11247_),
    .Y(_11248_));
 TAPCELL_ASAP7_75t_R PHY_254 ();
 AO21x1_ASAP7_75t_R _30941_ (.A1(_02481_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11250_));
 AOI22x1_ASAP7_75t_R _30942_ (.A1(_11123_),
    .A2(_11248_),
    .B1(_11250_),
    .B2(_01492_),
    .Y(_03914_));
 NAND2x1_ASAP7_75t_R _30943_ (.A(_09676_),
    .B(_11198_),
    .Y(_11251_));
 OA211x2_ASAP7_75t_R _30944_ (.A1(_02484_),
    .A2(_11198_),
    .B(_11251_),
    .C(_11123_),
    .Y(_11252_));
 AOI21x1_ASAP7_75t_R _30945_ (.A1(_01491_),
    .A2(_11107_),
    .B(_11252_),
    .Y(_03915_));
 NOR2x1_ASAP7_75t_R _30946_ (.A(_01490_),
    .B(_02483_),
    .Y(_11253_));
 NOR2x1_ASAP7_75t_R _30947_ (.A(_09683_),
    .B(_11148_),
    .Y(_11254_));
 AO21x1_ASAP7_75t_R _30948_ (.A1(_11120_),
    .A2(_11253_),
    .B(_11254_),
    .Y(_11255_));
 AO21x1_ASAP7_75t_R _30949_ (.A1(_02483_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11256_));
 AOI22x1_ASAP7_75t_R _30950_ (.A1(_11123_),
    .A2(_11255_),
    .B1(_11256_),
    .B2(_01490_),
    .Y(_03916_));
 NAND2x1_ASAP7_75t_R _30951_ (.A(_09691_),
    .B(_11101_),
    .Y(_11257_));
 OA211x2_ASAP7_75t_R _30952_ (.A1(_02486_),
    .A2(_11156_),
    .B(_11257_),
    .C(_11123_),
    .Y(_11258_));
 AOI21x1_ASAP7_75t_R _30953_ (.A1(_01489_),
    .A2(_11107_),
    .B(_11258_),
    .Y(_03917_));
 AO21x1_ASAP7_75t_R _30954_ (.A1(_02485_),
    .A2(_11144_),
    .B(_11107_),
    .Y(_11259_));
 NAND2x1_ASAP7_75t_R _30955_ (.A(_01488_),
    .B(_11259_),
    .Y(_11260_));
 OR4x1_ASAP7_75t_R _30956_ (.A(_01488_),
    .B(_02485_),
    .C(_11107_),
    .D(_11101_),
    .Y(_11261_));
 OA211x2_ASAP7_75t_R _30957_ (.A1(_09698_),
    .A2(_11106_),
    .B(_11260_),
    .C(_11261_),
    .Y(_03918_));
 INVx5_ASAP7_75t_R _30958_ (.A(net3517),
    .Y(_11262_));
 NAND2x1_ASAP7_75t_R _30959_ (.A(_13514_),
    .B(_13522_),
    .Y(_11263_));
 AND4x2_ASAP7_75t_R _30960_ (.A(_11263_),
    .B(net305),
    .C(net310),
    .D(_05634_),
    .Y(_11264_));
 AND2x4_ASAP7_75t_R _30961_ (.A(_11155_),
    .B(_11264_),
    .Y(_11265_));
 NAND2x2_ASAP7_75t_R _30962_ (.A(_11141_),
    .B(_11265_),
    .Y(_11266_));
 INVx1_ASAP7_75t_R _30963_ (.A(_05657_),
    .Y(_11267_));
 OR3x4_ASAP7_75t_R _30964_ (.A(_11267_),
    .B(_07929_),
    .C(_11147_),
    .Y(_11268_));
 AND4x1_ASAP7_75t_R _30965_ (.A(net302),
    .B(_11077_),
    .C(_09443_),
    .D(_11264_),
    .Y(_11269_));
 AND4x2_ASAP7_75t_R _30966_ (.A(_01315_),
    .B(_05752_),
    .C(net3038),
    .D(_05746_),
    .Y(_11270_));
 AND3x1_ASAP7_75t_R _30967_ (.A(_06655_),
    .B(_07543_),
    .C(_11270_),
    .Y(_11271_));
 OR2x4_ASAP7_75t_R _30968_ (.A(_11269_),
    .B(_11271_),
    .Y(_11272_));
 OA211x2_ASAP7_75t_R _30969_ (.A1(_11262_),
    .A2(_11266_),
    .B(_11268_),
    .C(_11272_),
    .Y(_11273_));
 NAND2x2_ASAP7_75t_R _30970_ (.A(_11272_),
    .B(_11268_),
    .Y(_11274_));
 AND2x6_ASAP7_75t_R _30971_ (.A(_11096_),
    .B(_11265_),
    .Y(_11275_));
 TAPCELL_ASAP7_75t_R PHY_253 ();
 AO21x1_ASAP7_75t_R _30973_ (.A1(_11262_),
    .A2(_11275_),
    .B(_00660_),
    .Y(_11277_));
 OA22x2_ASAP7_75t_R _30974_ (.A1(\cs_registers_i.mhpmcounter[2][0] ),
    .A2(_11273_),
    .B1(_11274_),
    .B2(_11277_),
    .Y(_03919_));
 AND3x1_ASAP7_75t_R _30975_ (.A(_06655_),
    .B(_07543_),
    .C(_11270_),
    .Y(_11278_));
 AND3x1_ASAP7_75t_R _30976_ (.A(net310),
    .B(_05634_),
    .C(_05699_),
    .Y(_11279_));
 AND4x1_ASAP7_75t_R _30977_ (.A(net302),
    .B(_07438_),
    .C(_11279_),
    .D(_09443_),
    .Y(_11280_));
 OR3x1_ASAP7_75t_R _30978_ (.A(_11267_),
    .B(_07929_),
    .C(_11119_),
    .Y(_11281_));
 OA21x2_ASAP7_75t_R _30979_ (.A1(_11278_),
    .A2(_11280_),
    .B(_11281_),
    .Y(_11282_));
 TAPCELL_ASAP7_75t_R PHY_252 ();
 NAND2x2_ASAP7_75t_R _30981_ (.A(_11096_),
    .B(_11265_),
    .Y(_11284_));
 OAI21x1_ASAP7_75t_R _30982_ (.A1(_06951_),
    .A2(_06976_),
    .B(_09443_),
    .Y(_11285_));
 OR3x4_ASAP7_75t_R _30983_ (.A(_07929_),
    .B(_11285_),
    .C(_11099_),
    .Y(_11286_));
 TAPCELL_ASAP7_75t_R PHY_251 ();
 NOR2x1_ASAP7_75t_R _30985_ (.A(net3647),
    .B(_11286_),
    .Y(_11288_));
 AO21x1_ASAP7_75t_R _30986_ (.A1(_02392_),
    .A2(_11284_),
    .B(_11288_),
    .Y(_11289_));
 NAND2x1_ASAP7_75t_R _30987_ (.A(_11282_),
    .B(_11289_),
    .Y(_11290_));
 OA21x2_ASAP7_75t_R _30988_ (.A1(\cs_registers_i.mhpmcounter[2][1] ),
    .A2(_11282_),
    .B(_11290_),
    .Y(_03920_));
 TAPCELL_ASAP7_75t_R PHY_250 ();
 AND2x6_ASAP7_75t_R _30990_ (.A(_11141_),
    .B(_11265_),
    .Y(_11292_));
 TAPCELL_ASAP7_75t_R PHY_249 ();
 TAPCELL_ASAP7_75t_R PHY_248 ();
 NAND2x1_ASAP7_75t_R _30993_ (.A(_11159_),
    .B(_11275_),
    .Y(_11295_));
 TAPCELL_ASAP7_75t_R PHY_247 ();
 OA211x2_ASAP7_75t_R _30995_ (.A1(_02394_),
    .A2(_11292_),
    .B(_11295_),
    .C(_11282_),
    .Y(_11297_));
 AOI21x1_ASAP7_75t_R _30996_ (.A1(_01486_),
    .A2(_11274_),
    .B(_11297_),
    .Y(_03921_));
 INVx1_ASAP7_75t_R _30997_ (.A(_02393_),
    .Y(_11298_));
 NOR3x2_ASAP7_75t_R _30998_ (.B(_11111_),
    .C(_11119_),
    .Y(_11299_),
    .A(_07929_));
 TAPCELL_ASAP7_75t_R PHY_246 ();
 TAPCELL_ASAP7_75t_R PHY_245 ();
 OA21x2_ASAP7_75t_R _31001_ (.A1(_11298_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11302_));
 TAPCELL_ASAP7_75t_R PHY_244 ();
 TAPCELL_ASAP7_75t_R PHY_243 ();
 AND3x1_ASAP7_75t_R _31004_ (.A(_01485_),
    .B(_11298_),
    .C(_11286_),
    .Y(_11305_));
 AOI21x1_ASAP7_75t_R _31005_ (.A1(net3563),
    .A2(_11292_),
    .B(_11305_),
    .Y(_11306_));
 TAPCELL_ASAP7_75t_R PHY_242 ();
 OAI22x1_ASAP7_75t_R _31007_ (.A1(_01485_),
    .A2(_11302_),
    .B1(_11306_),
    .B2(_11274_),
    .Y(_03922_));
 OR2x2_ASAP7_75t_R _31008_ (.A(net3378),
    .B(_11284_),
    .Y(_11308_));
 OA211x2_ASAP7_75t_R _31009_ (.A1(_02396_),
    .A2(_11292_),
    .B(_11308_),
    .C(_11282_),
    .Y(_11309_));
 AOI21x1_ASAP7_75t_R _31010_ (.A1(_01484_),
    .A2(_11274_),
    .B(_11309_),
    .Y(_03923_));
 INVx1_ASAP7_75t_R _31011_ (.A(_02395_),
    .Y(_11310_));
 AND3x1_ASAP7_75t_R _31012_ (.A(_01483_),
    .B(_11310_),
    .C(_11284_),
    .Y(_11311_));
 AOI21x1_ASAP7_75t_R _31013_ (.A1(net3632),
    .A2(_11275_),
    .B(_11311_),
    .Y(_11312_));
 TAPCELL_ASAP7_75t_R PHY_241 ();
 OA21x2_ASAP7_75t_R _31015_ (.A1(_11310_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11314_));
 OAI22x1_ASAP7_75t_R _31016_ (.A1(_11274_),
    .A2(_11312_),
    .B1(_11314_),
    .B2(_01483_),
    .Y(_03924_));
 NAND2x1_ASAP7_75t_R _31017_ (.A(_09504_),
    .B(_11299_),
    .Y(_11315_));
 OA211x2_ASAP7_75t_R _31018_ (.A1(_02398_),
    .A2(_11292_),
    .B(_11315_),
    .C(_11282_),
    .Y(_11316_));
 AOI21x1_ASAP7_75t_R _31019_ (.A1(_01482_),
    .A2(_11274_),
    .B(_11316_),
    .Y(_03925_));
 INVx1_ASAP7_75t_R _31020_ (.A(_02397_),
    .Y(_11317_));
 AND3x1_ASAP7_75t_R _31021_ (.A(_01481_),
    .B(_11317_),
    .C(_11266_),
    .Y(_11318_));
 AOI21x1_ASAP7_75t_R _31022_ (.A1(net3654),
    .A2(_11292_),
    .B(_11318_),
    .Y(_11319_));
 OA21x2_ASAP7_75t_R _31023_ (.A1(_11317_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11320_));
 OAI22x1_ASAP7_75t_R _31024_ (.A1(_11274_),
    .A2(_11319_),
    .B1(_11320_),
    .B2(_01481_),
    .Y(_03926_));
 NAND2x1_ASAP7_75t_R _31025_ (.A(_09518_),
    .B(_11299_),
    .Y(_11321_));
 OA211x2_ASAP7_75t_R _31026_ (.A1(_02400_),
    .A2(_11292_),
    .B(_11321_),
    .C(_11282_),
    .Y(_11322_));
 AOI21x1_ASAP7_75t_R _31027_ (.A1(_01480_),
    .A2(_11274_),
    .B(_11322_),
    .Y(_03927_));
 INVx1_ASAP7_75t_R _31028_ (.A(_02399_),
    .Y(_11323_));
 OA21x2_ASAP7_75t_R _31029_ (.A1(_11323_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11324_));
 AND3x1_ASAP7_75t_R _31030_ (.A(_01479_),
    .B(_11323_),
    .C(_11286_),
    .Y(_11325_));
 AOI21x1_ASAP7_75t_R _31031_ (.A1(net3716),
    .A2(_11292_),
    .B(_11325_),
    .Y(_11326_));
 OAI22x1_ASAP7_75t_R _31032_ (.A1(_01479_),
    .A2(_11324_),
    .B1(_11326_),
    .B2(_11274_),
    .Y(_03928_));
 NOR2x2_ASAP7_75t_R _31033_ (.A(_07929_),
    .B(_11285_),
    .Y(_11327_));
 AO21x1_ASAP7_75t_R _31034_ (.A1(_11155_),
    .A2(_11327_),
    .B(_02402_),
    .Y(_11328_));
 NAND2x1_ASAP7_75t_R _31035_ (.A(_09531_),
    .B(_11275_),
    .Y(_11329_));
 AND3x1_ASAP7_75t_R _31036_ (.A(_11282_),
    .B(_11328_),
    .C(_11329_),
    .Y(_11330_));
 AOI21x1_ASAP7_75t_R _31037_ (.A1(_01478_),
    .A2(_11274_),
    .B(_11330_),
    .Y(_03929_));
 INVx1_ASAP7_75t_R _31038_ (.A(_02401_),
    .Y(_11331_));
 OA21x2_ASAP7_75t_R _31039_ (.A1(_11331_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11332_));
 AND3x1_ASAP7_75t_R _31040_ (.A(_01477_),
    .B(_11331_),
    .C(_11286_),
    .Y(_11333_));
 AOI21x1_ASAP7_75t_R _31041_ (.A1(_09538_),
    .A2(_11292_),
    .B(_11333_),
    .Y(_11334_));
 OAI22x1_ASAP7_75t_R _31042_ (.A1(_01477_),
    .A2(_11332_),
    .B1(_11334_),
    .B2(_11274_),
    .Y(_03930_));
 AND2x4_ASAP7_75t_R _31043_ (.A(_11155_),
    .B(_11327_),
    .Y(_11335_));
 NAND2x2_ASAP7_75t_R _31044_ (.A(net3673),
    .B(_11335_),
    .Y(_11336_));
 OA211x2_ASAP7_75t_R _31045_ (.A1(_02404_),
    .A2(_11292_),
    .B(_11336_),
    .C(_11282_),
    .Y(_11337_));
 AOI21x1_ASAP7_75t_R _31046_ (.A1(_01476_),
    .A2(_11274_),
    .B(_11337_),
    .Y(_03931_));
 INVx1_ASAP7_75t_R _31047_ (.A(_02403_),
    .Y(_11338_));
 AND3x1_ASAP7_75t_R _31048_ (.A(_01475_),
    .B(_11338_),
    .C(_11286_),
    .Y(_11339_));
 AOI21x1_ASAP7_75t_R _31049_ (.A1(net3707),
    .A2(_11292_),
    .B(_11339_),
    .Y(_11340_));
 OA21x2_ASAP7_75t_R _31050_ (.A1(_11338_),
    .A2(_11292_),
    .B(_11282_),
    .Y(_11341_));
 OAI22x1_ASAP7_75t_R _31051_ (.A1(_11274_),
    .A2(_11340_),
    .B1(_11341_),
    .B2(_01475_),
    .Y(_03932_));
 NAND2x1_ASAP7_75t_R _31052_ (.A(net3541),
    .B(_11275_),
    .Y(_11342_));
 OA211x2_ASAP7_75t_R _31053_ (.A1(_02406_),
    .A2(_11292_),
    .B(_11342_),
    .C(_11282_),
    .Y(_11343_));
 AOI21x1_ASAP7_75t_R _31054_ (.A1(_01474_),
    .A2(_11274_),
    .B(_11343_),
    .Y(_03933_));
 INVx1_ASAP7_75t_R _31055_ (.A(_02405_),
    .Y(_11344_));
 OA21x2_ASAP7_75t_R _31056_ (.A1(_11344_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11345_));
 AND3x1_ASAP7_75t_R _31057_ (.A(_01473_),
    .B(_11344_),
    .C(_11286_),
    .Y(_11346_));
 AOI21x1_ASAP7_75t_R _31058_ (.A1(net3747),
    .A2(_11292_),
    .B(_11346_),
    .Y(_11347_));
 OAI22x1_ASAP7_75t_R _31059_ (.A1(_01473_),
    .A2(_11345_),
    .B1(_11347_),
    .B2(_11274_),
    .Y(_03934_));
 AO21x1_ASAP7_75t_R _31060_ (.A1(_11155_),
    .A2(_11327_),
    .B(_02408_),
    .Y(_11348_));
 NAND2x2_ASAP7_75t_R _31061_ (.A(net3604),
    .B(_11275_),
    .Y(_11349_));
 AND3x1_ASAP7_75t_R _31062_ (.A(_11282_),
    .B(_11348_),
    .C(_11349_),
    .Y(_11350_));
 AOI21x1_ASAP7_75t_R _31063_ (.A1(_01472_),
    .A2(_11274_),
    .B(_11350_),
    .Y(_03935_));
 INVx1_ASAP7_75t_R _31064_ (.A(_02407_),
    .Y(_11351_));
 OA21x2_ASAP7_75t_R _31065_ (.A1(_11351_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11352_));
 AND3x1_ASAP7_75t_R _31066_ (.A(_01471_),
    .B(_11351_),
    .C(_11286_),
    .Y(_11353_));
 AOI21x1_ASAP7_75t_R _31067_ (.A1(net3660),
    .A2(_11335_),
    .B(_11353_),
    .Y(_11354_));
 OAI22x1_ASAP7_75t_R _31068_ (.A1(_01471_),
    .A2(_11352_),
    .B1(_11354_),
    .B2(_11274_),
    .Y(_03936_));
 AO21x1_ASAP7_75t_R _31069_ (.A1(_11155_),
    .A2(_11327_),
    .B(_02410_),
    .Y(_11355_));
 OR2x2_ASAP7_75t_R _31070_ (.A(net3571),
    .B(_11284_),
    .Y(_11356_));
 AND3x1_ASAP7_75t_R _31071_ (.A(_11282_),
    .B(_11355_),
    .C(_11356_),
    .Y(_11357_));
 AOI21x1_ASAP7_75t_R _31072_ (.A1(_01470_),
    .A2(_11274_),
    .B(_11357_),
    .Y(_03937_));
 INVx1_ASAP7_75t_R _31073_ (.A(_02409_),
    .Y(_11358_));
 AND3x1_ASAP7_75t_R _31074_ (.A(_01469_),
    .B(_11358_),
    .C(_11286_),
    .Y(_11359_));
 AOI21x1_ASAP7_75t_R _31075_ (.A1(net3721),
    .A2(_11292_),
    .B(_11359_),
    .Y(_11360_));
 OA21x2_ASAP7_75t_R _31076_ (.A1(_11358_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11361_));
 OAI22x1_ASAP7_75t_R _31077_ (.A1(_11274_),
    .A2(_11360_),
    .B1(_11361_),
    .B2(_01469_),
    .Y(_03938_));
 OR2x2_ASAP7_75t_R _31078_ (.A(_09615_),
    .B(_11266_),
    .Y(_11362_));
 OA211x2_ASAP7_75t_R _31079_ (.A1(_02412_),
    .A2(_11292_),
    .B(_11362_),
    .C(_11282_),
    .Y(_11363_));
 AOI21x1_ASAP7_75t_R _31080_ (.A1(_01468_),
    .A2(_11274_),
    .B(_11363_),
    .Y(_03939_));
 INVx1_ASAP7_75t_R _31081_ (.A(_02411_),
    .Y(_11364_));
 OAI21x1_ASAP7_75t_R _31082_ (.A1(_11364_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11365_));
 AND3x1_ASAP7_75t_R _31083_ (.A(_01467_),
    .B(_11364_),
    .C(_11286_),
    .Y(_11366_));
 AO21x1_ASAP7_75t_R _31084_ (.A1(_09623_),
    .A2(_11335_),
    .B(_11366_),
    .Y(_11367_));
 AO22x1_ASAP7_75t_R _31085_ (.A1(_06021_),
    .A2(_11365_),
    .B1(_11367_),
    .B2(_11282_),
    .Y(_03940_));
 NAND2x1_ASAP7_75t_R _31086_ (.A(_09631_),
    .B(_11275_),
    .Y(_11368_));
 OA211x2_ASAP7_75t_R _31087_ (.A1(_02414_),
    .A2(_11292_),
    .B(_11368_),
    .C(_11282_),
    .Y(_11369_));
 AOI21x1_ASAP7_75t_R _31088_ (.A1(_01466_),
    .A2(_11274_),
    .B(_11369_),
    .Y(_03941_));
 INVx1_ASAP7_75t_R _31089_ (.A(_02413_),
    .Y(_11370_));
 AND3x1_ASAP7_75t_R _31090_ (.A(_01465_),
    .B(_11370_),
    .C(_11284_),
    .Y(_11371_));
 AOI21x1_ASAP7_75t_R _31091_ (.A1(_09638_),
    .A2(_11275_),
    .B(_11371_),
    .Y(_11372_));
 OA21x2_ASAP7_75t_R _31092_ (.A1(_11370_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11373_));
 OAI22x1_ASAP7_75t_R _31093_ (.A1(_11274_),
    .A2(_11372_),
    .B1(_11373_),
    .B2(_01465_),
    .Y(_03942_));
 NOR2x1_ASAP7_75t_R _31094_ (.A(_02416_),
    .B(_11275_),
    .Y(_11374_));
 AND5x2_ASAP7_75t_R _31095_ (.A(_09442_),
    .B(_07530_),
    .C(_09443_),
    .D(_09647_),
    .E(_11100_),
    .Y(_11375_));
 OR2x2_ASAP7_75t_R _31096_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(_11282_),
    .Y(_11376_));
 OA31x2_ASAP7_75t_R _31097_ (.A1(_11274_),
    .A2(_11374_),
    .A3(_11375_),
    .B1(_11376_),
    .Y(_03943_));
 INVx1_ASAP7_75t_R _31098_ (.A(_02415_),
    .Y(_11377_));
 OA21x2_ASAP7_75t_R _31099_ (.A1(_11377_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11378_));
 AND3x1_ASAP7_75t_R _31100_ (.A(_01463_),
    .B(_11377_),
    .C(_11286_),
    .Y(_11379_));
 AOI21x1_ASAP7_75t_R _31101_ (.A1(net3639),
    .A2(_11292_),
    .B(_11379_),
    .Y(_11380_));
 OAI22x1_ASAP7_75t_R _31102_ (.A1(_01463_),
    .A2(_11378_),
    .B1(_11380_),
    .B2(_11274_),
    .Y(_03944_));
 OR2x2_ASAP7_75t_R _31103_ (.A(_09661_),
    .B(_11284_),
    .Y(_11381_));
 OA21x2_ASAP7_75t_R _31104_ (.A1(_02418_),
    .A2(_11292_),
    .B(_11381_),
    .Y(_11382_));
 NAND2x1_ASAP7_75t_R _31105_ (.A(_11282_),
    .B(_11382_),
    .Y(_11383_));
 OA21x2_ASAP7_75t_R _31106_ (.A1(\cs_registers_i.mhpmcounter[2][26] ),
    .A2(_11282_),
    .B(_11383_),
    .Y(_03945_));
 INVx1_ASAP7_75t_R _31107_ (.A(_02417_),
    .Y(_11384_));
 OA21x2_ASAP7_75t_R _31108_ (.A1(_11384_),
    .A2(_11292_),
    .B(_11282_),
    .Y(_11385_));
 AND3x1_ASAP7_75t_R _31109_ (.A(_01461_),
    .B(_11384_),
    .C(_11286_),
    .Y(_11386_));
 AOI21x1_ASAP7_75t_R _31110_ (.A1(net3594),
    .A2(_11292_),
    .B(_11386_),
    .Y(_11387_));
 OAI22x1_ASAP7_75t_R _31111_ (.A1(_01461_),
    .A2(_11385_),
    .B1(_11387_),
    .B2(_11274_),
    .Y(_03946_));
 NAND2x1_ASAP7_75t_R _31112_ (.A(_09676_),
    .B(_11275_),
    .Y(_11388_));
 OA211x2_ASAP7_75t_R _31113_ (.A1(_02420_),
    .A2(_11292_),
    .B(_11388_),
    .C(_11282_),
    .Y(_11389_));
 AOI21x1_ASAP7_75t_R _31114_ (.A1(_01460_),
    .A2(_11274_),
    .B(_11389_),
    .Y(_03947_));
 INVx1_ASAP7_75t_R _31115_ (.A(_02419_),
    .Y(_11390_));
 AND3x1_ASAP7_75t_R _31116_ (.A(_01459_),
    .B(_11390_),
    .C(_11286_),
    .Y(_11391_));
 AO21x1_ASAP7_75t_R _31117_ (.A1(_09683_),
    .A2(_11292_),
    .B(_11391_),
    .Y(_11392_));
 OAI21x1_ASAP7_75t_R _31118_ (.A1(_11390_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11393_));
 AO32x1_ASAP7_75t_R _31119_ (.A1(_11272_),
    .A2(_11268_),
    .A3(_11392_),
    .B1(_11393_),
    .B2(_06025_),
    .Y(_03948_));
 NAND2x1_ASAP7_75t_R _31120_ (.A(_09691_),
    .B(_11335_),
    .Y(_11394_));
 OA211x2_ASAP7_75t_R _31121_ (.A1(_02422_),
    .A2(_11292_),
    .B(_11394_),
    .C(_11282_),
    .Y(_11395_));
 AOI21x1_ASAP7_75t_R _31122_ (.A1(_01458_),
    .A2(_11274_),
    .B(_11395_),
    .Y(_03949_));
 INVx1_ASAP7_75t_R _31123_ (.A(_02421_),
    .Y(_11396_));
 AND3x1_ASAP7_75t_R _31124_ (.A(_01457_),
    .B(_11396_),
    .C(_11286_),
    .Y(_11397_));
 AO21x1_ASAP7_75t_R _31125_ (.A1(_09698_),
    .A2(_11335_),
    .B(_11397_),
    .Y(_11398_));
 TAPCELL_ASAP7_75t_R PHY_240 ();
 OAI21x1_ASAP7_75t_R _31127_ (.A1(_11396_),
    .A2(_11299_),
    .B(_11282_),
    .Y(_11400_));
 INVx1_ASAP7_75t_R _31128_ (.A(_01457_),
    .Y(_11401_));
 AO32x1_ASAP7_75t_R _31129_ (.A1(_11272_),
    .A2(_11268_),
    .A3(_11398_),
    .B1(_11400_),
    .B2(_11401_),
    .Y(_03950_));
 AND3x2_ASAP7_75t_R _31130_ (.A(_05693_),
    .B(_06960_),
    .C(_11130_),
    .Y(_11402_));
 NAND2x2_ASAP7_75t_R _31131_ (.A(_11402_),
    .B(_11141_),
    .Y(_11403_));
 NAND2x1_ASAP7_75t_R _31132_ (.A(_01456_),
    .B(_11403_),
    .Y(_11404_));
 OAI21x1_ASAP7_75t_R _31133_ (.A1(_06212_),
    .A2(_06216_),
    .B(_06385_),
    .Y(_11405_));
 AND3x4_ASAP7_75t_R _31134_ (.A(_06271_),
    .B(_06932_),
    .C(_11405_),
    .Y(_11406_));
 AO21x2_ASAP7_75t_R _31135_ (.A1(_06230_),
    .A2(_06931_),
    .B(_05724_),
    .Y(_11407_));
 OR2x6_ASAP7_75t_R _31136_ (.A(_11406_),
    .B(_11407_),
    .Y(_11408_));
 TAPCELL_ASAP7_75t_R PHY_239 ();
 TAPCELL_ASAP7_75t_R PHY_238 ();
 OR4x1_ASAP7_75t_R _31139_ (.A(_07740_),
    .B(_11285_),
    .C(_09538_),
    .D(_09548_),
    .Y(_11411_));
 AND3x1_ASAP7_75t_R _31140_ (.A(_06301_),
    .B(_11408_),
    .C(_11411_),
    .Y(_11412_));
 TAPCELL_ASAP7_75t_R PHY_237 ();
 OR3x4_ASAP7_75t_R _31142_ (.A(_01718_),
    .B(_06221_),
    .C(_06300_),
    .Y(_11414_));
 TAPCELL_ASAP7_75t_R PHY_236 ();
 OAI22x1_ASAP7_75t_R _31144_ (.A1(_02140_),
    .A2(_11408_),
    .B1(_11414_),
    .B2(_02107_),
    .Y(_11416_));
 AO21x1_ASAP7_75t_R _31145_ (.A1(_11404_),
    .A2(_11412_),
    .B(_11416_),
    .Y(_03951_));
 INVx1_ASAP7_75t_R _31146_ (.A(_01455_),
    .Y(_11417_));
 AO21x1_ASAP7_75t_R _31147_ (.A1(_11402_),
    .A2(_11141_),
    .B(_11417_),
    .Y(_11418_));
 OAI22x1_ASAP7_75t_R _31148_ (.A1(_17810_),
    .A2(_11408_),
    .B1(_11414_),
    .B2(_02106_),
    .Y(_11419_));
 AO21x1_ASAP7_75t_R _31149_ (.A1(_11412_),
    .A2(_11418_),
    .B(_11419_),
    .Y(_03952_));
 AO21x1_ASAP7_75t_R _31150_ (.A1(_06887_),
    .A2(_02105_),
    .B(_06301_),
    .Y(_11420_));
 INVx1_ASAP7_75t_R _31151_ (.A(_11403_),
    .Y(_11421_));
 INVx2_ASAP7_75t_R _31152_ (.A(_11406_),
    .Y(_11422_));
 NAND2x2_ASAP7_75t_R _31153_ (.A(_11408_),
    .B(_11414_),
    .Y(_11423_));
 OA21x2_ASAP7_75t_R _31154_ (.A1(_02105_),
    .A2(_11422_),
    .B(_11423_),
    .Y(_11424_));
 OR3x1_ASAP7_75t_R _31155_ (.A(_01454_),
    .B(_11421_),
    .C(_11424_),
    .Y(_11425_));
 OA211x2_ASAP7_75t_R _31156_ (.A1(_01453_),
    .A2(_11408_),
    .B(_11420_),
    .C(_11425_),
    .Y(_11426_));
 OAI21x1_ASAP7_75t_R _31157_ (.A1(_11182_),
    .A2(_11403_),
    .B(_11426_),
    .Y(_03953_));
 AO21x1_ASAP7_75t_R _31158_ (.A1(_11402_),
    .A2(_11141_),
    .B(_06236_),
    .Y(_11427_));
 OA211x2_ASAP7_75t_R _31159_ (.A1(net3544),
    .A2(_11403_),
    .B(_11427_),
    .C(_11408_),
    .Y(_11428_));
 NOR2x1_ASAP7_75t_R _31160_ (.A(_01454_),
    .B(_06301_),
    .Y(_11429_));
 AO21x1_ASAP7_75t_R _31161_ (.A1(_06301_),
    .A2(_11428_),
    .B(_11429_),
    .Y(_03954_));
 INVx1_ASAP7_75t_R _31162_ (.A(_01452_),
    .Y(_11430_));
 NAND2x2_ASAP7_75t_R _31163_ (.A(_05776_),
    .B(_05777_),
    .Y(_11431_));
 TAPCELL_ASAP7_75t_R PHY_235 ();
 TAPCELL_ASAP7_75t_R PHY_234 ();
 TAPCELL_ASAP7_75t_R PHY_233 ();
 AO21x1_ASAP7_75t_R _31167_ (.A1(_05454_),
    .A2(_05943_),
    .B(_13886_),
    .Y(_11435_));
 TAPCELL_ASAP7_75t_R PHY_232 ();
 OA211x2_ASAP7_75t_R _31169_ (.A1(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A2(_06752_),
    .B(_11435_),
    .C(_05779_),
    .Y(_11437_));
 AO21x1_ASAP7_75t_R _31170_ (.A1(_11430_),
    .A2(_11431_),
    .B(_11437_),
    .Y(_03955_));
 INVx1_ASAP7_75t_R _31171_ (.A(_01451_),
    .Y(_11438_));
 AO21x1_ASAP7_75t_R _31172_ (.A1(_05454_),
    .A2(_05943_),
    .B(net2252),
    .Y(_11439_));
 OA211x2_ASAP7_75t_R _31173_ (.A1(net296),
    .A2(_06752_),
    .B(_11439_),
    .C(_05779_),
    .Y(_11440_));
 AO21x1_ASAP7_75t_R _31174_ (.A1(_11438_),
    .A2(_11431_),
    .B(_11440_),
    .Y(_03956_));
 TAPCELL_ASAP7_75t_R PHY_231 ();
 TAPCELL_ASAP7_75t_R PHY_230 ();
 AO21x1_ASAP7_75t_R _31177_ (.A1(_05454_),
    .A2(_05943_),
    .B(_06838_),
    .Y(_11443_));
 OA211x2_ASAP7_75t_R _31178_ (.A1(_05792_),
    .A2(_06752_),
    .B(_11443_),
    .C(_05779_),
    .Y(_11444_));
 AOI21x1_ASAP7_75t_R _31179_ (.A1(_01450_),
    .A2(_11431_),
    .B(_11444_),
    .Y(_03957_));
 TAPCELL_ASAP7_75t_R PHY_229 ();
 NAND2x1_ASAP7_75t_R _31181_ (.A(_14233_),
    .B(_06752_),
    .Y(_11446_));
 OA211x2_ASAP7_75t_R _31182_ (.A1(_06317_),
    .A2(_06752_),
    .B(_11446_),
    .C(_05779_),
    .Y(_11447_));
 AOI21x1_ASAP7_75t_R _31183_ (.A1(_01449_),
    .A2(_11431_),
    .B(_11447_),
    .Y(_03958_));
 NAND2x1_ASAP7_75t_R _31184_ (.A(net2221),
    .B(_06752_),
    .Y(_11448_));
 OA211x2_ASAP7_75t_R _31185_ (.A1(_05791_),
    .A2(_06752_),
    .B(_11448_),
    .C(_05779_),
    .Y(_11449_));
 AOI21x1_ASAP7_75t_R _31186_ (.A1(_01448_),
    .A2(_11431_),
    .B(_11449_),
    .Y(_03959_));
 AO21x1_ASAP7_75t_R _31187_ (.A1(_05454_),
    .A2(_05943_),
    .B(_14355_),
    .Y(_11450_));
 OA211x2_ASAP7_75t_R _31188_ (.A1(net176),
    .A2(_06752_),
    .B(_11450_),
    .C(_05779_),
    .Y(_11451_));
 AO21x1_ASAP7_75t_R _31189_ (.A1(_15106_),
    .A2(_11431_),
    .B(_11451_),
    .Y(_03960_));
 AO21x1_ASAP7_75t_R _31190_ (.A1(_05454_),
    .A2(_05943_),
    .B(_05567_),
    .Y(_11452_));
 OA211x2_ASAP7_75t_R _31191_ (.A1(_05793_),
    .A2(_06752_),
    .B(_11452_),
    .C(_05779_),
    .Y(_11453_));
 AOI21x1_ASAP7_75t_R _31192_ (.A1(_01446_),
    .A2(_11431_),
    .B(_11453_),
    .Y(_03961_));
 INVx1_ASAP7_75t_R _31193_ (.A(_01445_),
    .Y(_11454_));
 AO21x1_ASAP7_75t_R _31194_ (.A1(_05454_),
    .A2(_05943_),
    .B(_14479_),
    .Y(_11455_));
 OA211x2_ASAP7_75t_R _31195_ (.A1(net178),
    .A2(_06752_),
    .B(_11455_),
    .C(_05779_),
    .Y(_11456_));
 AO21x1_ASAP7_75t_R _31196_ (.A1(_11454_),
    .A2(_11431_),
    .B(_11456_),
    .Y(_03962_));
 INVx1_ASAP7_75t_R _31197_ (.A(_01444_),
    .Y(_11457_));
 AO21x1_ASAP7_75t_R _31198_ (.A1(_05454_),
    .A2(_05943_),
    .B(_14539_),
    .Y(_11458_));
 OA211x2_ASAP7_75t_R _31199_ (.A1(net179),
    .A2(_06752_),
    .B(_11458_),
    .C(_05779_),
    .Y(_11459_));
 AO21x1_ASAP7_75t_R _31200_ (.A1(_11457_),
    .A2(_11431_),
    .B(_11459_),
    .Y(_03963_));
 AO21x1_ASAP7_75t_R _31201_ (.A1(_05454_),
    .A2(_05943_),
    .B(_14597_),
    .Y(_11460_));
 OA211x2_ASAP7_75t_R _31202_ (.A1(net180),
    .A2(_06752_),
    .B(_11460_),
    .C(_05779_),
    .Y(_11461_));
 AO21x1_ASAP7_75t_R _31203_ (.A1(_15283_),
    .A2(_11431_),
    .B(_11461_),
    .Y(_03964_));
 AO21x1_ASAP7_75t_R _31204_ (.A1(_05454_),
    .A2(_05943_),
    .B(_14651_),
    .Y(_11462_));
 OA211x2_ASAP7_75t_R _31205_ (.A1(_05797_),
    .A2(_06752_),
    .B(_11462_),
    .C(_05779_),
    .Y(_11463_));
 AOI21x1_ASAP7_75t_R _31206_ (.A1(_01442_),
    .A2(_11431_),
    .B(_11463_),
    .Y(_03965_));
 AO21x1_ASAP7_75t_R _31207_ (.A1(_05454_),
    .A2(_05943_),
    .B(_05898_),
    .Y(_11464_));
 OA211x2_ASAP7_75t_R _31208_ (.A1(net152),
    .A2(_06752_),
    .B(_11464_),
    .C(_05779_),
    .Y(_11465_));
 AO21x1_ASAP7_75t_R _31209_ (.A1(_15405_),
    .A2(_11431_),
    .B(_11465_),
    .Y(_03966_));
 NAND2x1_ASAP7_75t_R _31210_ (.A(_15487_),
    .B(_06752_),
    .Y(_11466_));
 OA211x2_ASAP7_75t_R _31211_ (.A1(_05796_),
    .A2(_06752_),
    .B(_11466_),
    .C(_05779_),
    .Y(_11467_));
 AOI21x1_ASAP7_75t_R _31212_ (.A1(_02221_),
    .A2(_11431_),
    .B(_11467_),
    .Y(_03967_));
 OR2x2_ASAP7_75t_R _31213_ (.A(_15590_),
    .B(_05944_),
    .Y(_11468_));
 OA211x2_ASAP7_75t_R _31214_ (.A1(_06428_),
    .A2(_06752_),
    .B(_11468_),
    .C(_05779_),
    .Y(_11469_));
 AOI21x1_ASAP7_75t_R _31215_ (.A1(_02220_),
    .A2(_11431_),
    .B(_11469_),
    .Y(_03968_));
 OR2x2_ASAP7_75t_R _31216_ (.A(_15723_),
    .B(_05944_),
    .Y(_11470_));
 OA211x2_ASAP7_75t_R _31217_ (.A1(_15778_),
    .A2(_06752_),
    .B(_11470_),
    .C(_05779_),
    .Y(_11471_));
 AOI21x1_ASAP7_75t_R _31218_ (.A1(_02219_),
    .A2(_11431_),
    .B(_11471_),
    .Y(_03969_));
 TAPCELL_ASAP7_75t_R PHY_228 ();
 NAND2x1_ASAP7_75t_R _31220_ (.A(net156),
    .B(_05944_),
    .Y(_11473_));
 OA211x2_ASAP7_75t_R _31221_ (.A1(_15839_),
    .A2(_05944_),
    .B(_11473_),
    .C(_05779_),
    .Y(_11474_));
 AOI21x1_ASAP7_75t_R _31222_ (.A1(_02218_),
    .A2(_11431_),
    .B(_11474_),
    .Y(_03970_));
 NAND2x1_ASAP7_75t_R _31223_ (.A(net157),
    .B(_05944_),
    .Y(_11475_));
 TAPCELL_ASAP7_75t_R PHY_227 ();
 OA211x2_ASAP7_75t_R _31225_ (.A1(_15972_),
    .A2(_05944_),
    .B(_11475_),
    .C(_05779_),
    .Y(_11477_));
 AOI21x1_ASAP7_75t_R _31226_ (.A1(_02217_),
    .A2(_11431_),
    .B(_11477_),
    .Y(_03971_));
 TAPCELL_ASAP7_75t_R PHY_226 ();
 NAND2x1_ASAP7_75t_R _31228_ (.A(net2255),
    .B(_05944_),
    .Y(_11479_));
 OA211x2_ASAP7_75t_R _31229_ (.A1(_16087_),
    .A2(_05944_),
    .B(_11479_),
    .C(_05779_),
    .Y(_11480_));
 AOI21x1_ASAP7_75t_R _31230_ (.A1(_02216_),
    .A2(_11431_),
    .B(_11480_),
    .Y(_03972_));
 NAND2x1_ASAP7_75t_R _31231_ (.A(_16213_),
    .B(_06752_),
    .Y(_11481_));
 OA211x2_ASAP7_75t_R _31232_ (.A1(_16263_),
    .A2(_06752_),
    .B(_11481_),
    .C(_05779_),
    .Y(_11482_));
 AOI21x1_ASAP7_75t_R _31233_ (.A1(_02215_),
    .A2(_11431_),
    .B(_11482_),
    .Y(_03973_));
 NAND2x1_ASAP7_75t_R _31234_ (.A(_16324_),
    .B(_06752_),
    .Y(_11483_));
 OA211x2_ASAP7_75t_R _31235_ (.A1(_06472_),
    .A2(_06752_),
    .B(_11483_),
    .C(_05779_),
    .Y(_11484_));
 AOI21x1_ASAP7_75t_R _31236_ (.A1(_02214_),
    .A2(_11431_),
    .B(_11484_),
    .Y(_03974_));
 NAND2x1_ASAP7_75t_R _31237_ (.A(_16456_),
    .B(_06752_),
    .Y(_11485_));
 OA211x2_ASAP7_75t_R _31238_ (.A1(_16509_),
    .A2(_06752_),
    .B(_11485_),
    .C(_05779_),
    .Y(_11486_));
 AOI21x1_ASAP7_75t_R _31239_ (.A1(_02213_),
    .A2(_11431_),
    .B(_11486_),
    .Y(_03975_));
 NAND2x1_ASAP7_75t_R _31240_ (.A(net162),
    .B(_05944_),
    .Y(_11487_));
 OA211x2_ASAP7_75t_R _31241_ (.A1(net2181),
    .A2(_05944_),
    .B(_11487_),
    .C(_05779_),
    .Y(_11488_));
 AOI21x1_ASAP7_75t_R _31242_ (.A1(_02212_),
    .A2(_11431_),
    .B(_11488_),
    .Y(_03976_));
 NAND2x1_ASAP7_75t_R _31243_ (.A(net163),
    .B(_05944_),
    .Y(_11489_));
 OA211x2_ASAP7_75t_R _31244_ (.A1(_16679_),
    .A2(_05944_),
    .B(_11489_),
    .C(_05779_),
    .Y(_11490_));
 AOI21x1_ASAP7_75t_R _31245_ (.A1(_02211_),
    .A2(_11431_),
    .B(_11490_),
    .Y(_03977_));
 NAND2x1_ASAP7_75t_R _31246_ (.A(_04576_),
    .B(_06752_),
    .Y(_11491_));
 OA211x2_ASAP7_75t_R _31247_ (.A1(_06498_),
    .A2(_06752_),
    .B(_11491_),
    .C(_05779_),
    .Y(_11492_));
 AOI21x1_ASAP7_75t_R _31248_ (.A1(_02210_),
    .A2(_11431_),
    .B(_11492_),
    .Y(_03978_));
 NAND2x1_ASAP7_75t_R _31249_ (.A(_04697_),
    .B(_06752_),
    .Y(_11493_));
 OA211x2_ASAP7_75t_R _31250_ (.A1(_04747_),
    .A2(_06752_),
    .B(_11493_),
    .C(_05779_),
    .Y(_11494_));
 AOI21x1_ASAP7_75t_R _31251_ (.A1(_02209_),
    .A2(_11431_),
    .B(_11494_),
    .Y(_03979_));
 OR2x2_ASAP7_75t_R _31252_ (.A(_04808_),
    .B(_05944_),
    .Y(_11495_));
 OA211x2_ASAP7_75t_R _31253_ (.A1(_06511_),
    .A2(_06752_),
    .B(_11495_),
    .C(_05779_),
    .Y(_11496_));
 AOI21x1_ASAP7_75t_R _31254_ (.A1(_02208_),
    .A2(_11431_),
    .B(_11496_),
    .Y(_03980_));
 NAND2x1_ASAP7_75t_R _31255_ (.A(_04916_),
    .B(_06752_),
    .Y(_11497_));
 OA211x2_ASAP7_75t_R _31256_ (.A1(_04968_),
    .A2(_06752_),
    .B(_11497_),
    .C(_05779_),
    .Y(_11498_));
 AOI21x1_ASAP7_75t_R _31257_ (.A1(_02207_),
    .A2(_11431_),
    .B(_11498_),
    .Y(_03981_));
 NAND2x1_ASAP7_75t_R _31258_ (.A(net2158),
    .B(_05944_),
    .Y(_11499_));
 OA211x2_ASAP7_75t_R _31259_ (.A1(_05028_),
    .A2(_05944_),
    .B(_11499_),
    .C(_05779_),
    .Y(_11500_));
 AOI21x1_ASAP7_75t_R _31260_ (.A1(_02206_),
    .A2(_11431_),
    .B(_11500_),
    .Y(_03982_));
 NAND2x1_ASAP7_75t_R _31261_ (.A(net169),
    .B(_05944_),
    .Y(_11501_));
 OA211x2_ASAP7_75t_R _31262_ (.A1(_05136_),
    .A2(_05944_),
    .B(_11501_),
    .C(_05779_),
    .Y(_11502_));
 AOI21x1_ASAP7_75t_R _31263_ (.A1(_02205_),
    .A2(_11431_),
    .B(_11502_),
    .Y(_03983_));
 NAND2x1_ASAP7_75t_R _31264_ (.A(_05244_),
    .B(_06752_),
    .Y(_11503_));
 OA211x2_ASAP7_75t_R _31265_ (.A1(_06541_),
    .A2(_06752_),
    .B(_11503_),
    .C(_05779_),
    .Y(_11504_));
 AOI21x1_ASAP7_75t_R _31266_ (.A1(_02204_),
    .A2(_11431_),
    .B(_11504_),
    .Y(_03984_));
 OR2x2_ASAP7_75t_R _31267_ (.A(_05355_),
    .B(_05944_),
    .Y(_11505_));
 OA211x2_ASAP7_75t_R _31268_ (.A1(_05404_),
    .A2(_06752_),
    .B(_11505_),
    .C(_05779_),
    .Y(_11506_));
 AOI21x1_ASAP7_75t_R _31269_ (.A1(_02203_),
    .A2(_11431_),
    .B(_11506_),
    .Y(_03985_));
 INVx1_ASAP7_75t_R _31270_ (.A(_05943_),
    .Y(_11507_));
 OA211x2_ASAP7_75t_R _31271_ (.A1(net173),
    .A2(_11507_),
    .B(_05779_),
    .C(_05454_),
    .Y(_11508_));
 AO21x1_ASAP7_75t_R _31272_ (.A1(_08745_),
    .A2(_11431_),
    .B(_11508_),
    .Y(_03986_));
 OR3x4_ASAP7_75t_R _31273_ (.A(_06354_),
    .B(net2758),
    .C(_06565_),
    .Y(_11509_));
 TAPCELL_ASAP7_75t_R PHY_225 ();
 TAPCELL_ASAP7_75t_R PHY_224 ();
 TAPCELL_ASAP7_75t_R PHY_223 ();
 NAND2x1_ASAP7_75t_R _31277_ (.A(_02201_),
    .B(_11509_),
    .Y(_11513_));
 OA21x2_ASAP7_75t_R _31278_ (.A1(net239),
    .A2(_11509_),
    .B(_11513_),
    .Y(_03987_));
 NAND2x1_ASAP7_75t_R _31279_ (.A(_02200_),
    .B(_11509_),
    .Y(_11514_));
 OA21x2_ASAP7_75t_R _31280_ (.A1(net242),
    .A2(_11509_),
    .B(_11514_),
    .Y(_03988_));
 NAND2x1_ASAP7_75t_R _31281_ (.A(_02199_),
    .B(_11509_),
    .Y(_11515_));
 OA21x2_ASAP7_75t_R _31282_ (.A1(net243),
    .A2(_11509_),
    .B(_11515_),
    .Y(_03989_));
 NAND2x1_ASAP7_75t_R _31283_ (.A(_02198_),
    .B(_11509_),
    .Y(_11516_));
 OA21x2_ASAP7_75t_R _31284_ (.A1(net244),
    .A2(_11509_),
    .B(_11516_),
    .Y(_03990_));
 NAND2x1_ASAP7_75t_R _31285_ (.A(_02197_),
    .B(_11509_),
    .Y(_11517_));
 OA21x2_ASAP7_75t_R _31286_ (.A1(net245),
    .A2(_11509_),
    .B(_11517_),
    .Y(_03991_));
 NAND2x1_ASAP7_75t_R _31287_ (.A(_02196_),
    .B(_11509_),
    .Y(_11518_));
 OA21x2_ASAP7_75t_R _31288_ (.A1(net246),
    .A2(_11509_),
    .B(_11518_),
    .Y(_03992_));
 NAND2x1_ASAP7_75t_R _31289_ (.A(_02195_),
    .B(_11509_),
    .Y(_11519_));
 OA21x2_ASAP7_75t_R _31290_ (.A1(net247),
    .A2(_11509_),
    .B(_11519_),
    .Y(_03993_));
 NAND2x1_ASAP7_75t_R _31291_ (.A(_02194_),
    .B(_11509_),
    .Y(_11520_));
 OA21x2_ASAP7_75t_R _31292_ (.A1(net248),
    .A2(_11509_),
    .B(_11520_),
    .Y(_03994_));
 NAND2x1_ASAP7_75t_R _31293_ (.A(_02193_),
    .B(_11509_),
    .Y(_11521_));
 OA21x2_ASAP7_75t_R _31294_ (.A1(net219),
    .A2(_11509_),
    .B(_11521_),
    .Y(_03995_));
 NAND2x1_ASAP7_75t_R _31295_ (.A(_02192_),
    .B(_11509_),
    .Y(_11522_));
 OA21x2_ASAP7_75t_R _31296_ (.A1(net220),
    .A2(_11509_),
    .B(_11522_),
    .Y(_03996_));
 TAPCELL_ASAP7_75t_R PHY_222 ();
 TAPCELL_ASAP7_75t_R PHY_221 ();
 NAND2x1_ASAP7_75t_R _31299_ (.A(_02191_),
    .B(_11509_),
    .Y(_11525_));
 OA21x2_ASAP7_75t_R _31300_ (.A1(net221),
    .A2(_11509_),
    .B(_11525_),
    .Y(_03997_));
 NAND2x1_ASAP7_75t_R _31301_ (.A(_02190_),
    .B(_11509_),
    .Y(_11526_));
 OA21x2_ASAP7_75t_R _31302_ (.A1(net222),
    .A2(_11509_),
    .B(_11526_),
    .Y(_03998_));
 NAND2x1_ASAP7_75t_R _31303_ (.A(_02189_),
    .B(_11509_),
    .Y(_11527_));
 OA21x2_ASAP7_75t_R _31304_ (.A1(net223),
    .A2(_11509_),
    .B(_11527_),
    .Y(_03999_));
 NAND2x1_ASAP7_75t_R _31305_ (.A(_02188_),
    .B(_11509_),
    .Y(_11528_));
 OA21x2_ASAP7_75t_R _31306_ (.A1(net224),
    .A2(_11509_),
    .B(_11528_),
    .Y(_04000_));
 NAND2x1_ASAP7_75t_R _31307_ (.A(_02187_),
    .B(_11509_),
    .Y(_11529_));
 OA21x2_ASAP7_75t_R _31308_ (.A1(net225),
    .A2(_11509_),
    .B(_11529_),
    .Y(_04001_));
 NAND2x1_ASAP7_75t_R _31309_ (.A(_02186_),
    .B(_11509_),
    .Y(_11530_));
 OA21x2_ASAP7_75t_R _31310_ (.A1(net226),
    .A2(_11509_),
    .B(_11530_),
    .Y(_04002_));
 NAND2x1_ASAP7_75t_R _31311_ (.A(_02185_),
    .B(_11509_),
    .Y(_11531_));
 OA21x2_ASAP7_75t_R _31312_ (.A1(net227),
    .A2(_11509_),
    .B(_11531_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_R _31313_ (.A(_02184_),
    .B(_11509_),
    .Y(_11532_));
 OA21x2_ASAP7_75t_R _31314_ (.A1(net228),
    .A2(_11509_),
    .B(_11532_),
    .Y(_04004_));
 NAND2x1_ASAP7_75t_R _31315_ (.A(_02183_),
    .B(_11509_),
    .Y(_11533_));
 OA21x2_ASAP7_75t_R _31316_ (.A1(net229),
    .A2(_11509_),
    .B(_11533_),
    .Y(_04005_));
 NAND2x1_ASAP7_75t_R _31317_ (.A(_02182_),
    .B(_11509_),
    .Y(_11534_));
 OA21x2_ASAP7_75t_R _31318_ (.A1(net230),
    .A2(_11509_),
    .B(_11534_),
    .Y(_04006_));
 TAPCELL_ASAP7_75t_R PHY_220 ();
 TAPCELL_ASAP7_75t_R PHY_219 ();
 NAND2x1_ASAP7_75t_R _31321_ (.A(_02181_),
    .B(_11509_),
    .Y(_11537_));
 OA21x2_ASAP7_75t_R _31322_ (.A1(net231),
    .A2(_11509_),
    .B(_11537_),
    .Y(_04007_));
 NAND2x1_ASAP7_75t_R _31323_ (.A(_02180_),
    .B(_11509_),
    .Y(_11538_));
 OA21x2_ASAP7_75t_R _31324_ (.A1(net232),
    .A2(_11509_),
    .B(_11538_),
    .Y(_04008_));
 NAND2x1_ASAP7_75t_R _31325_ (.A(_02179_),
    .B(_11509_),
    .Y(_11539_));
 OA21x2_ASAP7_75t_R _31326_ (.A1(net233),
    .A2(_11509_),
    .B(_11539_),
    .Y(_04009_));
 NAND2x1_ASAP7_75t_R _31327_ (.A(_02178_),
    .B(_11509_),
    .Y(_11540_));
 OA21x2_ASAP7_75t_R _31328_ (.A1(net234),
    .A2(_11509_),
    .B(_11540_),
    .Y(_04010_));
 NAND2x1_ASAP7_75t_R _31329_ (.A(_02177_),
    .B(_11509_),
    .Y(_11541_));
 OA21x2_ASAP7_75t_R _31330_ (.A1(net235),
    .A2(_11509_),
    .B(_11541_),
    .Y(_04011_));
 NAND2x1_ASAP7_75t_R _31331_ (.A(_02176_),
    .B(_11509_),
    .Y(_11542_));
 OA21x2_ASAP7_75t_R _31332_ (.A1(net236),
    .A2(_11509_),
    .B(_11542_),
    .Y(_04012_));
 NAND2x1_ASAP7_75t_R _31333_ (.A(_02175_),
    .B(_11509_),
    .Y(_11543_));
 OA21x2_ASAP7_75t_R _31334_ (.A1(net237),
    .A2(_11509_),
    .B(_11543_),
    .Y(_04013_));
 NAND2x1_ASAP7_75t_R _31335_ (.A(_02174_),
    .B(_11509_),
    .Y(_11544_));
 OA21x2_ASAP7_75t_R _31336_ (.A1(net238),
    .A2(_11509_),
    .B(_11544_),
    .Y(_04014_));
 NAND2x1_ASAP7_75t_R _31337_ (.A(_02173_),
    .B(_11509_),
    .Y(_11545_));
 OA21x2_ASAP7_75t_R _31338_ (.A1(net240),
    .A2(_11509_),
    .B(_11545_),
    .Y(_04015_));
 NAND2x1_ASAP7_75t_R _31339_ (.A(_01729_),
    .B(_11509_),
    .Y(_11546_));
 OA21x2_ASAP7_75t_R _31340_ (.A1(net241),
    .A2(_11509_),
    .B(_11546_),
    .Y(_04016_));
 OA21x2_ASAP7_75t_R _31341_ (.A1(_11103_),
    .A2(_11105_),
    .B(_11122_),
    .Y(_11547_));
 TAPCELL_ASAP7_75t_R PHY_218 ();
 TAPCELL_ASAP7_75t_R PHY_217 ();
 AO21x2_ASAP7_75t_R _31344_ (.A1(_00661_),
    .A2(_11106_),
    .B(_11104_),
    .Y(_11550_));
 TAPCELL_ASAP7_75t_R PHY_216 ();
 OR2x2_ASAP7_75t_R _31346_ (.A(_02488_),
    .B(_11101_),
    .Y(_11552_));
 OA211x2_ASAP7_75t_R _31347_ (.A1(net3517),
    .A2(_11144_),
    .B(_11550_),
    .C(_11552_),
    .Y(_11553_));
 AOI21x1_ASAP7_75t_R _31348_ (.A1(_02172_),
    .A2(_11547_),
    .B(_11553_),
    .Y(_04017_));
 TAPCELL_ASAP7_75t_R PHY_215 ();
 OR3x1_ASAP7_75t_R _31350_ (.A(_02171_),
    .B(_02487_),
    .C(_11101_),
    .Y(_11555_));
 OAI21x1_ASAP7_75t_R _31351_ (.A1(net3647),
    .A2(_11120_),
    .B(_11555_),
    .Y(_11556_));
 TAPCELL_ASAP7_75t_R PHY_214 ();
 AO21x1_ASAP7_75t_R _31353_ (.A1(_02487_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11558_));
 AOI22x1_ASAP7_75t_R _31354_ (.A1(_11550_),
    .A2(_11556_),
    .B1(_11558_),
    .B2(_02171_),
    .Y(_04018_));
 TAPCELL_ASAP7_75t_R PHY_213 ();
 OA211x2_ASAP7_75t_R _31356_ (.A1(_02490_),
    .A2(_11156_),
    .B(_11161_),
    .C(_11550_),
    .Y(_11560_));
 AOI21x1_ASAP7_75t_R _31357_ (.A1(_02170_),
    .A2(_11547_),
    .B(_11560_),
    .Y(_04019_));
 NOR2x1_ASAP7_75t_R _31358_ (.A(_02169_),
    .B(_02489_),
    .Y(_11561_));
 AO21x1_ASAP7_75t_R _31359_ (.A1(_11144_),
    .A2(_11561_),
    .B(_11166_),
    .Y(_11562_));
 AO21x1_ASAP7_75t_R _31360_ (.A1(_02489_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11563_));
 AOI22x1_ASAP7_75t_R _31361_ (.A1(_11550_),
    .A2(_11562_),
    .B1(_11563_),
    .B2(_02169_),
    .Y(_04020_));
 NOR2x1_ASAP7_75t_R _31362_ (.A(_02492_),
    .B(_11156_),
    .Y(_11564_));
 OR3x1_ASAP7_75t_R _31363_ (.A(_11172_),
    .B(_11547_),
    .C(_11564_),
    .Y(_11565_));
 OA21x2_ASAP7_75t_R _31364_ (.A1(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .A2(_11550_),
    .B(_11565_),
    .Y(_04021_));
 NOR2x1_ASAP7_75t_R _31365_ (.A(_02167_),
    .B(_02491_),
    .Y(_11566_));
 AO21x1_ASAP7_75t_R _31366_ (.A1(_11144_),
    .A2(_11566_),
    .B(_11175_),
    .Y(_11567_));
 AO21x1_ASAP7_75t_R _31367_ (.A1(_02491_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11568_));
 AOI22x1_ASAP7_75t_R _31368_ (.A1(_11550_),
    .A2(_11567_),
    .B1(_11568_),
    .B2(_02167_),
    .Y(_04022_));
 OA211x2_ASAP7_75t_R _31369_ (.A1(_02494_),
    .A2(_11156_),
    .B(_11178_),
    .C(_11550_),
    .Y(_11569_));
 AOI21x1_ASAP7_75t_R _31370_ (.A1(_02166_),
    .A2(_11547_),
    .B(_11569_),
    .Y(_04023_));
 NOR2x1_ASAP7_75t_R _31371_ (.A(_02165_),
    .B(_02493_),
    .Y(_11570_));
 AO21x1_ASAP7_75t_R _31372_ (.A1(_11120_),
    .A2(_11570_),
    .B(_11183_),
    .Y(_11571_));
 AO21x1_ASAP7_75t_R _31373_ (.A1(_02493_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11572_));
 AOI22x1_ASAP7_75t_R _31374_ (.A1(_11550_),
    .A2(_11571_),
    .B1(_11572_),
    .B2(_02165_),
    .Y(_04024_));
 OA211x2_ASAP7_75t_R _31375_ (.A1(_02496_),
    .A2(_11156_),
    .B(_11186_),
    .C(_11550_),
    .Y(_11573_));
 AOI21x1_ASAP7_75t_R _31376_ (.A1(_02164_),
    .A2(_11547_),
    .B(_11573_),
    .Y(_04025_));
 NOR2x1_ASAP7_75t_R _31377_ (.A(_02163_),
    .B(_02495_),
    .Y(_11574_));
 AO21x1_ASAP7_75t_R _31378_ (.A1(_11144_),
    .A2(_11574_),
    .B(_11189_),
    .Y(_11575_));
 AO21x1_ASAP7_75t_R _31379_ (.A1(_02495_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11576_));
 AOI22x1_ASAP7_75t_R _31380_ (.A1(_11550_),
    .A2(_11575_),
    .B1(_11576_),
    .B2(_02163_),
    .Y(_04026_));
 OA211x2_ASAP7_75t_R _31381_ (.A1(_02498_),
    .A2(_11156_),
    .B(_11192_),
    .C(_11550_),
    .Y(_11577_));
 AOI21x1_ASAP7_75t_R _31382_ (.A1(_02162_),
    .A2(_11547_),
    .B(_11577_),
    .Y(_04027_));
 NOR2x1_ASAP7_75t_R _31383_ (.A(_02161_),
    .B(_02497_),
    .Y(_11578_));
 AO21x1_ASAP7_75t_R _31384_ (.A1(_11144_),
    .A2(_11578_),
    .B(_11195_),
    .Y(_11579_));
 AO21x1_ASAP7_75t_R _31385_ (.A1(_02497_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11580_));
 AOI22x1_ASAP7_75t_R _31386_ (.A1(_11550_),
    .A2(_11579_),
    .B1(_11580_),
    .B2(_02161_),
    .Y(_04028_));
 OA211x2_ASAP7_75t_R _31387_ (.A1(_02500_),
    .A2(_11198_),
    .B(_11200_),
    .C(_11550_),
    .Y(_11581_));
 AOI21x1_ASAP7_75t_R _31388_ (.A1(_02160_),
    .A2(_11547_),
    .B(_11581_),
    .Y(_04029_));
 NOR2x1_ASAP7_75t_R _31389_ (.A(_02159_),
    .B(_02499_),
    .Y(_11582_));
 AO21x1_ASAP7_75t_R _31390_ (.A1(_11120_),
    .A2(_11582_),
    .B(_11203_),
    .Y(_11583_));
 AO21x1_ASAP7_75t_R _31391_ (.A1(_02499_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11584_));
 AOI22x1_ASAP7_75t_R _31392_ (.A1(_11550_),
    .A2(_11583_),
    .B1(_11584_),
    .B2(_02159_),
    .Y(_04030_));
 OA211x2_ASAP7_75t_R _31393_ (.A1(_02502_),
    .A2(_11156_),
    .B(_11206_),
    .C(_11550_),
    .Y(_11585_));
 AOI21x1_ASAP7_75t_R _31394_ (.A1(_02158_),
    .A2(_11547_),
    .B(_11585_),
    .Y(_04031_));
 NOR2x1_ASAP7_75t_R _31395_ (.A(_02157_),
    .B(_02501_),
    .Y(_11586_));
 AO21x1_ASAP7_75t_R _31396_ (.A1(_11120_),
    .A2(_11586_),
    .B(_11209_),
    .Y(_11587_));
 AO21x1_ASAP7_75t_R _31397_ (.A1(_02501_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11588_));
 AOI22x1_ASAP7_75t_R _31398_ (.A1(_11550_),
    .A2(_11587_),
    .B1(_11588_),
    .B2(_02157_),
    .Y(_04032_));
 NOR2x1_ASAP7_75t_R _31399_ (.A(_02504_),
    .B(_11156_),
    .Y(_11589_));
 OR3x1_ASAP7_75t_R _31400_ (.A(_11213_),
    .B(_11547_),
    .C(_11589_),
    .Y(_11590_));
 OA21x2_ASAP7_75t_R _31401_ (.A1(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .A2(_11550_),
    .B(_11590_),
    .Y(_04033_));
 OR4x1_ASAP7_75t_R _31402_ (.A(_02155_),
    .B(_02503_),
    .C(_11107_),
    .D(_11156_),
    .Y(_11591_));
 AO21x1_ASAP7_75t_R _31403_ (.A1(_02503_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11592_));
 NAND2x1_ASAP7_75t_R _31404_ (.A(_02155_),
    .B(_11592_),
    .Y(_11593_));
 OA211x2_ASAP7_75t_R _31405_ (.A1(net3660),
    .A2(_11122_),
    .B(_11591_),
    .C(_11593_),
    .Y(_04034_));
 OA211x2_ASAP7_75t_R _31406_ (.A1(_02506_),
    .A2(_11198_),
    .B(_11550_),
    .C(_11220_),
    .Y(_11594_));
 AOI21x1_ASAP7_75t_R _31407_ (.A1(_02154_),
    .A2(_11547_),
    .B(_11594_),
    .Y(_04035_));
 NOR2x1_ASAP7_75t_R _31408_ (.A(_02153_),
    .B(_02505_),
    .Y(_11595_));
 AO21x1_ASAP7_75t_R _31409_ (.A1(_11144_),
    .A2(_11595_),
    .B(_11223_),
    .Y(_11596_));
 AO21x1_ASAP7_75t_R _31410_ (.A1(_02505_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11597_));
 AOI22x1_ASAP7_75t_R _31411_ (.A1(_11550_),
    .A2(_11596_),
    .B1(_11597_),
    .B2(_02153_),
    .Y(_04036_));
 OA211x2_ASAP7_75t_R _31412_ (.A1(_02508_),
    .A2(_11198_),
    .B(_11550_),
    .C(_11226_),
    .Y(_11598_));
 AOI21x1_ASAP7_75t_R _31413_ (.A1(_02152_),
    .A2(_11547_),
    .B(_11598_),
    .Y(_04037_));
 AO21x1_ASAP7_75t_R _31414_ (.A1(_02507_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11599_));
 NAND2x1_ASAP7_75t_R _31415_ (.A(_02151_),
    .B(_11599_),
    .Y(_11600_));
 OR4x1_ASAP7_75t_R _31416_ (.A(_02151_),
    .B(_02507_),
    .C(_11198_),
    .D(_11547_),
    .Y(_11601_));
 OA211x2_ASAP7_75t_R _31417_ (.A1(_09623_),
    .A2(_11122_),
    .B(_11600_),
    .C(_11601_),
    .Y(_04038_));
 OA211x2_ASAP7_75t_R _31418_ (.A1(_02510_),
    .A2(_11198_),
    .B(_11550_),
    .C(_11231_),
    .Y(_11602_));
 AOI21x1_ASAP7_75t_R _31419_ (.A1(_02150_),
    .A2(_11547_),
    .B(_11602_),
    .Y(_04039_));
 NOR2x1_ASAP7_75t_R _31420_ (.A(_02149_),
    .B(_02509_),
    .Y(_11603_));
 AO21x1_ASAP7_75t_R _31421_ (.A1(_11120_),
    .A2(_11603_),
    .B(_11234_),
    .Y(_11604_));
 AO21x1_ASAP7_75t_R _31422_ (.A1(_02509_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11605_));
 AOI22x1_ASAP7_75t_R _31423_ (.A1(_11550_),
    .A2(_11604_),
    .B1(_11605_),
    .B2(_02149_),
    .Y(_04040_));
 OR2x2_ASAP7_75t_R _31424_ (.A(_02512_),
    .B(_11156_),
    .Y(_11606_));
 OA211x2_ASAP7_75t_R _31425_ (.A1(_11237_),
    .A2(_11120_),
    .B(_11550_),
    .C(_11606_),
    .Y(_11607_));
 AOI21x1_ASAP7_75t_R _31426_ (.A1(_02148_),
    .A2(_11547_),
    .B(_11607_),
    .Y(_04041_));
 NOR2x1_ASAP7_75t_R _31427_ (.A(_02147_),
    .B(_02511_),
    .Y(_11608_));
 AO21x1_ASAP7_75t_R _31428_ (.A1(_11144_),
    .A2(_11608_),
    .B(_11241_),
    .Y(_11609_));
 AO21x1_ASAP7_75t_R _31429_ (.A1(_02511_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11610_));
 AOI22x1_ASAP7_75t_R _31430_ (.A1(_11550_),
    .A2(_11609_),
    .B1(_11610_),
    .B2(_02147_),
    .Y(_04042_));
 OA211x2_ASAP7_75t_R _31431_ (.A1(_02514_),
    .A2(_11156_),
    .B(_11550_),
    .C(_11244_),
    .Y(_11611_));
 AOI21x1_ASAP7_75t_R _31432_ (.A1(_02146_),
    .A2(_11547_),
    .B(_11611_),
    .Y(_04043_));
 NOR2x1_ASAP7_75t_R _31433_ (.A(_02145_),
    .B(_02513_),
    .Y(_11612_));
 AO21x1_ASAP7_75t_R _31434_ (.A1(_11120_),
    .A2(_11612_),
    .B(_11247_),
    .Y(_11613_));
 AO21x1_ASAP7_75t_R _31435_ (.A1(_02513_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11614_));
 AOI22x1_ASAP7_75t_R _31436_ (.A1(_11550_),
    .A2(_11613_),
    .B1(_11614_),
    .B2(_02145_),
    .Y(_04044_));
 OA211x2_ASAP7_75t_R _31437_ (.A1(_02516_),
    .A2(_11198_),
    .B(_11550_),
    .C(_11251_),
    .Y(_11615_));
 AOI21x1_ASAP7_75t_R _31438_ (.A1(_02144_),
    .A2(_11547_),
    .B(_11615_),
    .Y(_04045_));
 NOR2x1_ASAP7_75t_R _31439_ (.A(_02143_),
    .B(_02515_),
    .Y(_11616_));
 AO21x1_ASAP7_75t_R _31440_ (.A1(_11120_),
    .A2(_11616_),
    .B(_11254_),
    .Y(_11617_));
 AO21x1_ASAP7_75t_R _31441_ (.A1(_02515_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11618_));
 AOI22x1_ASAP7_75t_R _31442_ (.A1(_11550_),
    .A2(_11617_),
    .B1(_11618_),
    .B2(_02143_),
    .Y(_04046_));
 OA211x2_ASAP7_75t_R _31443_ (.A1(_02518_),
    .A2(_11156_),
    .B(_11550_),
    .C(_11257_),
    .Y(_11619_));
 AOI21x1_ASAP7_75t_R _31444_ (.A1(_02142_),
    .A2(_11547_),
    .B(_11619_),
    .Y(_04047_));
 AO21x1_ASAP7_75t_R _31445_ (.A1(_02517_),
    .A2(_11144_),
    .B(_11547_),
    .Y(_11620_));
 NAND2x1_ASAP7_75t_R _31446_ (.A(_02141_),
    .B(_11620_),
    .Y(_11621_));
 OR4x1_ASAP7_75t_R _31447_ (.A(_02141_),
    .B(_02517_),
    .C(_11101_),
    .D(_11547_),
    .Y(_11622_));
 OA211x2_ASAP7_75t_R _31448_ (.A1(_09698_),
    .A2(_11122_),
    .B(_11621_),
    .C(_11622_),
    .Y(_04048_));
 TAPCELL_ASAP7_75t_R PHY_212 ();
 AOI21x1_ASAP7_75t_R _31450_ (.A1(_05727_),
    .A2(_05728_),
    .B(_06300_),
    .Y(_11624_));
 AND2x2_ASAP7_75t_R _31451_ (.A(_01456_),
    .B(_06420_),
    .Y(_11625_));
 AO21x1_ASAP7_75t_R _31452_ (.A1(_01577_),
    .A2(_06366_),
    .B(_11625_),
    .Y(_11626_));
 AO21x1_ASAP7_75t_R _31453_ (.A1(_05727_),
    .A2(_05728_),
    .B(_06300_),
    .Y(_11627_));
 AND2x2_ASAP7_75t_R _31454_ (.A(_02140_),
    .B(_11627_),
    .Y(_11628_));
 AO21x1_ASAP7_75t_R _31455_ (.A1(_11624_),
    .A2(_11626_),
    .B(_11628_),
    .Y(_11629_));
 NAND2x1_ASAP7_75t_R _31456_ (.A(_11406_),
    .B(_11629_),
    .Y(_04049_));
 AND2x2_ASAP7_75t_R _31457_ (.A(_01455_),
    .B(_06420_),
    .Y(_11630_));
 AO21x1_ASAP7_75t_R _31458_ (.A1(_01576_),
    .A2(_06366_),
    .B(_11630_),
    .Y(_11631_));
 AND2x2_ASAP7_75t_R _31459_ (.A(_17810_),
    .B(_11627_),
    .Y(_11632_));
 AO21x1_ASAP7_75t_R _31460_ (.A1(_11624_),
    .A2(_11631_),
    .B(_11632_),
    .Y(_11633_));
 NAND2x1_ASAP7_75t_R _31461_ (.A(_11406_),
    .B(_11633_),
    .Y(_04050_));
 NAND3x2_ASAP7_75t_R _31462_ (.B(_11086_),
    .C(_11096_),
    .Y(_11634_),
    .A(_05693_));
 TAPCELL_ASAP7_75t_R PHY_211 ();
 TAPCELL_ASAP7_75t_R PHY_210 ();
 NAND2x1_ASAP7_75t_R _31465_ (.A(_02139_),
    .B(_11634_),
    .Y(_11637_));
 OA21x2_ASAP7_75t_R _31466_ (.A1(_11262_),
    .A2(_11634_),
    .B(_11637_),
    .Y(_04051_));
 NAND2x1_ASAP7_75t_R _31467_ (.A(_02138_),
    .B(_11634_),
    .Y(_11638_));
 OA21x2_ASAP7_75t_R _31468_ (.A1(net3647),
    .A2(_11634_),
    .B(_11638_),
    .Y(_04052_));
 NAND2x1_ASAP7_75t_R _31469_ (.A(_02137_),
    .B(_11634_),
    .Y(_11639_));
 OA21x2_ASAP7_75t_R _31470_ (.A1(_11159_),
    .A2(_11634_),
    .B(_11639_),
    .Y(_04053_));
 NAND2x1_ASAP7_75t_R _31471_ (.A(_02136_),
    .B(_11634_),
    .Y(_11640_));
 OA21x2_ASAP7_75t_R _31472_ (.A1(net3544),
    .A2(_11634_),
    .B(_11640_),
    .Y(_04054_));
 NAND2x1_ASAP7_75t_R _31473_ (.A(_02135_),
    .B(_11634_),
    .Y(_11641_));
 OA21x2_ASAP7_75t_R _31474_ (.A1(net3379),
    .A2(_11634_),
    .B(_11641_),
    .Y(_04055_));
 NAND2x1_ASAP7_75t_R _31475_ (.A(_02134_),
    .B(_11634_),
    .Y(_11642_));
 OA21x2_ASAP7_75t_R _31476_ (.A1(net3632),
    .A2(_11634_),
    .B(_11642_),
    .Y(_04056_));
 NAND2x1_ASAP7_75t_R _31477_ (.A(_02133_),
    .B(_11634_),
    .Y(_11643_));
 OA21x2_ASAP7_75t_R _31478_ (.A1(_09504_),
    .A2(_11634_),
    .B(_11643_),
    .Y(_04057_));
 NAND2x1_ASAP7_75t_R _31479_ (.A(_02132_),
    .B(_11634_),
    .Y(_11644_));
 OA21x2_ASAP7_75t_R _31480_ (.A1(net3654),
    .A2(_11634_),
    .B(_11644_),
    .Y(_04058_));
 NAND2x1_ASAP7_75t_R _31481_ (.A(_02131_),
    .B(_11634_),
    .Y(_11645_));
 OA21x2_ASAP7_75t_R _31482_ (.A1(net3725),
    .A2(_11634_),
    .B(_11645_),
    .Y(_04059_));
 TAPCELL_ASAP7_75t_R PHY_209 ();
 NAND2x1_ASAP7_75t_R _31484_ (.A(_02130_),
    .B(_11634_),
    .Y(_11647_));
 OA21x2_ASAP7_75t_R _31485_ (.A1(net3716),
    .A2(_11634_),
    .B(_11647_),
    .Y(_04060_));
 TAPCELL_ASAP7_75t_R PHY_208 ();
 NAND2x1_ASAP7_75t_R _31487_ (.A(_02129_),
    .B(_11634_),
    .Y(_11649_));
 OA21x2_ASAP7_75t_R _31488_ (.A1(net3736),
    .A2(_11634_),
    .B(_11649_),
    .Y(_04061_));
 NAND2x1_ASAP7_75t_R _31489_ (.A(_02128_),
    .B(_11634_),
    .Y(_11650_));
 OA21x2_ASAP7_75t_R _31490_ (.A1(_09538_),
    .A2(_11634_),
    .B(_11650_),
    .Y(_04062_));
 NAND2x1_ASAP7_75t_R _31491_ (.A(_02127_),
    .B(_11634_),
    .Y(_11651_));
 OA21x2_ASAP7_75t_R _31492_ (.A1(net3673),
    .A2(_11634_),
    .B(_11651_),
    .Y(_04063_));
 NAND2x1_ASAP7_75t_R _31493_ (.A(_02126_),
    .B(_11634_),
    .Y(_11652_));
 OA21x2_ASAP7_75t_R _31494_ (.A1(net3707),
    .A2(_11634_),
    .B(_11652_),
    .Y(_04064_));
 NAND2x1_ASAP7_75t_R _31495_ (.A(_02125_),
    .B(_11634_),
    .Y(_11653_));
 OA21x2_ASAP7_75t_R _31496_ (.A1(net3541),
    .A2(_11634_),
    .B(_11653_),
    .Y(_04065_));
 NAND2x1_ASAP7_75t_R _31497_ (.A(_02124_),
    .B(_11634_),
    .Y(_11654_));
 OA21x2_ASAP7_75t_R _31498_ (.A1(net3747),
    .A2(_11634_),
    .B(_11654_),
    .Y(_04066_));
 NAND2x1_ASAP7_75t_R _31499_ (.A(_02123_),
    .B(_11634_),
    .Y(_11655_));
 OA21x2_ASAP7_75t_R _31500_ (.A1(net3604),
    .A2(_11634_),
    .B(_11655_),
    .Y(_04067_));
 NAND2x1_ASAP7_75t_R _31501_ (.A(_02122_),
    .B(_11634_),
    .Y(_11656_));
 OA21x2_ASAP7_75t_R _31502_ (.A1(net3660),
    .A2(_11634_),
    .B(_11656_),
    .Y(_04068_));
 NAND2x1_ASAP7_75t_R _31503_ (.A(_02121_),
    .B(_11634_),
    .Y(_11657_));
 OA21x2_ASAP7_75t_R _31504_ (.A1(net3557),
    .A2(_11634_),
    .B(_11657_),
    .Y(_04069_));
 TAPCELL_ASAP7_75t_R PHY_207 ();
 NAND2x1_ASAP7_75t_R _31506_ (.A(_02120_),
    .B(_11634_),
    .Y(_11659_));
 OA21x2_ASAP7_75t_R _31507_ (.A1(net3721),
    .A2(_11634_),
    .B(_11659_),
    .Y(_04070_));
 TAPCELL_ASAP7_75t_R PHY_206 ();
 NAND2x1_ASAP7_75t_R _31509_ (.A(_02119_),
    .B(_11634_),
    .Y(_11661_));
 OA21x2_ASAP7_75t_R _31510_ (.A1(net3683),
    .A2(_11634_),
    .B(_11661_),
    .Y(_04071_));
 NAND2x1_ASAP7_75t_R _31511_ (.A(_02118_),
    .B(_11634_),
    .Y(_11662_));
 OA21x2_ASAP7_75t_R _31512_ (.A1(_09623_),
    .A2(_11634_),
    .B(_11662_),
    .Y(_04072_));
 NAND2x1_ASAP7_75t_R _31513_ (.A(_02117_),
    .B(_11634_),
    .Y(_11663_));
 OA21x2_ASAP7_75t_R _31514_ (.A1(net3691),
    .A2(_11634_),
    .B(_11663_),
    .Y(_04073_));
 NAND2x1_ASAP7_75t_R _31515_ (.A(_02116_),
    .B(_11634_),
    .Y(_11664_));
 OA21x2_ASAP7_75t_R _31516_ (.A1(_09638_),
    .A2(_11634_),
    .B(_11664_),
    .Y(_04074_));
 NAND2x1_ASAP7_75t_R _31517_ (.A(_08437_),
    .B(_11634_),
    .Y(_11665_));
 OR3x1_ASAP7_75t_R _31518_ (.A(net3531),
    .B(_09646_),
    .C(_11634_),
    .Y(_11666_));
 NAND2x1_ASAP7_75t_R _31519_ (.A(_11665_),
    .B(_11666_),
    .Y(_04075_));
 NAND2x1_ASAP7_75t_R _31520_ (.A(_02114_),
    .B(_11634_),
    .Y(_11667_));
 OA21x2_ASAP7_75t_R _31521_ (.A1(net3639),
    .A2(_11634_),
    .B(_11667_),
    .Y(_04076_));
 NAND2x1_ASAP7_75t_R _31522_ (.A(_02113_),
    .B(_11634_),
    .Y(_11668_));
 OA21x2_ASAP7_75t_R _31523_ (.A1(_09662_),
    .A2(_11634_),
    .B(_11668_),
    .Y(_04077_));
 NAND2x1_ASAP7_75t_R _31524_ (.A(_02112_),
    .B(_11634_),
    .Y(_11669_));
 OA21x2_ASAP7_75t_R _31525_ (.A1(net3594),
    .A2(_11634_),
    .B(_11669_),
    .Y(_04078_));
 NAND2x1_ASAP7_75t_R _31526_ (.A(_02111_),
    .B(_11634_),
    .Y(_11670_));
 OA21x2_ASAP7_75t_R _31527_ (.A1(_09676_),
    .A2(_11634_),
    .B(_11670_),
    .Y(_04079_));
 NAND2x1_ASAP7_75t_R _31528_ (.A(_02110_),
    .B(_11634_),
    .Y(_11671_));
 OA21x2_ASAP7_75t_R _31529_ (.A1(net3611),
    .A2(_11634_),
    .B(_11671_),
    .Y(_04080_));
 NAND2x1_ASAP7_75t_R _31530_ (.A(_02109_),
    .B(_11634_),
    .Y(_11672_));
 OA21x2_ASAP7_75t_R _31531_ (.A1(net3698),
    .A2(_11634_),
    .B(_11672_),
    .Y(_04081_));
 NAND2x1_ASAP7_75t_R _31532_ (.A(_02108_),
    .B(_11634_),
    .Y(_11673_));
 OA21x2_ASAP7_75t_R _31533_ (.A1(_09698_),
    .A2(_11634_),
    .B(_11673_),
    .Y(_04082_));
 TAPCELL_ASAP7_75t_R PHY_205 ();
 NOR2x2_ASAP7_75t_R _31535_ (.A(_11406_),
    .B(_11407_),
    .Y(_11675_));
 TAPCELL_ASAP7_75t_R PHY_204 ();
 TAPCELL_ASAP7_75t_R PHY_203 ();
 AND2x2_ASAP7_75t_R _31538_ (.A(_01456_),
    .B(_11675_),
    .Y(_11678_));
 AOI21x1_ASAP7_75t_R _31539_ (.A1(_02107_),
    .A2(_11408_),
    .B(_11678_),
    .Y(_04083_));
 TAPCELL_ASAP7_75t_R PHY_202 ();
 NAND2x1_ASAP7_75t_R _31541_ (.A(_02106_),
    .B(_11408_),
    .Y(_11680_));
 OA21x2_ASAP7_75t_R _31542_ (.A1(_11417_),
    .A2(_11408_),
    .B(_11680_),
    .Y(_04084_));
 AND2x2_ASAP7_75t_R _31543_ (.A(_01454_),
    .B(_11675_),
    .Y(_11681_));
 AOI21x1_ASAP7_75t_R _31544_ (.A1(_02105_),
    .A2(_11408_),
    .B(_11681_),
    .Y(_04085_));
 AND2x2_ASAP7_75t_R _31545_ (.A(_01913_),
    .B(_11675_),
    .Y(_11682_));
 AOI21x1_ASAP7_75t_R _31546_ (.A1(_02104_),
    .A2(_11408_),
    .B(_11682_),
    .Y(_04086_));
 INVx1_ASAP7_75t_R _31547_ (.A(_02103_),
    .Y(_11683_));
 TAPCELL_ASAP7_75t_R PHY_201 ();
 TAPCELL_ASAP7_75t_R PHY_200 ();
 TAPCELL_ASAP7_75t_R PHY_199 ();
 NAND2x1_ASAP7_75t_R _31551_ (.A(_01912_),
    .B(_11675_),
    .Y(_11687_));
 OA21x2_ASAP7_75t_R _31552_ (.A1(_11683_),
    .A2(_11675_),
    .B(_11687_),
    .Y(_04087_));
 AND2x2_ASAP7_75t_R _31553_ (.A(_01911_),
    .B(_11675_),
    .Y(_11688_));
 AOI21x1_ASAP7_75t_R _31554_ (.A1(_02102_),
    .A2(_11408_),
    .B(_11688_),
    .Y(_04088_));
 INVx1_ASAP7_75t_R _31555_ (.A(_01910_),
    .Y(_11689_));
 NAND2x1_ASAP7_75t_R _31556_ (.A(_02101_),
    .B(_11408_),
    .Y(_11690_));
 OA21x2_ASAP7_75t_R _31557_ (.A1(_11689_),
    .A2(_11408_),
    .B(_11690_),
    .Y(_04089_));
 AND2x2_ASAP7_75t_R _31558_ (.A(_01909_),
    .B(_11675_),
    .Y(_11691_));
 AOI21x1_ASAP7_75t_R _31559_ (.A1(_02100_),
    .A2(_11408_),
    .B(_11691_),
    .Y(_04090_));
 AND2x2_ASAP7_75t_R _31560_ (.A(_01908_),
    .B(_11675_),
    .Y(_11692_));
 AOI21x1_ASAP7_75t_R _31561_ (.A1(_02099_),
    .A2(_11408_),
    .B(_11692_),
    .Y(_04091_));
 AND4x1_ASAP7_75t_R _31562_ (.A(_13525_),
    .B(_05564_),
    .C(_05702_),
    .D(_11087_),
    .Y(_11693_));
 NAND2x2_ASAP7_75t_R _31563_ (.A(_11693_),
    .B(_11096_),
    .Y(_11694_));
 TAPCELL_ASAP7_75t_R PHY_198 ();
 TAPCELL_ASAP7_75t_R PHY_197 ();
 NAND2x1_ASAP7_75t_R _31566_ (.A(_02098_),
    .B(_11694_),
    .Y(_11697_));
 OA21x2_ASAP7_75t_R _31567_ (.A1(_11262_),
    .A2(_11694_),
    .B(_11697_),
    .Y(_04092_));
 NAND2x1_ASAP7_75t_R _31568_ (.A(_02097_),
    .B(_11694_),
    .Y(_11698_));
 OA21x2_ASAP7_75t_R _31569_ (.A1(net3647),
    .A2(_11694_),
    .B(_11698_),
    .Y(_04093_));
 NAND2x1_ASAP7_75t_R _31570_ (.A(_02096_),
    .B(_11694_),
    .Y(_11699_));
 OA21x2_ASAP7_75t_R _31571_ (.A1(_11159_),
    .A2(_11694_),
    .B(_11699_),
    .Y(_04094_));
 NAND2x1_ASAP7_75t_R _31572_ (.A(_02095_),
    .B(_11694_),
    .Y(_11700_));
 OA21x2_ASAP7_75t_R _31573_ (.A1(net3544),
    .A2(_11694_),
    .B(_11700_),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_R _31574_ (.A(_02094_),
    .B(_11694_),
    .Y(_11701_));
 OA21x2_ASAP7_75t_R _31575_ (.A1(net3379),
    .A2(_11694_),
    .B(_11701_),
    .Y(_04096_));
 NAND2x1_ASAP7_75t_R _31576_ (.A(_02093_),
    .B(_11694_),
    .Y(_11702_));
 OA21x2_ASAP7_75t_R _31577_ (.A1(net3632),
    .A2(_11694_),
    .B(_11702_),
    .Y(_04097_));
 NAND2x1_ASAP7_75t_R _31578_ (.A(_02092_),
    .B(_11694_),
    .Y(_11703_));
 OA21x2_ASAP7_75t_R _31579_ (.A1(_09504_),
    .A2(_11694_),
    .B(_11703_),
    .Y(_04098_));
 NAND2x1_ASAP7_75t_R _31580_ (.A(_02091_),
    .B(_11694_),
    .Y(_11704_));
 OA21x2_ASAP7_75t_R _31581_ (.A1(net3654),
    .A2(_11694_),
    .B(_11704_),
    .Y(_04099_));
 NAND2x1_ASAP7_75t_R _31582_ (.A(_02090_),
    .B(_11694_),
    .Y(_11705_));
 OA21x2_ASAP7_75t_R _31583_ (.A1(net3725),
    .A2(_11694_),
    .B(_11705_),
    .Y(_04100_));
 TAPCELL_ASAP7_75t_R PHY_196 ();
 NAND2x1_ASAP7_75t_R _31585_ (.A(_02089_),
    .B(_11694_),
    .Y(_11707_));
 OA21x2_ASAP7_75t_R _31586_ (.A1(net3716),
    .A2(_11694_),
    .B(_11707_),
    .Y(_04101_));
 TAPCELL_ASAP7_75t_R PHY_195 ();
 NAND2x1_ASAP7_75t_R _31588_ (.A(_02088_),
    .B(_11694_),
    .Y(_11709_));
 OA21x2_ASAP7_75t_R _31589_ (.A1(net3736),
    .A2(_11694_),
    .B(_11709_),
    .Y(_04102_));
 NAND2x1_ASAP7_75t_R _31590_ (.A(_02087_),
    .B(_11694_),
    .Y(_11710_));
 OA21x2_ASAP7_75t_R _31591_ (.A1(_09538_),
    .A2(_11694_),
    .B(_11710_),
    .Y(_04103_));
 NAND2x1_ASAP7_75t_R _31592_ (.A(_02086_),
    .B(_11694_),
    .Y(_11711_));
 OA21x2_ASAP7_75t_R _31593_ (.A1(net3673),
    .A2(_11694_),
    .B(_11711_),
    .Y(_04104_));
 NAND2x1_ASAP7_75t_R _31594_ (.A(_02085_),
    .B(_11694_),
    .Y(_11712_));
 OA21x2_ASAP7_75t_R _31595_ (.A1(net3707),
    .A2(_11694_),
    .B(_11712_),
    .Y(_04105_));
 NAND2x1_ASAP7_75t_R _31596_ (.A(_02084_),
    .B(_11694_),
    .Y(_11713_));
 OA21x2_ASAP7_75t_R _31597_ (.A1(net3541),
    .A2(_11694_),
    .B(_11713_),
    .Y(_04106_));
 NAND2x1_ASAP7_75t_R _31598_ (.A(_02083_),
    .B(_11694_),
    .Y(_11714_));
 OA21x2_ASAP7_75t_R _31599_ (.A1(net3747),
    .A2(_11694_),
    .B(_11714_),
    .Y(_04107_));
 NAND2x1_ASAP7_75t_R _31600_ (.A(_02082_),
    .B(_11694_),
    .Y(_11715_));
 OA21x2_ASAP7_75t_R _31601_ (.A1(net3604),
    .A2(_11694_),
    .B(_11715_),
    .Y(_04108_));
 NAND2x1_ASAP7_75t_R _31602_ (.A(_02081_),
    .B(_11694_),
    .Y(_11716_));
 OA21x2_ASAP7_75t_R _31603_ (.A1(net3660),
    .A2(_11694_),
    .B(_11716_),
    .Y(_04109_));
 NAND2x1_ASAP7_75t_R _31604_ (.A(_02080_),
    .B(_11694_),
    .Y(_11717_));
 OA21x2_ASAP7_75t_R _31605_ (.A1(net3557),
    .A2(_11694_),
    .B(_11717_),
    .Y(_04110_));
 TAPCELL_ASAP7_75t_R PHY_194 ();
 NAND2x1_ASAP7_75t_R _31607_ (.A(_02079_),
    .B(_11694_),
    .Y(_11719_));
 OA21x2_ASAP7_75t_R _31608_ (.A1(net3711),
    .A2(_11694_),
    .B(_11719_),
    .Y(_04111_));
 TAPCELL_ASAP7_75t_R PHY_193 ();
 NAND2x1_ASAP7_75t_R _31610_ (.A(_02078_),
    .B(_11694_),
    .Y(_11721_));
 OA21x2_ASAP7_75t_R _31611_ (.A1(_09616_),
    .A2(_11694_),
    .B(_11721_),
    .Y(_04112_));
 NAND2x1_ASAP7_75t_R _31612_ (.A(_02077_),
    .B(_11694_),
    .Y(_11722_));
 OA21x2_ASAP7_75t_R _31613_ (.A1(_09623_),
    .A2(_11694_),
    .B(_11722_),
    .Y(_04113_));
 NAND2x1_ASAP7_75t_R _31614_ (.A(_02076_),
    .B(_11694_),
    .Y(_11723_));
 OA21x2_ASAP7_75t_R _31615_ (.A1(net3691),
    .A2(_11694_),
    .B(_11723_),
    .Y(_04114_));
 NAND2x1_ASAP7_75t_R _31616_ (.A(_02075_),
    .B(_11694_),
    .Y(_11724_));
 OA21x2_ASAP7_75t_R _31617_ (.A1(_09638_),
    .A2(_11694_),
    .B(_11724_),
    .Y(_04115_));
 NOR2x1_ASAP7_75t_R _31618_ (.A(_07026_),
    .B(_11119_),
    .Y(_11725_));
 NOR2x1_ASAP7_75t_R _31619_ (.A(_02074_),
    .B(_11725_),
    .Y(_11726_));
 AO21x1_ASAP7_75t_R _31620_ (.A1(_09647_),
    .A2(_11725_),
    .B(_11726_),
    .Y(_04116_));
 NAND2x1_ASAP7_75t_R _31621_ (.A(_02073_),
    .B(_11694_),
    .Y(_11727_));
 OA21x2_ASAP7_75t_R _31622_ (.A1(net3644),
    .A2(_11694_),
    .B(_11727_),
    .Y(_04117_));
 NAND2x1_ASAP7_75t_R _31623_ (.A(_02072_),
    .B(_11694_),
    .Y(_11728_));
 OA21x2_ASAP7_75t_R _31624_ (.A1(_09662_),
    .A2(_11694_),
    .B(_11728_),
    .Y(_04118_));
 NAND2x1_ASAP7_75t_R _31625_ (.A(_02071_),
    .B(_11694_),
    .Y(_11729_));
 OA21x2_ASAP7_75t_R _31626_ (.A1(net3594),
    .A2(_11694_),
    .B(_11729_),
    .Y(_04119_));
 NAND2x1_ASAP7_75t_R _31627_ (.A(_02070_),
    .B(_11694_),
    .Y(_11730_));
 OA21x2_ASAP7_75t_R _31628_ (.A1(_09676_),
    .A2(_11694_),
    .B(_11730_),
    .Y(_04120_));
 NAND2x1_ASAP7_75t_R _31629_ (.A(_02069_),
    .B(_11694_),
    .Y(_11731_));
 OA21x2_ASAP7_75t_R _31630_ (.A1(net3611),
    .A2(_11694_),
    .B(_11731_),
    .Y(_04121_));
 NAND2x1_ASAP7_75t_R _31631_ (.A(_02068_),
    .B(_11694_),
    .Y(_11732_));
 OA21x2_ASAP7_75t_R _31632_ (.A1(_09691_),
    .A2(_11694_),
    .B(_11732_),
    .Y(_04122_));
 NAND2x1_ASAP7_75t_R _31633_ (.A(_02067_),
    .B(_11694_),
    .Y(_11733_));
 OA21x2_ASAP7_75t_R _31634_ (.A1(_09698_),
    .A2(_11694_),
    .B(_11733_),
    .Y(_04123_));
 NOR2x2_ASAP7_75t_R _31635_ (.A(_07008_),
    .B(_09445_),
    .Y(_11734_));
 TAPCELL_ASAP7_75t_R PHY_192 ();
 AND3x4_ASAP7_75t_R _31637_ (.A(_01714_),
    .B(_01715_),
    .C(_01716_),
    .Y(_11736_));
 TAPCELL_ASAP7_75t_R PHY_191 ();
 NOR2x2_ASAP7_75t_R _31639_ (.A(_11736_),
    .B(_11734_),
    .Y(_11738_));
 TAPCELL_ASAP7_75t_R PHY_190 ();
 INVx1_ASAP7_75t_R _31641_ (.A(_00095_),
    .Y(_11740_));
 AO22x1_ASAP7_75t_R _31642_ (.A1(net3422),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11740_),
    .Y(_11741_));
 AO21x1_ASAP7_75t_R _31643_ (.A1(net3725),
    .A2(_11734_),
    .B(_11741_),
    .Y(_04124_));
 INVx1_ASAP7_75t_R _31644_ (.A(_00098_),
    .Y(_11742_));
 AO22x1_ASAP7_75t_R _31645_ (.A1(net3126),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11742_),
    .Y(_11743_));
 AO21x1_ASAP7_75t_R _31646_ (.A1(net3716),
    .A2(_11734_),
    .B(_11743_),
    .Y(_04125_));
 INVx1_ASAP7_75t_R _31647_ (.A(_00101_),
    .Y(_11744_));
 AO22x1_ASAP7_75t_R _31648_ (.A1(net3026),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11744_),
    .Y(_11745_));
 AO21x1_ASAP7_75t_R _31649_ (.A1(net3736),
    .A2(_11734_),
    .B(_11745_),
    .Y(_04126_));
 AO22x1_ASAP7_75t_R _31650_ (.A1(net2922),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_06410_),
    .Y(_11746_));
 AO21x1_ASAP7_75t_R _31651_ (.A1(_09538_),
    .A2(_11734_),
    .B(_11746_),
    .Y(_04127_));
 INVx1_ASAP7_75t_R _31652_ (.A(_00656_),
    .Y(_11747_));
 AO22x1_ASAP7_75t_R _31653_ (.A1(net3460),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11747_),
    .Y(_11748_));
 AO21x1_ASAP7_75t_R _31654_ (.A1(net3673),
    .A2(_11734_),
    .B(_11748_),
    .Y(_04128_));
 INVx1_ASAP7_75t_R _31655_ (.A(_00108_),
    .Y(_11749_));
 AO22x1_ASAP7_75t_R _31656_ (.A1(net3253),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11749_),
    .Y(_11750_));
 AO21x1_ASAP7_75t_R _31657_ (.A1(net3707),
    .A2(_11734_),
    .B(_11750_),
    .Y(_04129_));
 INVx1_ASAP7_75t_R _31658_ (.A(_00111_),
    .Y(_11751_));
 AO22x1_ASAP7_75t_R _31659_ (.A1(net3475),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11751_),
    .Y(_11752_));
 AO21x1_ASAP7_75t_R _31660_ (.A1(net3541),
    .A2(_11734_),
    .B(_11752_),
    .Y(_04130_));
 AO22x1_ASAP7_75t_R _31661_ (.A1(net3452),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_08097_),
    .Y(_11753_));
 AO21x1_ASAP7_75t_R _31662_ (.A1(net3747),
    .A2(_11734_),
    .B(_11753_),
    .Y(_04131_));
 INVx1_ASAP7_75t_R _31663_ (.A(_00117_),
    .Y(_11754_));
 AO22x1_ASAP7_75t_R _31664_ (.A1(net3320),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11754_),
    .Y(_11755_));
 AO21x1_ASAP7_75t_R _31665_ (.A1(net3604),
    .A2(_11734_),
    .B(_11755_),
    .Y(_04132_));
 INVx1_ASAP7_75t_R _31666_ (.A(_00120_),
    .Y(_11756_));
 AO22x1_ASAP7_75t_R _31667_ (.A1(net3199),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11756_),
    .Y(_11757_));
 AO21x1_ASAP7_75t_R _31668_ (.A1(net3660),
    .A2(_11734_),
    .B(_11757_),
    .Y(_04133_));
 TAPCELL_ASAP7_75t_R PHY_189 ();
 TAPCELL_ASAP7_75t_R PHY_188 ();
 TAPCELL_ASAP7_75t_R PHY_187 ();
 INVx1_ASAP7_75t_R _31672_ (.A(_00123_),
    .Y(_11761_));
 AO22x1_ASAP7_75t_R _31673_ (.A1(net3336),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11761_),
    .Y(_11762_));
 AO21x1_ASAP7_75t_R _31674_ (.A1(net3573),
    .A2(_11734_),
    .B(_11762_),
    .Y(_04134_));
 INVx1_ASAP7_75t_R _31675_ (.A(_00126_),
    .Y(_11763_));
 AO22x1_ASAP7_75t_R _31676_ (.A1(net3430),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11763_),
    .Y(_11764_));
 AO21x1_ASAP7_75t_R _31677_ (.A1(net3721),
    .A2(_11734_),
    .B(_11764_),
    .Y(_04135_));
 INVx1_ASAP7_75t_R _31678_ (.A(_00129_),
    .Y(_11765_));
 AO22x1_ASAP7_75t_R _31679_ (.A1(net3276),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11765_),
    .Y(_11766_));
 AO21x1_ASAP7_75t_R _31680_ (.A1(net3683),
    .A2(_11734_),
    .B(_11766_),
    .Y(_04136_));
 INVx1_ASAP7_75t_R _31681_ (.A(_00132_),
    .Y(_11767_));
 AO22x1_ASAP7_75t_R _31682_ (.A1(net3344),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11767_),
    .Y(_11768_));
 AO21x1_ASAP7_75t_R _31683_ (.A1(net3678),
    .A2(_11734_),
    .B(_11768_),
    .Y(_04137_));
 INVx1_ASAP7_75t_R _31684_ (.A(_00135_),
    .Y(_11769_));
 AO22x1_ASAP7_75t_R _31685_ (.A1(net3220),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11769_),
    .Y(_11770_));
 AO21x1_ASAP7_75t_R _31686_ (.A1(net3691),
    .A2(_11734_),
    .B(_11770_),
    .Y(_04138_));
 INVx1_ASAP7_75t_R _31687_ (.A(_00138_),
    .Y(_11771_));
 AO22x1_ASAP7_75t_R _31688_ (.A1(net3215),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11771_),
    .Y(_11772_));
 AO21x1_ASAP7_75t_R _31689_ (.A1(_09638_),
    .A2(_11734_),
    .B(_11772_),
    .Y(_04139_));
 INVx1_ASAP7_75t_R _31690_ (.A(_00141_),
    .Y(_11773_));
 AO22x1_ASAP7_75t_R _31691_ (.A1(net3177),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11773_),
    .Y(_11774_));
 AO21x1_ASAP7_75t_R _31692_ (.A1(_09647_),
    .A2(_11734_),
    .B(_11774_),
    .Y(_04140_));
 AO22x1_ASAP7_75t_R _31693_ (.A1(net3366),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_08468_),
    .Y(_11775_));
 AO21x1_ASAP7_75t_R _31694_ (.A1(net3644),
    .A2(_11734_),
    .B(_11775_),
    .Y(_04141_));
 INVx1_ASAP7_75t_R _31695_ (.A(_00147_),
    .Y(_11776_));
 AO22x1_ASAP7_75t_R _31696_ (.A1(net3352),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11776_),
    .Y(_11777_));
 AO21x1_ASAP7_75t_R _31697_ (.A1(_09662_),
    .A2(_11734_),
    .B(_11777_),
    .Y(_04142_));
 INVx1_ASAP7_75t_R _31698_ (.A(_00150_),
    .Y(_11778_));
 AO22x1_ASAP7_75t_R _31699_ (.A1(net3328),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11778_),
    .Y(_11779_));
 AO21x1_ASAP7_75t_R _31700_ (.A1(net3594),
    .A2(_11734_),
    .B(_11779_),
    .Y(_04143_));
 INVx1_ASAP7_75t_R _31701_ (.A(_00153_),
    .Y(_11780_));
 AO22x1_ASAP7_75t_R _31702_ (.A1(net3245),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11780_),
    .Y(_11781_));
 AO21x1_ASAP7_75t_R _31703_ (.A1(_09676_),
    .A2(_11734_),
    .B(_11781_),
    .Y(_04144_));
 AO22x1_ASAP7_75t_R _31704_ (.A1(net3189),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_08584_),
    .Y(_11782_));
 AO21x1_ASAP7_75t_R _31705_ (.A1(net3611),
    .A2(_11734_),
    .B(_11782_),
    .Y(_04145_));
 INVx1_ASAP7_75t_R _31706_ (.A(_00159_),
    .Y(_11783_));
 AO22x1_ASAP7_75t_R _31707_ (.A1(net3229),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11783_),
    .Y(_11784_));
 AO21x1_ASAP7_75t_R _31708_ (.A1(net3698),
    .A2(_11734_),
    .B(_11784_),
    .Y(_04146_));
 INVx1_ASAP7_75t_R _31709_ (.A(_00161_),
    .Y(_11785_));
 AO22x1_ASAP7_75t_R _31710_ (.A1(net3268),
    .A2(_11736_),
    .B1(_11738_),
    .B2(_11785_),
    .Y(_11786_));
 AO21x1_ASAP7_75t_R _31711_ (.A1(_09698_),
    .A2(_11734_),
    .B(_11786_),
    .Y(_04147_));
 NAND3x1_ASAP7_75t_R _31712_ (.A(_06655_),
    .B(_07543_),
    .C(_11270_),
    .Y(_11787_));
 OA21x2_ASAP7_75t_R _31713_ (.A1(_11269_),
    .A2(_11787_),
    .B(_11268_),
    .Y(_11788_));
 CKINVDCx6p67_ASAP7_75t_R _31714_ (.A(_11788_),
    .Y(_11789_));
 TAPCELL_ASAP7_75t_R PHY_186 ();
 NOR2x1_ASAP7_75t_R _31716_ (.A(_02424_),
    .B(_11275_),
    .Y(_11791_));
 AO21x1_ASAP7_75t_R _31717_ (.A1(_11262_),
    .A2(_11275_),
    .B(_11791_),
    .Y(_11792_));
 OR2x2_ASAP7_75t_R _31718_ (.A(_11788_),
    .B(_11792_),
    .Y(_11793_));
 OA21x2_ASAP7_75t_R _31719_ (.A1(\cs_registers_i.mhpmcounter[2][32] ),
    .A2(_11789_),
    .B(_11793_),
    .Y(_04148_));
 NAND3x1_ASAP7_75t_R _31720_ (.A(_06655_),
    .B(_07543_),
    .C(_11270_),
    .Y(_11794_));
 OA21x2_ASAP7_75t_R _31721_ (.A1(_11794_),
    .A2(_11280_),
    .B(_11281_),
    .Y(_11795_));
 AO21x1_ASAP7_75t_R _31722_ (.A1(_02423_),
    .A2(_11286_),
    .B(_11795_),
    .Y(_11796_));
 OR3x1_ASAP7_75t_R _31723_ (.A(_02065_),
    .B(_02423_),
    .C(_11275_),
    .Y(_11797_));
 OAI21x1_ASAP7_75t_R _31724_ (.A1(net3647),
    .A2(_11284_),
    .B(_11797_),
    .Y(_11798_));
 AOI22x1_ASAP7_75t_R _31725_ (.A1(_02065_),
    .A2(_11796_),
    .B1(_11798_),
    .B2(_11789_),
    .Y(_04149_));
 TAPCELL_ASAP7_75t_R PHY_185 ();
 OAI21x1_ASAP7_75t_R _31727_ (.A1(_02426_),
    .A2(_11292_),
    .B(_11295_),
    .Y(_11800_));
 TAPCELL_ASAP7_75t_R PHY_184 ();
 NAND2x1_ASAP7_75t_R _31729_ (.A(_02064_),
    .B(_11788_),
    .Y(_11802_));
 OA21x2_ASAP7_75t_R _31730_ (.A1(_11788_),
    .A2(_11800_),
    .B(_11802_),
    .Y(_04150_));
 OR3x1_ASAP7_75t_R _31731_ (.A(_02063_),
    .B(_02425_),
    .C(_11275_),
    .Y(_11803_));
 OAI21x1_ASAP7_75t_R _31732_ (.A1(net3563),
    .A2(_11284_),
    .B(_11803_),
    .Y(_11804_));
 TAPCELL_ASAP7_75t_R PHY_183 ();
 AO21x1_ASAP7_75t_R _31734_ (.A1(_02425_),
    .A2(_11286_),
    .B(_11795_),
    .Y(_11806_));
 AOI22x1_ASAP7_75t_R _31735_ (.A1(_11789_),
    .A2(_11804_),
    .B1(_11806_),
    .B2(_02063_),
    .Y(_04151_));
 OAI21x1_ASAP7_75t_R _31736_ (.A1(_02428_),
    .A2(_11292_),
    .B(_11308_),
    .Y(_11807_));
 NAND2x1_ASAP7_75t_R _31737_ (.A(_02062_),
    .B(_11788_),
    .Y(_11808_));
 OA21x2_ASAP7_75t_R _31738_ (.A1(_11788_),
    .A2(_11807_),
    .B(_11808_),
    .Y(_04152_));
 OR3x1_ASAP7_75t_R _31739_ (.A(_02061_),
    .B(_02427_),
    .C(_11275_),
    .Y(_11809_));
 OAI21x1_ASAP7_75t_R _31740_ (.A1(net3632),
    .A2(_11284_),
    .B(_11809_),
    .Y(_11810_));
 AO21x1_ASAP7_75t_R _31741_ (.A1(_02427_),
    .A2(_11286_),
    .B(_11795_),
    .Y(_11811_));
 AOI22x1_ASAP7_75t_R _31742_ (.A1(_11789_),
    .A2(_11810_),
    .B1(_11811_),
    .B2(_02061_),
    .Y(_04153_));
 OAI21x1_ASAP7_75t_R _31743_ (.A1(_02430_),
    .A2(_11275_),
    .B(_11315_),
    .Y(_11812_));
 NAND2x1_ASAP7_75t_R _31744_ (.A(_02060_),
    .B(_11788_),
    .Y(_11813_));
 OA21x2_ASAP7_75t_R _31745_ (.A1(_11788_),
    .A2(_11812_),
    .B(_11813_),
    .Y(_04154_));
 INVx5_ASAP7_75t_R _31746_ (.A(_11795_),
    .Y(_11814_));
 OR3x4_ASAP7_75t_R _31747_ (.A(_07929_),
    .B(_11111_),
    .C(_11119_),
    .Y(_11815_));
 TAPCELL_ASAP7_75t_R PHY_182 ();
 TAPCELL_ASAP7_75t_R PHY_181 ();
 OR3x1_ASAP7_75t_R _31750_ (.A(_02059_),
    .B(_02429_),
    .C(_11299_),
    .Y(_11818_));
 OAI21x1_ASAP7_75t_R _31751_ (.A1(net3615),
    .A2(_11815_),
    .B(_11818_),
    .Y(_11819_));
 AO21x1_ASAP7_75t_R _31752_ (.A1(_02429_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11820_));
 AOI22x1_ASAP7_75t_R _31753_ (.A1(_11814_),
    .A2(_11819_),
    .B1(_11820_),
    .B2(_02059_),
    .Y(_04155_));
 OAI21x1_ASAP7_75t_R _31754_ (.A1(_02432_),
    .A2(_11275_),
    .B(_11321_),
    .Y(_11821_));
 NAND2x1_ASAP7_75t_R _31755_ (.A(_02058_),
    .B(_11788_),
    .Y(_11822_));
 OA21x2_ASAP7_75t_R _31756_ (.A1(_11788_),
    .A2(_11821_),
    .B(_11822_),
    .Y(_04156_));
 OR3x1_ASAP7_75t_R _31757_ (.A(_02057_),
    .B(_02431_),
    .C(_11299_),
    .Y(_11823_));
 OAI21x1_ASAP7_75t_R _31758_ (.A1(net3716),
    .A2(_11815_),
    .B(_11823_),
    .Y(_11824_));
 AO21x1_ASAP7_75t_R _31759_ (.A1(_02431_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11825_));
 AOI22x1_ASAP7_75t_R _31760_ (.A1(_11814_),
    .A2(_11824_),
    .B1(_11825_),
    .B2(_02057_),
    .Y(_04157_));
 OAI21x1_ASAP7_75t_R _31761_ (.A1(_02434_),
    .A2(_11299_),
    .B(_11329_),
    .Y(_11826_));
 NAND2x1_ASAP7_75t_R _31762_ (.A(_02056_),
    .B(_11788_),
    .Y(_11827_));
 OA21x2_ASAP7_75t_R _31763_ (.A1(_11788_),
    .A2(_11826_),
    .B(_11827_),
    .Y(_04158_));
 OR3x1_ASAP7_75t_R _31764_ (.A(_02055_),
    .B(_02433_),
    .C(_11299_),
    .Y(_11828_));
 OAI21x1_ASAP7_75t_R _31765_ (.A1(_09538_),
    .A2(_11815_),
    .B(_11828_),
    .Y(_11829_));
 AO21x1_ASAP7_75t_R _31766_ (.A1(_02433_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11830_));
 AOI22x1_ASAP7_75t_R _31767_ (.A1(_11814_),
    .A2(_11829_),
    .B1(_11830_),
    .B2(_02055_),
    .Y(_04159_));
 OAI21x1_ASAP7_75t_R _31768_ (.A1(_02436_),
    .A2(_11275_),
    .B(_11336_),
    .Y(_11831_));
 TAPCELL_ASAP7_75t_R PHY_180 ();
 NAND2x1_ASAP7_75t_R _31770_ (.A(_02054_),
    .B(_11788_),
    .Y(_11833_));
 OA21x2_ASAP7_75t_R _31771_ (.A1(_11788_),
    .A2(_11831_),
    .B(_11833_),
    .Y(_04160_));
 OR3x1_ASAP7_75t_R _31772_ (.A(_02053_),
    .B(_02435_),
    .C(_11299_),
    .Y(_11834_));
 OAI21x1_ASAP7_75t_R _31773_ (.A1(net3707),
    .A2(_11815_),
    .B(_11834_),
    .Y(_11835_));
 AO21x1_ASAP7_75t_R _31774_ (.A1(_02435_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11836_));
 AOI22x1_ASAP7_75t_R _31775_ (.A1(_11814_),
    .A2(net3708),
    .B1(_11836_),
    .B2(_02053_),
    .Y(_04161_));
 OAI21x1_ASAP7_75t_R _31776_ (.A1(_02438_),
    .A2(_11299_),
    .B(_11342_),
    .Y(_11837_));
 NAND2x1_ASAP7_75t_R _31777_ (.A(_02052_),
    .B(_11788_),
    .Y(_11838_));
 OA21x2_ASAP7_75t_R _31778_ (.A1(_11788_),
    .A2(_11837_),
    .B(_11838_),
    .Y(_04162_));
 INVx1_ASAP7_75t_R _31779_ (.A(_02437_),
    .Y(_11839_));
 AND3x1_ASAP7_75t_R _31780_ (.A(_02051_),
    .B(_11839_),
    .C(_11286_),
    .Y(_11840_));
 AO21x1_ASAP7_75t_R _31781_ (.A1(net3747),
    .A2(_11275_),
    .B(_11840_),
    .Y(_11841_));
 AO21x1_ASAP7_75t_R _31782_ (.A1(_02437_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11842_));
 INVx1_ASAP7_75t_R _31783_ (.A(_02051_),
    .Y(_11843_));
 AO22x1_ASAP7_75t_R _31784_ (.A1(_11789_),
    .A2(_11841_),
    .B1(_11842_),
    .B2(_11843_),
    .Y(_04163_));
 OAI21x1_ASAP7_75t_R _31785_ (.A1(_02440_),
    .A2(_11299_),
    .B(_11349_),
    .Y(_11844_));
 NAND2x1_ASAP7_75t_R _31786_ (.A(_02050_),
    .B(_11788_),
    .Y(_11845_));
 OA21x2_ASAP7_75t_R _31787_ (.A1(_11788_),
    .A2(_11844_),
    .B(_11845_),
    .Y(_04164_));
 INVx1_ASAP7_75t_R _31788_ (.A(_02049_),
    .Y(_11846_));
 AO21x1_ASAP7_75t_R _31789_ (.A1(_02439_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11847_));
 INVx1_ASAP7_75t_R _31790_ (.A(_02439_),
    .Y(_11848_));
 AND3x1_ASAP7_75t_R _31791_ (.A(_02049_),
    .B(_11848_),
    .C(_11286_),
    .Y(_11849_));
 AO21x1_ASAP7_75t_R _31792_ (.A1(net3660),
    .A2(_11299_),
    .B(_11849_),
    .Y(_11850_));
 AO22x1_ASAP7_75t_R _31793_ (.A1(_11846_),
    .A2(_11847_),
    .B1(_11850_),
    .B2(_11789_),
    .Y(_04165_));
 OAI21x1_ASAP7_75t_R _31794_ (.A1(_02442_),
    .A2(_11299_),
    .B(_11356_),
    .Y(_11851_));
 NAND2x1_ASAP7_75t_R _31795_ (.A(_02048_),
    .B(_11788_),
    .Y(_11852_));
 OA21x2_ASAP7_75t_R _31796_ (.A1(_11788_),
    .A2(_11851_),
    .B(_11852_),
    .Y(_04166_));
 INVx1_ASAP7_75t_R _31797_ (.A(_02441_),
    .Y(_11853_));
 AND3x1_ASAP7_75t_R _31798_ (.A(_02047_),
    .B(_11853_),
    .C(_11286_),
    .Y(_11854_));
 AO21x1_ASAP7_75t_R _31799_ (.A1(net3711),
    .A2(_11275_),
    .B(_11854_),
    .Y(_11855_));
 AO21x1_ASAP7_75t_R _31800_ (.A1(_02441_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11856_));
 INVx1_ASAP7_75t_R _31801_ (.A(_02047_),
    .Y(_11857_));
 AO22x1_ASAP7_75t_R _31802_ (.A1(_11789_),
    .A2(_11855_),
    .B1(_11856_),
    .B2(_11857_),
    .Y(_04167_));
 OAI21x1_ASAP7_75t_R _31803_ (.A1(_02444_),
    .A2(_11299_),
    .B(_11362_),
    .Y(_11858_));
 NAND2x1_ASAP7_75t_R _31804_ (.A(_02046_),
    .B(_11788_),
    .Y(_11859_));
 OA21x2_ASAP7_75t_R _31805_ (.A1(_11788_),
    .A2(_11858_),
    .B(_11859_),
    .Y(_04168_));
 INVx1_ASAP7_75t_R _31806_ (.A(_02045_),
    .Y(_11860_));
 AO21x1_ASAP7_75t_R _31807_ (.A1(_02443_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11861_));
 INVx1_ASAP7_75t_R _31808_ (.A(_02443_),
    .Y(_11862_));
 AND3x1_ASAP7_75t_R _31809_ (.A(_02045_),
    .B(_11862_),
    .C(_11286_),
    .Y(_11863_));
 AO21x1_ASAP7_75t_R _31810_ (.A1(_09623_),
    .A2(_11299_),
    .B(_11863_),
    .Y(_11864_));
 AO22x1_ASAP7_75t_R _31811_ (.A1(_11860_),
    .A2(_11861_),
    .B1(_11864_),
    .B2(_11789_),
    .Y(_04169_));
 OAI21x1_ASAP7_75t_R _31812_ (.A1(_02446_),
    .A2(_11299_),
    .B(_11368_),
    .Y(_11865_));
 NAND2x1_ASAP7_75t_R _31813_ (.A(_02044_),
    .B(_11788_),
    .Y(_11866_));
 OA21x2_ASAP7_75t_R _31814_ (.A1(_11788_),
    .A2(_11865_),
    .B(_11866_),
    .Y(_04170_));
 OR3x1_ASAP7_75t_R _31815_ (.A(_02043_),
    .B(_02445_),
    .C(_11299_),
    .Y(_11867_));
 OAI21x1_ASAP7_75t_R _31816_ (.A1(_09638_),
    .A2(_11815_),
    .B(_11867_),
    .Y(_11868_));
 AO21x1_ASAP7_75t_R _31817_ (.A1(_02445_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11869_));
 AOI22x1_ASAP7_75t_R _31818_ (.A1(_11814_),
    .A2(_11868_),
    .B1(_11869_),
    .B2(_02043_),
    .Y(_04171_));
 NOR2x1_ASAP7_75t_R _31819_ (.A(_02448_),
    .B(_11275_),
    .Y(_11870_));
 NAND2x1_ASAP7_75t_R _31820_ (.A(_02042_),
    .B(_11788_),
    .Y(_11871_));
 OA31x2_ASAP7_75t_R _31821_ (.A1(_11375_),
    .A2(_11788_),
    .A3(_11870_),
    .B1(_11871_),
    .Y(_04172_));
 INVx1_ASAP7_75t_R _31822_ (.A(_02041_),
    .Y(_11872_));
 AO21x1_ASAP7_75t_R _31823_ (.A1(_02447_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11873_));
 INVx1_ASAP7_75t_R _31824_ (.A(_02447_),
    .Y(_11874_));
 AND3x1_ASAP7_75t_R _31825_ (.A(_02041_),
    .B(_11874_),
    .C(_11286_),
    .Y(_11875_));
 AO21x1_ASAP7_75t_R _31826_ (.A1(net3639),
    .A2(_11275_),
    .B(_11875_),
    .Y(_11876_));
 AO22x1_ASAP7_75t_R _31827_ (.A1(_11872_),
    .A2(_11873_),
    .B1(_11876_),
    .B2(_11789_),
    .Y(_04173_));
 OAI21x1_ASAP7_75t_R _31828_ (.A1(_02450_),
    .A2(_11299_),
    .B(_11381_),
    .Y(_11877_));
 NAND2x1_ASAP7_75t_R _31829_ (.A(_02040_),
    .B(_11788_),
    .Y(_11878_));
 OA21x2_ASAP7_75t_R _31830_ (.A1(_11788_),
    .A2(_11877_),
    .B(_11878_),
    .Y(_04174_));
 INVx1_ASAP7_75t_R _31831_ (.A(_02039_),
    .Y(_11879_));
 AO21x1_ASAP7_75t_R _31832_ (.A1(_02449_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11880_));
 INVx1_ASAP7_75t_R _31833_ (.A(_02449_),
    .Y(_11881_));
 AND3x1_ASAP7_75t_R _31834_ (.A(_02039_),
    .B(_11881_),
    .C(_11286_),
    .Y(_11882_));
 AO21x1_ASAP7_75t_R _31835_ (.A1(net3594),
    .A2(_11275_),
    .B(_11882_),
    .Y(_11883_));
 AO22x1_ASAP7_75t_R _31836_ (.A1(_11879_),
    .A2(_11880_),
    .B1(_11883_),
    .B2(_11789_),
    .Y(_04175_));
 OAI21x1_ASAP7_75t_R _31837_ (.A1(_02452_),
    .A2(_11299_),
    .B(_11388_),
    .Y(_11884_));
 NAND2x1_ASAP7_75t_R _31838_ (.A(_02038_),
    .B(_11788_),
    .Y(_11885_));
 OA21x2_ASAP7_75t_R _31839_ (.A1(_11788_),
    .A2(_11884_),
    .B(_11885_),
    .Y(_04176_));
 OR3x1_ASAP7_75t_R _31840_ (.A(_02037_),
    .B(_02451_),
    .C(_11299_),
    .Y(_11886_));
 OAI21x1_ASAP7_75t_R _31841_ (.A1(net3611),
    .A2(_11815_),
    .B(_11886_),
    .Y(_11887_));
 AO21x1_ASAP7_75t_R _31842_ (.A1(_02451_),
    .A2(_11815_),
    .B(_11795_),
    .Y(_11888_));
 AOI22x1_ASAP7_75t_R _31843_ (.A1(_11814_),
    .A2(_11887_),
    .B1(_11888_),
    .B2(_02037_),
    .Y(_04177_));
 OAI21x1_ASAP7_75t_R _31844_ (.A1(_02454_),
    .A2(_11275_),
    .B(_11394_),
    .Y(_11889_));
 NAND2x1_ASAP7_75t_R _31845_ (.A(_02036_),
    .B(_11788_),
    .Y(_11890_));
 OA21x2_ASAP7_75t_R _31846_ (.A1(_11788_),
    .A2(_11889_),
    .B(_11890_),
    .Y(_04178_));
 OR3x1_ASAP7_75t_R _31847_ (.A(_02035_),
    .B(_02453_),
    .C(_11299_),
    .Y(_11891_));
 OAI21x1_ASAP7_75t_R _31848_ (.A1(_09698_),
    .A2(_11815_),
    .B(_11891_),
    .Y(_11892_));
 AO21x1_ASAP7_75t_R _31849_ (.A1(_02453_),
    .A2(_11286_),
    .B(_11795_),
    .Y(_11893_));
 AOI22x1_ASAP7_75t_R _31850_ (.A1(_11789_),
    .A2(_11892_),
    .B1(_11893_),
    .B2(_02035_),
    .Y(_04179_));
 NAND3x2_ASAP7_75t_R _31851_ (.B(_11087_),
    .C(_11096_),
    .Y(_11894_),
    .A(_05693_));
 TAPCELL_ASAP7_75t_R PHY_179 ();
 NAND2x1_ASAP7_75t_R _31853_ (.A(_02034_),
    .B(_11894_),
    .Y(_11896_));
 OA21x2_ASAP7_75t_R _31854_ (.A1(_11159_),
    .A2(_11894_),
    .B(_11896_),
    .Y(_04180_));
 NAND2x1_ASAP7_75t_R _31855_ (.A(_02033_),
    .B(_11894_),
    .Y(_11897_));
 OA21x2_ASAP7_75t_R _31856_ (.A1(_09538_),
    .A2(_11894_),
    .B(_11897_),
    .Y(_04181_));
 NAND2x1_ASAP7_75t_R _31857_ (.A(_02032_),
    .B(_11894_),
    .Y(_11898_));
 OA21x2_ASAP7_75t_R _31858_ (.A1(net3673),
    .A2(_11894_),
    .B(_11898_),
    .Y(_04182_));
 NAND2x1_ASAP7_75t_R _31859_ (.A(_02031_),
    .B(_11894_),
    .Y(_11899_));
 OA21x2_ASAP7_75t_R _31860_ (.A1(net3707),
    .A2(_11894_),
    .B(_11899_),
    .Y(_04183_));
 NAND2x1_ASAP7_75t_R _31861_ (.A(_02030_),
    .B(_11894_),
    .Y(_11900_));
 OA21x2_ASAP7_75t_R _31862_ (.A1(net3747),
    .A2(_11894_),
    .B(_11900_),
    .Y(_04184_));
 INVx1_ASAP7_75t_R _31863_ (.A(_05746_),
    .Y(_11901_));
 AO221x2_ASAP7_75t_R _31864_ (.A1(_01719_),
    .A2(_01725_),
    .B1(_11901_),
    .B2(_13459_),
    .C(_06214_),
    .Y(_11902_));
 TAPCELL_ASAP7_75t_R PHY_178 ();
 TAPCELL_ASAP7_75t_R PHY_177 ();
 TAPCELL_ASAP7_75t_R PHY_176 ();
 TAPCELL_ASAP7_75t_R PHY_175 ();
 AND2x2_ASAP7_75t_R _31869_ (.A(_00385_),
    .B(_01746_),
    .Y(_11907_));
 AO21x1_ASAP7_75t_R _31870_ (.A1(_05659_),
    .A2(_01723_),
    .B(_11907_),
    .Y(_11908_));
 OR4x1_ASAP7_75t_R _31871_ (.A(_01312_),
    .B(_06207_),
    .C(_06211_),
    .D(_11908_),
    .Y(_11909_));
 OAI21x1_ASAP7_75t_R _31872_ (.A1(_01641_),
    .A2(_11902_),
    .B(_11909_),
    .Y(_11910_));
 AND2x2_ASAP7_75t_R _31873_ (.A(_01311_),
    .B(_05557_),
    .Y(_11911_));
 AND4x2_ASAP7_75t_R _31874_ (.A(net310),
    .B(_05634_),
    .C(_05667_),
    .D(_11096_),
    .Y(_11912_));
 AND2x6_ASAP7_75t_R _31875_ (.A(_11086_),
    .B(_11912_),
    .Y(_11913_));
 TAPCELL_ASAP7_75t_R PHY_174 ();
 INVx1_ASAP7_75t_R _31877_ (.A(_02029_),
    .Y(_11915_));
 NAND2x2_ASAP7_75t_R _31878_ (.A(_11086_),
    .B(_11912_),
    .Y(_11916_));
 TAPCELL_ASAP7_75t_R PHY_173 ();
 AND3x1_ASAP7_75t_R _31880_ (.A(_11915_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11918_));
 AO221x1_ASAP7_75t_R _31881_ (.A1(_11910_),
    .A2(_11911_),
    .B1(_11913_),
    .B2(_11262_),
    .C(_11918_),
    .Y(_04185_));
 AND2x6_ASAP7_75t_R _31882_ (.A(_06385_),
    .B(_11675_),
    .Y(_11919_));
 TAPCELL_ASAP7_75t_R PHY_172 ();
 TAPCELL_ASAP7_75t_R PHY_171 ();
 TAPCELL_ASAP7_75t_R PHY_170 ();
 TAPCELL_ASAP7_75t_R PHY_169 ();
 TAPCELL_ASAP7_75t_R PHY_168 ();
 XNOR2x1_ASAP7_75t_R _31888_ (.B(_01720_),
    .Y(_11925_),
    .A(_01722_));
 TAPCELL_ASAP7_75t_R PHY_167 ();
 TAPCELL_ASAP7_75t_R PHY_166 ();
 TAPCELL_ASAP7_75t_R PHY_165 ();
 TAPCELL_ASAP7_75t_R PHY_164 ();
 AND2x2_ASAP7_75t_R _31893_ (.A(_00385_),
    .B(_00163_),
    .Y(_11930_));
 AO21x1_ASAP7_75t_R _31894_ (.A1(_05659_),
    .A2(_00164_),
    .B(_11930_),
    .Y(_11931_));
 TAPCELL_ASAP7_75t_R PHY_163 ();
 OA222x2_ASAP7_75t_R _31896_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01640_),
    .C1(_11931_),
    .C2(_01312_),
    .Y(_11933_));
 AOI21x1_ASAP7_75t_R _31897_ (.A1(_06211_),
    .A2(_11925_),
    .B(_11933_),
    .Y(_11934_));
 INVx1_ASAP7_75t_R _31898_ (.A(_02028_),
    .Y(_11935_));
 TAPCELL_ASAP7_75t_R PHY_162 ();
 AND3x1_ASAP7_75t_R _31900_ (.A(_11935_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11937_));
 AO221x1_ASAP7_75t_R _31901_ (.A1(net3647),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11934_),
    .C(_11937_),
    .Y(_04186_));
 TAPCELL_ASAP7_75t_R PHY_161 ();
 AND2x2_ASAP7_75t_R _31903_ (.A(_00385_),
    .B(_00165_),
    .Y(_11939_));
 AO21x1_ASAP7_75t_R _31904_ (.A1(_05659_),
    .A2(_00166_),
    .B(_11939_),
    .Y(_11940_));
 OAI22x1_ASAP7_75t_R _31905_ (.A1(_01639_),
    .A2(_11902_),
    .B1(_11940_),
    .B2(_01312_),
    .Y(_11941_));
 CKINVDCx16_ASAP7_75t_R _31906_ (.A(_01722_),
    .Y(_11942_));
 TAPCELL_ASAP7_75t_R PHY_160 ();
 NAND2x1_ASAP7_75t_R _31908_ (.A(_00167_),
    .B(_11942_),
    .Y(_11944_));
 OA211x2_ASAP7_75t_R _31909_ (.A1(\cs_registers_i.pc_id_i[2] ),
    .A2(_11942_),
    .B(_06211_),
    .C(_11944_),
    .Y(_11945_));
 AO21x2_ASAP7_75t_R _31910_ (.A1(_06205_),
    .A2(_11941_),
    .B(_11945_),
    .Y(_11946_));
 INVx1_ASAP7_75t_R _31911_ (.A(_02027_),
    .Y(_11947_));
 AND3x1_ASAP7_75t_R _31912_ (.A(_11947_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11948_));
 AO221x1_ASAP7_75t_R _31913_ (.A1(_11159_),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11946_),
    .C(_11948_),
    .Y(_04187_));
 TAPCELL_ASAP7_75t_R PHY_159 ();
 AND2x2_ASAP7_75t_R _31915_ (.A(_00385_),
    .B(_00168_),
    .Y(_11950_));
 AO21x1_ASAP7_75t_R _31916_ (.A1(_05659_),
    .A2(_00169_),
    .B(_11950_),
    .Y(_11951_));
 OAI22x1_ASAP7_75t_R _31917_ (.A1(_01638_),
    .A2(_11902_),
    .B1(_11951_),
    .B2(_01312_),
    .Y(_11952_));
 TAPCELL_ASAP7_75t_R PHY_158 ();
 TAPCELL_ASAP7_75t_R PHY_157 ();
 NAND2x1_ASAP7_75t_R _31920_ (.A(_11942_),
    .B(_00171_),
    .Y(_11955_));
 OA211x2_ASAP7_75t_R _31921_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[3] ),
    .B(_06211_),
    .C(_11955_),
    .Y(_11956_));
 AO21x1_ASAP7_75t_R _31922_ (.A1(_06205_),
    .A2(_11952_),
    .B(_11956_),
    .Y(_11957_));
 INVx1_ASAP7_75t_R _31923_ (.A(_02026_),
    .Y(_11958_));
 AND3x1_ASAP7_75t_R _31924_ (.A(_11958_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11959_));
 AO221x1_ASAP7_75t_R _31925_ (.A1(net3544),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11957_),
    .C(_11959_),
    .Y(_04188_));
 NOR2x1_ASAP7_75t_R _31926_ (.A(_01722_),
    .B(_02520_),
    .Y(_11960_));
 XNOR2x2_ASAP7_75t_R _31927_ (.A(_15051_),
    .B(_11960_),
    .Y(_11961_));
 AND2x2_ASAP7_75t_R _31928_ (.A(_00385_),
    .B(_00172_),
    .Y(_11962_));
 AO21x1_ASAP7_75t_R _31929_ (.A1(_05659_),
    .A2(_00173_),
    .B(_11962_),
    .Y(_11963_));
 OA222x2_ASAP7_75t_R _31930_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01637_),
    .C1(_11963_),
    .C2(_01312_),
    .Y(_11964_));
 AOI21x1_ASAP7_75t_R _31931_ (.A1(_06211_),
    .A2(_11961_),
    .B(_11964_),
    .Y(_11965_));
 INVx1_ASAP7_75t_R _31932_ (.A(_02025_),
    .Y(_11966_));
 AND3x1_ASAP7_75t_R _31933_ (.A(_11966_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11967_));
 AO221x1_ASAP7_75t_R _31934_ (.A1(net3379),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11965_),
    .C(_11967_),
    .Y(_04189_));
 AND2x2_ASAP7_75t_R _31935_ (.A(_00385_),
    .B(_00175_),
    .Y(_11968_));
 AO21x1_ASAP7_75t_R _31936_ (.A1(_05659_),
    .A2(_00176_),
    .B(_11968_),
    .Y(_11969_));
 OAI22x1_ASAP7_75t_R _31937_ (.A1(_01636_),
    .A2(_11902_),
    .B1(_11969_),
    .B2(_01312_),
    .Y(_11970_));
 TAPCELL_ASAP7_75t_R PHY_156 ();
 NAND2x1_ASAP7_75t_R _31939_ (.A(_11942_),
    .B(_00178_),
    .Y(_11972_));
 OA211x2_ASAP7_75t_R _31940_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[5] ),
    .B(_06211_),
    .C(_11972_),
    .Y(_11973_));
 AO21x2_ASAP7_75t_R _31941_ (.A1(_06205_),
    .A2(_11970_),
    .B(_11973_),
    .Y(_11974_));
 INVx1_ASAP7_75t_R _31942_ (.A(_02024_),
    .Y(_11975_));
 AND3x1_ASAP7_75t_R _31943_ (.A(_11975_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11976_));
 AO221x1_ASAP7_75t_R _31944_ (.A1(net3632),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11974_),
    .C(_11976_),
    .Y(_04190_));
 INVx1_ASAP7_75t_R _31945_ (.A(_02023_),
    .Y(_11977_));
 NOR2x1_ASAP7_75t_R _31946_ (.A(_01722_),
    .B(_02521_),
    .Y(_11978_));
 XNOR2x1_ASAP7_75t_R _31947_ (.B(_11978_),
    .Y(_11979_),
    .A(_15169_));
 AND2x2_ASAP7_75t_R _31948_ (.A(_00278_),
    .B(_00385_),
    .Y(_11980_));
 AO21x1_ASAP7_75t_R _31949_ (.A1(_05659_),
    .A2(_00179_),
    .B(_11980_),
    .Y(_11981_));
 OA222x2_ASAP7_75t_R _31950_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01635_),
    .C1(_11981_),
    .C2(_01312_),
    .Y(_11982_));
 AOI21x1_ASAP7_75t_R _31951_ (.A1(_06211_),
    .A2(_11979_),
    .B(_11982_),
    .Y(_11983_));
 AO32x1_ASAP7_75t_R _31952_ (.A1(_11977_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_11983_),
    .Y(_11984_));
 AO21x1_ASAP7_75t_R _31953_ (.A1(_09504_),
    .A2(_11913_),
    .B(_11984_),
    .Y(_04191_));
 AND2x2_ASAP7_75t_R _31954_ (.A(_00323_),
    .B(_00385_),
    .Y(_11985_));
 AO21x1_ASAP7_75t_R _31955_ (.A1(_05659_),
    .A2(_00181_),
    .B(_11985_),
    .Y(_11986_));
 OAI22x1_ASAP7_75t_R _31956_ (.A1(_01634_),
    .A2(_11902_),
    .B1(_11986_),
    .B2(_01312_),
    .Y(_11987_));
 NAND2x1_ASAP7_75t_R _31957_ (.A(_11942_),
    .B(_00183_),
    .Y(_11988_));
 OA211x2_ASAP7_75t_R _31958_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[7] ),
    .B(_06211_),
    .C(_11988_),
    .Y(_11989_));
 AO21x1_ASAP7_75t_R _31959_ (.A1(_06205_),
    .A2(_11987_),
    .B(_11989_),
    .Y(_11990_));
 INVx1_ASAP7_75t_R _31960_ (.A(_02022_),
    .Y(_11991_));
 AND3x1_ASAP7_75t_R _31961_ (.A(_11991_),
    .B(_11408_),
    .C(_11916_),
    .Y(_11992_));
 AO221x1_ASAP7_75t_R _31962_ (.A1(net3654),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_11990_),
    .C(_11992_),
    .Y(_04192_));
 INVx1_ASAP7_75t_R _31963_ (.A(_02021_),
    .Y(_11993_));
 OR2x2_ASAP7_75t_R _31964_ (.A(_01722_),
    .B(_02522_),
    .Y(_11994_));
 XNOR2x1_ASAP7_75t_R _31965_ (.B(_11994_),
    .Y(_11995_),
    .A(_00186_));
 AND2x2_ASAP7_75t_R _31966_ (.A(_00385_),
    .B(_00184_),
    .Y(_11996_));
 AO21x1_ASAP7_75t_R _31967_ (.A1(_05659_),
    .A2(_00185_),
    .B(_11996_),
    .Y(_11997_));
 OA222x2_ASAP7_75t_R _31968_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01633_),
    .C1(_11997_),
    .C2(_01312_),
    .Y(_11998_));
 AOI21x1_ASAP7_75t_R _31969_ (.A1(_06211_),
    .A2(_11995_),
    .B(_11998_),
    .Y(_11999_));
 AO32x1_ASAP7_75t_R _31970_ (.A1(_11993_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_11999_),
    .Y(_12000_));
 AO21x1_ASAP7_75t_R _31971_ (.A1(net3725),
    .A2(_11913_),
    .B(_12000_),
    .Y(_04193_));
 AND2x2_ASAP7_75t_R _31972_ (.A(_00385_),
    .B(_00187_),
    .Y(_12001_));
 AO21x1_ASAP7_75t_R _31973_ (.A1(_05659_),
    .A2(_00188_),
    .B(_12001_),
    .Y(_12002_));
 OAI22x1_ASAP7_75t_R _31974_ (.A1(_01632_),
    .A2(_11902_),
    .B1(_12002_),
    .B2(_01312_),
    .Y(_12003_));
 NAND2x1_ASAP7_75t_R _31975_ (.A(_11942_),
    .B(_00190_),
    .Y(_12004_));
 OA211x2_ASAP7_75t_R _31976_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[9] ),
    .B(_06211_),
    .C(_12004_),
    .Y(_12005_));
 AO21x1_ASAP7_75t_R _31977_ (.A1(_06205_),
    .A2(_12003_),
    .B(_12005_),
    .Y(_12006_));
 INVx1_ASAP7_75t_R _31978_ (.A(_02020_),
    .Y(_12007_));
 AND3x1_ASAP7_75t_R _31979_ (.A(_12007_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12008_));
 AO221x1_ASAP7_75t_R _31980_ (.A1(net3716),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12006_),
    .C(_12008_),
    .Y(_04194_));
 NOR2x1_ASAP7_75t_R _31981_ (.A(_01722_),
    .B(_02523_),
    .Y(_12009_));
 XNOR2x1_ASAP7_75t_R _31982_ (.B(_12009_),
    .Y(_12010_),
    .A(_15398_));
 AND2x2_ASAP7_75t_R _31983_ (.A(_00385_),
    .B(_00191_),
    .Y(_12011_));
 AO21x1_ASAP7_75t_R _31984_ (.A1(_05659_),
    .A2(_00192_),
    .B(_12011_),
    .Y(_12012_));
 OA222x2_ASAP7_75t_R _31985_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01631_),
    .C1(_12012_),
    .C2(_01312_),
    .Y(_12013_));
 AOI21x1_ASAP7_75t_R _31986_ (.A1(_06211_),
    .A2(_12010_),
    .B(_12013_),
    .Y(_12014_));
 INVx1_ASAP7_75t_R _31987_ (.A(_02019_),
    .Y(_12015_));
 TAPCELL_ASAP7_75t_R PHY_155 ();
 AND3x1_ASAP7_75t_R _31989_ (.A(_12015_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12017_));
 AO221x1_ASAP7_75t_R _31990_ (.A1(net3736),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12014_),
    .C(_12017_),
    .Y(_04195_));
 AND2x2_ASAP7_75t_R _31991_ (.A(_00385_),
    .B(_00194_),
    .Y(_12018_));
 AO21x1_ASAP7_75t_R _31992_ (.A1(_05659_),
    .A2(_00195_),
    .B(_12018_),
    .Y(_12019_));
 OAI22x1_ASAP7_75t_R _31993_ (.A1(_01630_),
    .A2(_11902_),
    .B1(_12019_),
    .B2(_01312_),
    .Y(_12020_));
 NAND2x1_ASAP7_75t_R _31994_ (.A(_11942_),
    .B(_00197_),
    .Y(_12021_));
 OA211x2_ASAP7_75t_R _31995_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[11] ),
    .B(_06211_),
    .C(_12021_),
    .Y(_12022_));
 AO21x1_ASAP7_75t_R _31996_ (.A1(_06205_),
    .A2(_12020_),
    .B(_12022_),
    .Y(_12023_));
 INVx1_ASAP7_75t_R _31997_ (.A(_02018_),
    .Y(_12024_));
 AND3x1_ASAP7_75t_R _31998_ (.A(_12024_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12025_));
 AO221x1_ASAP7_75t_R _31999_ (.A1(_09538_),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12023_),
    .C(_12025_),
    .Y(_04196_));
 INVx1_ASAP7_75t_R _32000_ (.A(_02017_),
    .Y(_12026_));
 OR2x2_ASAP7_75t_R _32001_ (.A(_01722_),
    .B(_02524_),
    .Y(_12027_));
 XNOR2x1_ASAP7_75t_R _32002_ (.B(_12027_),
    .Y(_12028_),
    .A(_00199_));
 AND2x2_ASAP7_75t_R _32003_ (.A(_00281_),
    .B(_00385_),
    .Y(_12029_));
 AO21x1_ASAP7_75t_R _32004_ (.A1(_05659_),
    .A2(_00198_),
    .B(_12029_),
    .Y(_12030_));
 OA222x2_ASAP7_75t_R _32005_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01629_),
    .C1(_12030_),
    .C2(_01312_),
    .Y(_12031_));
 AOI21x1_ASAP7_75t_R _32006_ (.A1(_06211_),
    .A2(_12028_),
    .B(_12031_),
    .Y(_12032_));
 AO32x1_ASAP7_75t_R _32007_ (.A1(_12026_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_12032_),
    .Y(_12033_));
 AO21x1_ASAP7_75t_R _32008_ (.A1(net3673),
    .A2(_11913_),
    .B(_12033_),
    .Y(_04197_));
 AND2x2_ASAP7_75t_R _32009_ (.A(_00282_),
    .B(_00385_),
    .Y(_12034_));
 AO21x1_ASAP7_75t_R _32010_ (.A1(_05659_),
    .A2(_00200_),
    .B(_12034_),
    .Y(_12035_));
 OAI22x1_ASAP7_75t_R _32011_ (.A1(_01628_),
    .A2(_11902_),
    .B1(_12035_),
    .B2(_01312_),
    .Y(_12036_));
 NAND2x1_ASAP7_75t_R _32012_ (.A(_11942_),
    .B(_00202_),
    .Y(_12037_));
 OA211x2_ASAP7_75t_R _32013_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[13] ),
    .B(_06211_),
    .C(_12037_),
    .Y(_12038_));
 AO21x1_ASAP7_75t_R _32014_ (.A1(_06205_),
    .A2(_12036_),
    .B(_12038_),
    .Y(_12039_));
 INVx1_ASAP7_75t_R _32015_ (.A(_02016_),
    .Y(_12040_));
 AND3x1_ASAP7_75t_R _32016_ (.A(_12040_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12041_));
 AO221x1_ASAP7_75t_R _32017_ (.A1(net3707),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12039_),
    .C(_12041_),
    .Y(_04198_));
 TAPCELL_ASAP7_75t_R PHY_154 ();
 NOR2x1_ASAP7_75t_R _32019_ (.A(_01722_),
    .B(_02525_),
    .Y(_12043_));
 XNOR2x1_ASAP7_75t_R _32020_ (.B(_12043_),
    .Y(_12044_),
    .A(_15775_));
 AND2x2_ASAP7_75t_R _32021_ (.A(_00279_),
    .B(_00385_),
    .Y(_12045_));
 AO21x1_ASAP7_75t_R _32022_ (.A1(_05659_),
    .A2(_00203_),
    .B(_12045_),
    .Y(_12046_));
 OA222x2_ASAP7_75t_R _32023_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01627_),
    .C1(_12046_),
    .C2(_01312_),
    .Y(_12047_));
 AOI21x1_ASAP7_75t_R _32024_ (.A1(_06211_),
    .A2(_12044_),
    .B(_12047_),
    .Y(_12048_));
 INVx1_ASAP7_75t_R _32025_ (.A(_02015_),
    .Y(_12049_));
 TAPCELL_ASAP7_75t_R PHY_153 ();
 AND3x1_ASAP7_75t_R _32027_ (.A(_12049_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12051_));
 AO221x1_ASAP7_75t_R _32028_ (.A1(net3541),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12048_),
    .C(_12051_),
    .Y(_04199_));
 AND2x2_ASAP7_75t_R _32029_ (.A(_00290_),
    .B(_00385_),
    .Y(_12052_));
 AO21x1_ASAP7_75t_R _32030_ (.A1(_05659_),
    .A2(_00205_),
    .B(_12052_),
    .Y(_12053_));
 OAI22x1_ASAP7_75t_R _32031_ (.A1(_01626_),
    .A2(_11902_),
    .B1(_12053_),
    .B2(_01312_),
    .Y(_12054_));
 NAND2x1_ASAP7_75t_R _32032_ (.A(_11942_),
    .B(_00207_),
    .Y(_12055_));
 OA211x2_ASAP7_75t_R _32033_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[15] ),
    .B(_06211_),
    .C(_12055_),
    .Y(_12056_));
 AO21x1_ASAP7_75t_R _32034_ (.A1(_06205_),
    .A2(_12054_),
    .B(_12056_),
    .Y(_12057_));
 INVx1_ASAP7_75t_R _32035_ (.A(_02014_),
    .Y(_12058_));
 AND3x1_ASAP7_75t_R _32036_ (.A(_12058_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12059_));
 AO221x1_ASAP7_75t_R _32037_ (.A1(net3747),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12057_),
    .C(_12059_),
    .Y(_04200_));
 TAPCELL_ASAP7_75t_R PHY_152 ();
 OR2x2_ASAP7_75t_R _32039_ (.A(_01722_),
    .B(_02526_),
    .Y(_12061_));
 XNOR2x1_ASAP7_75t_R _32040_ (.B(_12061_),
    .Y(_12062_),
    .A(_00208_));
 NAND2x2_ASAP7_75t_R _32041_ (.A(_00385_),
    .B(_06214_),
    .Y(_12063_));
 TAPCELL_ASAP7_75t_R PHY_151 ();
 OA222x2_ASAP7_75t_R _32043_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01625_),
    .C1(_12063_),
    .C2(net2214),
    .Y(_12065_));
 AOI21x1_ASAP7_75t_R _32044_ (.A1(_06211_),
    .A2(_12062_),
    .B(_12065_),
    .Y(_12066_));
 INVx1_ASAP7_75t_R _32045_ (.A(_02013_),
    .Y(_12067_));
 AND3x1_ASAP7_75t_R _32046_ (.A(_12067_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12068_));
 AO221x1_ASAP7_75t_R _32047_ (.A1(net3604),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12066_),
    .C(_12068_),
    .Y(_04201_));
 INVx1_ASAP7_75t_R _32048_ (.A(_02012_),
    .Y(_12069_));
 OAI22x1_ASAP7_75t_R _32049_ (.A1(_01624_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(net2303),
    .Y(_12070_));
 NAND2x1_ASAP7_75t_R _32050_ (.A(_11942_),
    .B(_00210_),
    .Y(_12071_));
 OA211x2_ASAP7_75t_R _32051_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[17] ),
    .B(_06211_),
    .C(_12071_),
    .Y(_12072_));
 AO21x1_ASAP7_75t_R _32052_ (.A1(_06205_),
    .A2(_12070_),
    .B(_12072_),
    .Y(_12073_));
 AO32x1_ASAP7_75t_R _32053_ (.A1(_12069_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_12073_),
    .Y(_12074_));
 AO21x1_ASAP7_75t_R _32054_ (.A1(net3660),
    .A2(_11913_),
    .B(_12074_),
    .Y(_04202_));
 OR2x2_ASAP7_75t_R _32055_ (.A(_01722_),
    .B(_02527_),
    .Y(_12075_));
 XNOR2x1_ASAP7_75t_R _32056_ (.B(_12075_),
    .Y(_12076_),
    .A(_00211_));
 OA222x2_ASAP7_75t_R _32057_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01623_),
    .C1(_12063_),
    .C2(_00287_),
    .Y(_12077_));
 AOI21x1_ASAP7_75t_R _32058_ (.A1(_06211_),
    .A2(_12076_),
    .B(_12077_),
    .Y(_12078_));
 INVx1_ASAP7_75t_R _32059_ (.A(_02011_),
    .Y(_12079_));
 AND3x1_ASAP7_75t_R _32060_ (.A(_12079_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12080_));
 AO221x1_ASAP7_75t_R _32061_ (.A1(net3557),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12078_),
    .C(_12080_),
    .Y(_04203_));
 OAI22x1_ASAP7_75t_R _32062_ (.A1(_01622_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(_00286_),
    .Y(_12081_));
 NAND2x1_ASAP7_75t_R _32063_ (.A(_11942_),
    .B(_00213_),
    .Y(_12082_));
 OA211x2_ASAP7_75t_R _32064_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[19] ),
    .B(_06211_),
    .C(_12082_),
    .Y(_12083_));
 AO21x1_ASAP7_75t_R _32065_ (.A1(_06205_),
    .A2(_12081_),
    .B(_12083_),
    .Y(_12084_));
 INVx1_ASAP7_75t_R _32066_ (.A(_02010_),
    .Y(_12085_));
 AND3x1_ASAP7_75t_R _32067_ (.A(_12085_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12086_));
 AO221x1_ASAP7_75t_R _32068_ (.A1(net3711),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12084_),
    .C(_12086_),
    .Y(_04204_));
 OR2x2_ASAP7_75t_R _32069_ (.A(_01722_),
    .B(_02528_),
    .Y(_12087_));
 XNOR2x1_ASAP7_75t_R _32070_ (.B(_12087_),
    .Y(_12088_),
    .A(_00214_));
 OA222x2_ASAP7_75t_R _32071_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01621_),
    .C1(_12063_),
    .C2(net375),
    .Y(_12089_));
 AOI21x1_ASAP7_75t_R _32072_ (.A1(_06211_),
    .A2(_12088_),
    .B(_12089_),
    .Y(_12090_));
 INVx1_ASAP7_75t_R _32073_ (.A(_02009_),
    .Y(_12091_));
 AND3x1_ASAP7_75t_R _32074_ (.A(_12091_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12092_));
 AO221x1_ASAP7_75t_R _32075_ (.A1(_09616_),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12090_),
    .C(_12092_),
    .Y(_04205_));
 INVx1_ASAP7_75t_R _32076_ (.A(_02008_),
    .Y(_12093_));
 OAI22x1_ASAP7_75t_R _32077_ (.A1(_01620_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(net2277),
    .Y(_12094_));
 NAND2x1_ASAP7_75t_R _32078_ (.A(_11942_),
    .B(_00216_),
    .Y(_12095_));
 OA211x2_ASAP7_75t_R _32079_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[21] ),
    .B(_06211_),
    .C(_12095_),
    .Y(_12096_));
 AO21x1_ASAP7_75t_R _32080_ (.A1(_06205_),
    .A2(_12094_),
    .B(_12096_),
    .Y(_12097_));
 AO32x1_ASAP7_75t_R _32081_ (.A1(_12093_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_12097_),
    .Y(_12098_));
 AO21x1_ASAP7_75t_R _32082_ (.A1(net3678),
    .A2(_11913_),
    .B(_12098_),
    .Y(_04206_));
 OR2x2_ASAP7_75t_R _32083_ (.A(_01722_),
    .B(_02529_),
    .Y(_12099_));
 XNOR2x1_ASAP7_75t_R _32084_ (.B(_12099_),
    .Y(_12100_),
    .A(_00217_));
 OA222x2_ASAP7_75t_R _32085_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01619_),
    .C1(_12063_),
    .C2(net2363),
    .Y(_12101_));
 AOI21x1_ASAP7_75t_R _32086_ (.A1(_06211_),
    .A2(_12100_),
    .B(_12101_),
    .Y(_12102_));
 INVx1_ASAP7_75t_R _32087_ (.A(_02007_),
    .Y(_12103_));
 AND3x1_ASAP7_75t_R _32088_ (.A(_12103_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12104_));
 AO221x1_ASAP7_75t_R _32089_ (.A1(net3691),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12102_),
    .C(_12104_),
    .Y(_04207_));
 OR3x1_ASAP7_75t_R _32090_ (.A(_06319_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12105_));
 OA222x2_ASAP7_75t_R _32091_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01618_),
    .C1(_12063_),
    .C2(net333),
    .Y(_12106_));
 OR2x2_ASAP7_75t_R _32092_ (.A(_01722_),
    .B(_00219_),
    .Y(_12107_));
 OA211x2_ASAP7_75t_R _32093_ (.A1(_11942_),
    .A2(_00218_),
    .B(_06211_),
    .C(_12107_),
    .Y(_12108_));
 OR3x2_ASAP7_75t_R _32094_ (.A(_12105_),
    .B(_12106_),
    .C(_12108_),
    .Y(_12109_));
 TAPCELL_ASAP7_75t_R PHY_150 ();
 OR3x1_ASAP7_75t_R _32096_ (.A(_02006_),
    .B(_11675_),
    .C(_11913_),
    .Y(_12111_));
 OA211x2_ASAP7_75t_R _32097_ (.A1(net3580),
    .A2(_11916_),
    .B(_12109_),
    .C(_12111_),
    .Y(_12112_));
 INVx1_ASAP7_75t_R _32098_ (.A(net3581),
    .Y(_04208_));
 OR2x2_ASAP7_75t_R _32099_ (.A(_01722_),
    .B(_02530_),
    .Y(_12113_));
 XNOR2x1_ASAP7_75t_R _32100_ (.B(_12113_),
    .Y(_12114_),
    .A(_00220_));
 OA222x2_ASAP7_75t_R _32101_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01617_),
    .C1(_12063_),
    .C2(_00244_),
    .Y(_12115_));
 AO21x1_ASAP7_75t_R _32102_ (.A1(_06211_),
    .A2(_12114_),
    .B(_12115_),
    .Y(_12116_));
 OR2x2_ASAP7_75t_R _32103_ (.A(_12105_),
    .B(_12116_),
    .Y(_12117_));
 OR3x1_ASAP7_75t_R _32104_ (.A(_02005_),
    .B(_11675_),
    .C(_11913_),
    .Y(_12118_));
 OR3x1_ASAP7_75t_R _32105_ (.A(net3531),
    .B(_09646_),
    .C(_11916_),
    .Y(_12119_));
 NAND3x1_ASAP7_75t_R _32106_ (.A(_12117_),
    .B(_12118_),
    .C(_12119_),
    .Y(_04209_));
 OAI22x1_ASAP7_75t_R _32107_ (.A1(_01616_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(_01743_),
    .Y(_12120_));
 NAND2x1_ASAP7_75t_R _32108_ (.A(_11942_),
    .B(_00222_),
    .Y(_12121_));
 OA211x2_ASAP7_75t_R _32109_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[25] ),
    .B(_06211_),
    .C(_12121_),
    .Y(_12122_));
 AO21x1_ASAP7_75t_R _32110_ (.A1(_06205_),
    .A2(_12120_),
    .B(_12122_),
    .Y(_12123_));
 INVx1_ASAP7_75t_R _32111_ (.A(_02004_),
    .Y(_12124_));
 AND3x1_ASAP7_75t_R _32112_ (.A(_12124_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12125_));
 AO221x1_ASAP7_75t_R _32113_ (.A1(net3639),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12123_),
    .C(_12125_),
    .Y(_04210_));
 OR2x2_ASAP7_75t_R _32114_ (.A(_01722_),
    .B(_02531_),
    .Y(_12126_));
 XNOR2x1_ASAP7_75t_R _32115_ (.B(_12126_),
    .Y(_12127_),
    .A(_00223_));
 OA222x2_ASAP7_75t_R _32116_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01615_),
    .C1(_12063_),
    .C2(_00283_),
    .Y(_12128_));
 AOI21x1_ASAP7_75t_R _32117_ (.A1(_06211_),
    .A2(_12127_),
    .B(_12128_),
    .Y(_12129_));
 INVx1_ASAP7_75t_R _32118_ (.A(_02003_),
    .Y(_12130_));
 AND3x1_ASAP7_75t_R _32119_ (.A(_12130_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12131_));
 AO221x1_ASAP7_75t_R _32120_ (.A1(_09662_),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12129_),
    .C(_12131_),
    .Y(_04211_));
 OAI22x1_ASAP7_75t_R _32121_ (.A1(_01614_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(_01742_),
    .Y(_12132_));
 NAND2x1_ASAP7_75t_R _32122_ (.A(_11942_),
    .B(_00225_),
    .Y(_12133_));
 OA211x2_ASAP7_75t_R _32123_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[27] ),
    .B(_06211_),
    .C(_12133_),
    .Y(_12134_));
 AO21x1_ASAP7_75t_R _32124_ (.A1(_06205_),
    .A2(_12132_),
    .B(_12134_),
    .Y(_12135_));
 INVx1_ASAP7_75t_R _32125_ (.A(_02002_),
    .Y(_12136_));
 AND3x1_ASAP7_75t_R _32126_ (.A(_12136_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12137_));
 AO221x1_ASAP7_75t_R _32127_ (.A1(net3594),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12135_),
    .C(_12137_),
    .Y(_04212_));
 OR2x2_ASAP7_75t_R _32128_ (.A(_01722_),
    .B(_02532_),
    .Y(_12138_));
 XNOR2x1_ASAP7_75t_R _32129_ (.B(_12138_),
    .Y(_12139_),
    .A(_00226_));
 OA222x2_ASAP7_75t_R _32130_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_01741_),
    .B2(_12063_),
    .C1(_11902_),
    .C2(_01613_),
    .Y(_12140_));
 AOI21x1_ASAP7_75t_R _32131_ (.A1(_06211_),
    .A2(_12139_),
    .B(_12140_),
    .Y(_12141_));
 INVx1_ASAP7_75t_R _32132_ (.A(_02001_),
    .Y(_12142_));
 AND3x1_ASAP7_75t_R _32133_ (.A(_12142_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12143_));
 AO221x1_ASAP7_75t_R _32134_ (.A1(_09676_),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12141_),
    .C(_12143_),
    .Y(_04213_));
 OAI22x1_ASAP7_75t_R _32135_ (.A1(_01612_),
    .A2(_11902_),
    .B1(_12063_),
    .B2(_01740_),
    .Y(_12144_));
 NAND2x1_ASAP7_75t_R _32136_ (.A(_11942_),
    .B(_00228_),
    .Y(_12145_));
 OA211x2_ASAP7_75t_R _32137_ (.A1(_11942_),
    .A2(\cs_registers_i.pc_id_i[29] ),
    .B(_06211_),
    .C(_12145_),
    .Y(_12146_));
 AO21x1_ASAP7_75t_R _32138_ (.A1(_06205_),
    .A2(_12144_),
    .B(_12146_),
    .Y(_12147_));
 INVx1_ASAP7_75t_R _32139_ (.A(_02000_),
    .Y(_12148_));
 AND3x1_ASAP7_75t_R _32140_ (.A(_12148_),
    .B(_11408_),
    .C(_11916_),
    .Y(_12149_));
 AO221x1_ASAP7_75t_R _32141_ (.A1(net3611),
    .A2(_11913_),
    .B1(_11919_),
    .B2(_12147_),
    .C(_12149_),
    .Y(_04214_));
 INVx1_ASAP7_75t_R _32142_ (.A(_01999_),
    .Y(_12150_));
 NOR2x1_ASAP7_75t_R _32143_ (.A(_01722_),
    .B(_02533_),
    .Y(_12151_));
 XNOR2x1_ASAP7_75t_R _32144_ (.B(_12151_),
    .Y(_12152_),
    .A(_05401_));
 OA222x2_ASAP7_75t_R _32145_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_01739_),
    .B2(_12063_),
    .C1(_11902_),
    .C2(_01611_),
    .Y(_12153_));
 AOI21x1_ASAP7_75t_R _32146_ (.A1(_06211_),
    .A2(_12152_),
    .B(_12153_),
    .Y(_12154_));
 AO32x1_ASAP7_75t_R _32147_ (.A1(_12150_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_12154_),
    .Y(_12155_));
 AO21x1_ASAP7_75t_R _32148_ (.A1(net3698),
    .A2(_11913_),
    .B(_12155_),
    .Y(_04215_));
 INVx1_ASAP7_75t_R _32149_ (.A(_01998_),
    .Y(_12156_));
 OR4x1_ASAP7_75t_R _32150_ (.A(_01722_),
    .B(_00227_),
    .C(_00229_),
    .D(_06094_),
    .Y(_12157_));
 XNOR2x1_ASAP7_75t_R _32151_ (.B(_12157_),
    .Y(_12158_),
    .A(_00230_));
 OA222x2_ASAP7_75t_R _32152_ (.A1(_01317_),
    .A2(_01721_),
    .B1(_11902_),
    .B2(_01610_),
    .C1(_12063_),
    .C2(_00280_),
    .Y(_12159_));
 AOI21x1_ASAP7_75t_R _32153_ (.A1(_06211_),
    .A2(_12158_),
    .B(_12159_),
    .Y(_12160_));
 AO32x1_ASAP7_75t_R _32154_ (.A1(_12156_),
    .A2(_11408_),
    .A3(_11916_),
    .B1(_11919_),
    .B2(_12160_),
    .Y(_12161_));
 AO21x1_ASAP7_75t_R _32155_ (.A1(_09698_),
    .A2(_11913_),
    .B(_12161_),
    .Y(_04216_));
 NAND2x1_ASAP7_75t_R _32156_ (.A(_01997_),
    .B(_11403_),
    .Y(_12162_));
 OA21x2_ASAP7_75t_R _32157_ (.A1(_09623_),
    .A2(_11403_),
    .B(_12162_),
    .Y(_04217_));
 NAND2x1_ASAP7_75t_R _32158_ (.A(_01996_),
    .B(_11403_),
    .Y(_12163_));
 OA21x2_ASAP7_75t_R _32159_ (.A1(net3660),
    .A2(_11403_),
    .B(_12163_),
    .Y(_04218_));
 NAND2x2_ASAP7_75t_R _32160_ (.A(_11087_),
    .B(_11912_),
    .Y(_12164_));
 TAPCELL_ASAP7_75t_R PHY_149 ();
 TAPCELL_ASAP7_75t_R PHY_148 ();
 NAND2x1_ASAP7_75t_R _32163_ (.A(_01995_),
    .B(_12164_),
    .Y(_12167_));
 OA21x2_ASAP7_75t_R _32164_ (.A1(_11262_),
    .A2(_12164_),
    .B(_12167_),
    .Y(_04219_));
 NAND2x1_ASAP7_75t_R _32165_ (.A(_01994_),
    .B(_12164_),
    .Y(_12168_));
 OA21x2_ASAP7_75t_R _32166_ (.A1(net3647),
    .A2(_12164_),
    .B(_12168_),
    .Y(_04220_));
 NAND2x1_ASAP7_75t_R _32167_ (.A(_01993_),
    .B(_12164_),
    .Y(_12169_));
 OA21x2_ASAP7_75t_R _32168_ (.A1(_11159_),
    .A2(_12164_),
    .B(_12169_),
    .Y(_04221_));
 NAND2x1_ASAP7_75t_R _32169_ (.A(_01992_),
    .B(_12164_),
    .Y(_12170_));
 OA21x2_ASAP7_75t_R _32170_ (.A1(net3544),
    .A2(_12164_),
    .B(_12170_),
    .Y(_04222_));
 NAND2x1_ASAP7_75t_R _32171_ (.A(_01991_),
    .B(_12164_),
    .Y(_12171_));
 OA21x2_ASAP7_75t_R _32172_ (.A1(net3379),
    .A2(_12164_),
    .B(_12171_),
    .Y(_04223_));
 NAND2x1_ASAP7_75t_R _32173_ (.A(_01990_),
    .B(_12164_),
    .Y(_12172_));
 OA21x2_ASAP7_75t_R _32174_ (.A1(net3632),
    .A2(_12164_),
    .B(_12172_),
    .Y(_04224_));
 NAND2x1_ASAP7_75t_R _32175_ (.A(_01989_),
    .B(_12164_),
    .Y(_12173_));
 OA21x2_ASAP7_75t_R _32176_ (.A1(_09504_),
    .A2(_12164_),
    .B(_12173_),
    .Y(_04225_));
 NAND2x1_ASAP7_75t_R _32177_ (.A(_01988_),
    .B(_12164_),
    .Y(_12174_));
 OA21x2_ASAP7_75t_R _32178_ (.A1(net3615),
    .A2(_12164_),
    .B(_12174_),
    .Y(_04226_));
 TAPCELL_ASAP7_75t_R PHY_147 ();
 NAND2x1_ASAP7_75t_R _32180_ (.A(_01987_),
    .B(_12164_),
    .Y(_12176_));
 OA21x2_ASAP7_75t_R _32181_ (.A1(net3725),
    .A2(_12164_),
    .B(_12176_),
    .Y(_04227_));
 NAND2x1_ASAP7_75t_R _32182_ (.A(_01986_),
    .B(_12164_),
    .Y(_12177_));
 OA21x2_ASAP7_75t_R _32183_ (.A1(net3716),
    .A2(_12164_),
    .B(_12177_),
    .Y(_04228_));
 TAPCELL_ASAP7_75t_R PHY_146 ();
 NAND2x1_ASAP7_75t_R _32185_ (.A(_01985_),
    .B(_12164_),
    .Y(_12179_));
 OA21x2_ASAP7_75t_R _32186_ (.A1(net3736),
    .A2(_12164_),
    .B(_12179_),
    .Y(_04229_));
 NAND2x1_ASAP7_75t_R _32187_ (.A(_01984_),
    .B(_12164_),
    .Y(_12180_));
 OA21x2_ASAP7_75t_R _32188_ (.A1(_09538_),
    .A2(_12164_),
    .B(_12180_),
    .Y(_04230_));
 NAND2x1_ASAP7_75t_R _32189_ (.A(_01983_),
    .B(_12164_),
    .Y(_12181_));
 OA21x2_ASAP7_75t_R _32190_ (.A1(net3673),
    .A2(_12164_),
    .B(_12181_),
    .Y(_04231_));
 NAND2x1_ASAP7_75t_R _32191_ (.A(_01982_),
    .B(_12164_),
    .Y(_12182_));
 OA21x2_ASAP7_75t_R _32192_ (.A1(net3707),
    .A2(_12164_),
    .B(_12182_),
    .Y(_04232_));
 NAND2x1_ASAP7_75t_R _32193_ (.A(_01981_),
    .B(_12164_),
    .Y(_12183_));
 OA21x2_ASAP7_75t_R _32194_ (.A1(net3541),
    .A2(_12164_),
    .B(_12183_),
    .Y(_04233_));
 NAND2x1_ASAP7_75t_R _32195_ (.A(_01980_),
    .B(_12164_),
    .Y(_12184_));
 OA21x2_ASAP7_75t_R _32196_ (.A1(net3747),
    .A2(_12164_),
    .B(_12184_),
    .Y(_04234_));
 NAND2x1_ASAP7_75t_R _32197_ (.A(_01979_),
    .B(_12164_),
    .Y(_12185_));
 OA21x2_ASAP7_75t_R _32198_ (.A1(net3604),
    .A2(_12164_),
    .B(_12185_),
    .Y(_04235_));
 NAND2x1_ASAP7_75t_R _32199_ (.A(_01978_),
    .B(_12164_),
    .Y(_12186_));
 OA21x2_ASAP7_75t_R _32200_ (.A1(net3660),
    .A2(_12164_),
    .B(_12186_),
    .Y(_04236_));
 TAPCELL_ASAP7_75t_R PHY_145 ();
 NAND2x1_ASAP7_75t_R _32202_ (.A(_01977_),
    .B(_12164_),
    .Y(_12188_));
 OA21x2_ASAP7_75t_R _32203_ (.A1(net3557),
    .A2(_12164_),
    .B(_12188_),
    .Y(_04237_));
 NAND2x1_ASAP7_75t_R _32204_ (.A(_01976_),
    .B(_12164_),
    .Y(_12189_));
 OA21x2_ASAP7_75t_R _32205_ (.A1(net3721),
    .A2(_12164_),
    .B(_12189_),
    .Y(_04238_));
 TAPCELL_ASAP7_75t_R PHY_144 ();
 NAND2x1_ASAP7_75t_R _32207_ (.A(_01975_),
    .B(_12164_),
    .Y(_12191_));
 OA21x2_ASAP7_75t_R _32208_ (.A1(net3683),
    .A2(_12164_),
    .B(_12191_),
    .Y(_04239_));
 NAND2x1_ASAP7_75t_R _32209_ (.A(_01974_),
    .B(_12164_),
    .Y(_12192_));
 OA21x2_ASAP7_75t_R _32210_ (.A1(_09623_),
    .A2(_12164_),
    .B(_12192_),
    .Y(_04240_));
 NAND2x1_ASAP7_75t_R _32211_ (.A(_01973_),
    .B(_12164_),
    .Y(_12193_));
 OA21x2_ASAP7_75t_R _32212_ (.A1(net3691),
    .A2(_12164_),
    .B(_12193_),
    .Y(_04241_));
 NAND2x1_ASAP7_75t_R _32213_ (.A(_01972_),
    .B(_12164_),
    .Y(_12194_));
 OA21x2_ASAP7_75t_R _32214_ (.A1(_09638_),
    .A2(_12164_),
    .B(_12194_),
    .Y(_04242_));
 INVx1_ASAP7_75t_R _32215_ (.A(_01971_),
    .Y(_12195_));
 NOR3x1_ASAP7_75t_R _32216_ (.A(net3531),
    .B(_09646_),
    .C(_12164_),
    .Y(_12196_));
 AO21x1_ASAP7_75t_R _32217_ (.A1(_12195_),
    .A2(_12164_),
    .B(_12196_),
    .Y(_04243_));
 NAND2x1_ASAP7_75t_R _32218_ (.A(_01970_),
    .B(_12164_),
    .Y(_12197_));
 OA21x2_ASAP7_75t_R _32219_ (.A1(net3639),
    .A2(_12164_),
    .B(_12197_),
    .Y(_04244_));
 NAND2x1_ASAP7_75t_R _32220_ (.A(_01969_),
    .B(_12164_),
    .Y(_12198_));
 OA21x2_ASAP7_75t_R _32221_ (.A1(_09662_),
    .A2(_12164_),
    .B(_12198_),
    .Y(_04245_));
 NAND2x1_ASAP7_75t_R _32222_ (.A(_01968_),
    .B(_12164_),
    .Y(_12199_));
 OA21x2_ASAP7_75t_R _32223_ (.A1(net3594),
    .A2(_12164_),
    .B(_12199_),
    .Y(_04246_));
 NAND2x1_ASAP7_75t_R _32224_ (.A(_01967_),
    .B(_12164_),
    .Y(_12200_));
 OA21x2_ASAP7_75t_R _32225_ (.A1(_09676_),
    .A2(_12164_),
    .B(_12200_),
    .Y(_04247_));
 NAND2x1_ASAP7_75t_R _32226_ (.A(_01966_),
    .B(_12164_),
    .Y(_12201_));
 OA21x2_ASAP7_75t_R _32227_ (.A1(net3611),
    .A2(_12164_),
    .B(_12201_),
    .Y(_04248_));
 NAND2x1_ASAP7_75t_R _32228_ (.A(_01965_),
    .B(_12164_),
    .Y(_12202_));
 OA21x2_ASAP7_75t_R _32229_ (.A1(_09691_),
    .A2(_12164_),
    .B(_12202_),
    .Y(_04249_));
 NAND2x1_ASAP7_75t_R _32230_ (.A(_01964_),
    .B(_12164_),
    .Y(_12203_));
 OA21x2_ASAP7_75t_R _32231_ (.A1(_09698_),
    .A2(_12164_),
    .B(_12203_),
    .Y(_04250_));
 AND3x1_ASAP7_75t_R _32232_ (.A(_05647_),
    .B(_05707_),
    .C(_07450_),
    .Y(_12204_));
 INVx1_ASAP7_75t_R _32233_ (.A(_12204_),
    .Y(_12205_));
 NOR2x2_ASAP7_75t_R _32234_ (.A(_11119_),
    .B(_12205_),
    .Y(_12206_));
 TAPCELL_ASAP7_75t_R PHY_143 ();
 TAPCELL_ASAP7_75t_R PHY_142 ();
 NOR2x1_ASAP7_75t_R _32237_ (.A(_01963_),
    .B(_12206_),
    .Y(_12209_));
 AO21x1_ASAP7_75t_R _32238_ (.A1(net3604),
    .A2(_12206_),
    .B(_12209_),
    .Y(_04251_));
 NOR2x1_ASAP7_75t_R _32239_ (.A(_01962_),
    .B(_12206_),
    .Y(_12210_));
 AO21x1_ASAP7_75t_R _32240_ (.A1(net3660),
    .A2(_12206_),
    .B(_12210_),
    .Y(_04252_));
 TAPCELL_ASAP7_75t_R PHY_141 ();
 NOR2x1_ASAP7_75t_R _32242_ (.A(_01961_),
    .B(_12206_),
    .Y(_12212_));
 AO21x1_ASAP7_75t_R _32243_ (.A1(net3557),
    .A2(_12206_),
    .B(_12212_),
    .Y(_04253_));
 NOR2x1_ASAP7_75t_R _32244_ (.A(_01960_),
    .B(_12206_),
    .Y(_12213_));
 AO21x1_ASAP7_75t_R _32245_ (.A1(net3711),
    .A2(_12206_),
    .B(_12213_),
    .Y(_04254_));
 NOR2x1_ASAP7_75t_R _32246_ (.A(_01959_),
    .B(_12206_),
    .Y(_12214_));
 AO21x1_ASAP7_75t_R _32247_ (.A1(net3683),
    .A2(_12206_),
    .B(_12214_),
    .Y(_04255_));
 NOR2x1_ASAP7_75t_R _32248_ (.A(_01958_),
    .B(_12206_),
    .Y(_12215_));
 AO21x1_ASAP7_75t_R _32249_ (.A1(net3678),
    .A2(_12206_),
    .B(_12215_),
    .Y(_04256_));
 NOR2x1_ASAP7_75t_R _32250_ (.A(_01957_),
    .B(_12206_),
    .Y(_12216_));
 AO21x1_ASAP7_75t_R _32251_ (.A1(net3691),
    .A2(_12206_),
    .B(_12216_),
    .Y(_04257_));
 NOR2x1_ASAP7_75t_R _32252_ (.A(_01956_),
    .B(_12206_),
    .Y(_12217_));
 AO21x1_ASAP7_75t_R _32253_ (.A1(_09638_),
    .A2(_12206_),
    .B(_12217_),
    .Y(_04258_));
 NAND2x1_ASAP7_75t_R _32254_ (.A(_11096_),
    .B(_12204_),
    .Y(_12218_));
 AND2x2_ASAP7_75t_R _32255_ (.A(_06256_),
    .B(_12218_),
    .Y(_12219_));
 AO21x1_ASAP7_75t_R _32256_ (.A1(_09647_),
    .A2(_12206_),
    .B(_12219_),
    .Y(_04259_));
 NOR2x1_ASAP7_75t_R _32257_ (.A(_01954_),
    .B(_12206_),
    .Y(_12220_));
 AO21x1_ASAP7_75t_R _32258_ (.A1(net3639),
    .A2(_12206_),
    .B(_12220_),
    .Y(_04260_));
 NOR2x1_ASAP7_75t_R _32259_ (.A(_01953_),
    .B(_12206_),
    .Y(_12221_));
 AO21x1_ASAP7_75t_R _32260_ (.A1(_09662_),
    .A2(_12206_),
    .B(_12221_),
    .Y(_04261_));
 NOR2x1_ASAP7_75t_R _32261_ (.A(_01952_),
    .B(_12206_),
    .Y(_12222_));
 AO21x1_ASAP7_75t_R _32262_ (.A1(net3594),
    .A2(_12206_),
    .B(_12222_),
    .Y(_04262_));
 NOR2x1_ASAP7_75t_R _32263_ (.A(_01951_),
    .B(_12206_),
    .Y(_12223_));
 AO21x1_ASAP7_75t_R _32264_ (.A1(_09676_),
    .A2(_12206_),
    .B(_12223_),
    .Y(_04263_));
 NOR2x1_ASAP7_75t_R _32265_ (.A(_01950_),
    .B(_12206_),
    .Y(_12224_));
 AO21x1_ASAP7_75t_R _32266_ (.A1(net3611),
    .A2(_12206_),
    .B(_12224_),
    .Y(_04264_));
 NOR2x1_ASAP7_75t_R _32267_ (.A(_01949_),
    .B(_12206_),
    .Y(_12225_));
 AO21x1_ASAP7_75t_R _32268_ (.A1(net3698),
    .A2(_12206_),
    .B(_12225_),
    .Y(_04265_));
 NOR2x1_ASAP7_75t_R _32269_ (.A(_01948_),
    .B(_12206_),
    .Y(_12226_));
 AO21x1_ASAP7_75t_R _32270_ (.A1(_09538_),
    .A2(_12206_),
    .B(_12226_),
    .Y(_04266_));
 NOR2x1_ASAP7_75t_R _32271_ (.A(_01947_),
    .B(_12206_),
    .Y(_12227_));
 AO21x1_ASAP7_75t_R _32272_ (.A1(net3615),
    .A2(_12206_),
    .B(_12227_),
    .Y(_04267_));
 NOR2x1_ASAP7_75t_R _32273_ (.A(_01946_),
    .B(_12206_),
    .Y(_12228_));
 AO21x1_ASAP7_75t_R _32274_ (.A1(net3544),
    .A2(_12206_),
    .B(_12228_),
    .Y(_04268_));
 AND3x1_ASAP7_75t_R _32275_ (.A(_05601_),
    .B(_05630_),
    .C(_11078_),
    .Y(_12229_));
 NAND2x1_ASAP7_75t_R _32276_ (.A(_07440_),
    .B(_12229_),
    .Y(_12230_));
 AND2x6_ASAP7_75t_R _32277_ (.A(_11408_),
    .B(_11414_),
    .Y(_12231_));
 OAI21x1_ASAP7_75t_R _32278_ (.A1(_11285_),
    .A2(_12230_),
    .B(_12231_),
    .Y(_12232_));
 TAPCELL_ASAP7_75t_R PHY_140 ();
 OAI22x1_ASAP7_75t_R _32280_ (.A1(_01907_),
    .A2(_11414_),
    .B1(_12232_),
    .B2(_01945_),
    .Y(_04269_));
 OA21x2_ASAP7_75t_R _32281_ (.A1(_11285_),
    .A2(_12230_),
    .B(_12231_),
    .Y(_12234_));
 TAPCELL_ASAP7_75t_R PHY_139 ();
 NAND2x1_ASAP7_75t_R _32283_ (.A(_09452_),
    .B(_11414_),
    .Y(_12236_));
 OR2x2_ASAP7_75t_R _32284_ (.A(_01906_),
    .B(_11414_),
    .Y(_12237_));
 AND4x1_ASAP7_75t_R _32285_ (.A(_11406_),
    .B(_12232_),
    .C(_12236_),
    .D(_12237_),
    .Y(_12238_));
 AO221x1_ASAP7_75t_R _32286_ (.A1(_09461_),
    .A2(_11675_),
    .B1(_12234_),
    .B2(_01944_),
    .C(_12238_),
    .Y(_12239_));
 INVx1_ASAP7_75t_R _32287_ (.A(_12239_),
    .Y(_04270_));
 NOR2x2_ASAP7_75t_R _32288_ (.A(_01718_),
    .B(_06301_),
    .Y(_12240_));
 TAPCELL_ASAP7_75t_R PHY_138 ();
 AND3x1_ASAP7_75t_R _32290_ (.A(net3526),
    .B(_11406_),
    .C(_11414_),
    .Y(_12242_));
 AO21x1_ASAP7_75t_R _32291_ (.A1(_01905_),
    .A2(_12240_),
    .B(_12242_),
    .Y(_12243_));
 TAPCELL_ASAP7_75t_R PHY_137 ();
 NAND2x1_ASAP7_75t_R _32293_ (.A(_11159_),
    .B(_11407_),
    .Y(_12245_));
 OA211x2_ASAP7_75t_R _32294_ (.A1(_09468_),
    .A2(_11407_),
    .B(_12245_),
    .C(_11422_),
    .Y(_12246_));
 OR3x1_ASAP7_75t_R _32295_ (.A(_12234_),
    .B(_12243_),
    .C(_12246_),
    .Y(_12247_));
 OAI21x1_ASAP7_75t_R _32296_ (.A1(_01943_),
    .A2(_12232_),
    .B(_12247_),
    .Y(_04271_));
 INVx1_ASAP7_75t_R _32297_ (.A(_01942_),
    .Y(_12248_));
 TAPCELL_ASAP7_75t_R PHY_136 ();
 TAPCELL_ASAP7_75t_R PHY_135 ();
 TAPCELL_ASAP7_75t_R PHY_134 ();
 TAPCELL_ASAP7_75t_R PHY_133 ();
 AOI22x1_ASAP7_75t_R _32302_ (.A1(_09480_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_01904_),
    .Y(_12253_));
 OA211x2_ASAP7_75t_R _32303_ (.A1(net3544),
    .A2(_11423_),
    .B(_12232_),
    .C(_12253_),
    .Y(_12254_));
 AO21x1_ASAP7_75t_R _32304_ (.A1(_12248_),
    .A2(_12234_),
    .B(_12254_),
    .Y(_04272_));
 INVx1_ASAP7_75t_R _32305_ (.A(_01941_),
    .Y(_12255_));
 AOI22x1_ASAP7_75t_R _32306_ (.A1(_09488_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_01903_),
    .Y(_12256_));
 OA211x2_ASAP7_75t_R _32307_ (.A1(net3379),
    .A2(_11423_),
    .B(_12232_),
    .C(_12256_),
    .Y(_12257_));
 AO21x1_ASAP7_75t_R _32308_ (.A1(_12255_),
    .A2(_12234_),
    .B(_12257_),
    .Y(_04273_));
 TAPCELL_ASAP7_75t_R PHY_132 ();
 TAPCELL_ASAP7_75t_R PHY_131 ();
 TAPCELL_ASAP7_75t_R PHY_130 ();
 INVx1_ASAP7_75t_R _32312_ (.A(_01902_),
    .Y(_12261_));
 AO22x1_ASAP7_75t_R _32313_ (.A1(_09498_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12261_),
    .Y(_12262_));
 AO21x1_ASAP7_75t_R _32314_ (.A1(net3632),
    .A2(_12231_),
    .B(_12262_),
    .Y(_12263_));
 NAND2x1_ASAP7_75t_R _32315_ (.A(_01940_),
    .B(_12234_),
    .Y(_12264_));
 OA21x2_ASAP7_75t_R _32316_ (.A1(_12234_),
    .A2(_12263_),
    .B(_12264_),
    .Y(_04274_));
 INVx1_ASAP7_75t_R _32317_ (.A(_01939_),
    .Y(_12265_));
 INVx1_ASAP7_75t_R _32318_ (.A(_01901_),
    .Y(_12266_));
 AO221x1_ASAP7_75t_R _32319_ (.A1(_09506_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12266_),
    .C(_12234_),
    .Y(_12267_));
 AO21x1_ASAP7_75t_R _32320_ (.A1(_09504_),
    .A2(_12231_),
    .B(_12267_),
    .Y(_12268_));
 OA21x2_ASAP7_75t_R _32321_ (.A1(_12265_),
    .A2(_12232_),
    .B(_12268_),
    .Y(_04275_));
 TAPCELL_ASAP7_75t_R PHY_129 ();
 INVx1_ASAP7_75t_R _32323_ (.A(_01900_),
    .Y(_12270_));
 AO22x1_ASAP7_75t_R _32324_ (.A1(_09514_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12270_),
    .Y(_12271_));
 AO21x1_ASAP7_75t_R _32325_ (.A1(net3615),
    .A2(_12231_),
    .B(_12271_),
    .Y(_12272_));
 NAND2x1_ASAP7_75t_R _32326_ (.A(_01938_),
    .B(_12234_),
    .Y(_12273_));
 OA21x2_ASAP7_75t_R _32327_ (.A1(_12234_),
    .A2(_12272_),
    .B(_12273_),
    .Y(_04276_));
 INVx1_ASAP7_75t_R _32328_ (.A(_01899_),
    .Y(_12274_));
 AO221x1_ASAP7_75t_R _32329_ (.A1(_09520_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12274_),
    .C(_12234_),
    .Y(_12275_));
 AO21x1_ASAP7_75t_R _32330_ (.A1(_09518_),
    .A2(_12231_),
    .B(_12275_),
    .Y(_12276_));
 OA21x2_ASAP7_75t_R _32331_ (.A1(_06381_),
    .A2(_12232_),
    .B(_12276_),
    .Y(_04277_));
 INVx1_ASAP7_75t_R _32332_ (.A(_01898_),
    .Y(_12277_));
 AO22x1_ASAP7_75t_R _32333_ (.A1(_09526_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12277_),
    .Y(_12278_));
 AO21x1_ASAP7_75t_R _32334_ (.A1(_09524_),
    .A2(_12231_),
    .B(_12278_),
    .Y(_12279_));
 NAND2x1_ASAP7_75t_R _32335_ (.A(_01936_),
    .B(_12234_),
    .Y(_12280_));
 OA21x2_ASAP7_75t_R _32336_ (.A1(_12234_),
    .A2(_12279_),
    .B(_12280_),
    .Y(_04278_));
 TAPCELL_ASAP7_75t_R PHY_128 ();
 INVx1_ASAP7_75t_R _32338_ (.A(_01897_),
    .Y(_12282_));
 AO22x1_ASAP7_75t_R _32339_ (.A1(_09533_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12282_),
    .Y(_12283_));
 AO21x1_ASAP7_75t_R _32340_ (.A1(_09531_),
    .A2(_12231_),
    .B(_12283_),
    .Y(_12284_));
 NAND2x1_ASAP7_75t_R _32341_ (.A(_01935_),
    .B(_12234_),
    .Y(_12285_));
 OA21x2_ASAP7_75t_R _32342_ (.A1(_12234_),
    .A2(_12284_),
    .B(_12285_),
    .Y(_04279_));
 INVx1_ASAP7_75t_R _32343_ (.A(_01896_),
    .Y(_12286_));
 AO22x1_ASAP7_75t_R _32344_ (.A1(_09541_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12286_),
    .Y(_12287_));
 AO21x1_ASAP7_75t_R _32345_ (.A1(_09538_),
    .A2(_12231_),
    .B(_12287_),
    .Y(_12288_));
 NAND2x1_ASAP7_75t_R _32346_ (.A(_01934_),
    .B(_12234_),
    .Y(_12289_));
 OA21x2_ASAP7_75t_R _32347_ (.A1(_12234_),
    .A2(_12288_),
    .B(_12289_),
    .Y(_04280_));
 INVx1_ASAP7_75t_R _32348_ (.A(_01933_),
    .Y(_12290_));
 INVx1_ASAP7_75t_R _32349_ (.A(_01895_),
    .Y(_12291_));
 AO221x1_ASAP7_75t_R _32350_ (.A1(_09551_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12291_),
    .C(_12234_),
    .Y(_12292_));
 AO21x1_ASAP7_75t_R _32351_ (.A1(net3673),
    .A2(_12231_),
    .B(_12292_),
    .Y(_12293_));
 OA21x2_ASAP7_75t_R _32352_ (.A1(_12290_),
    .A2(_12232_),
    .B(_12293_),
    .Y(_04281_));
 INVx1_ASAP7_75t_R _32353_ (.A(_01894_),
    .Y(_12294_));
 AO22x1_ASAP7_75t_R _32354_ (.A1(_09560_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12294_),
    .Y(_12295_));
 AO21x1_ASAP7_75t_R _32355_ (.A1(net3707),
    .A2(_12231_),
    .B(_12295_),
    .Y(_12296_));
 NAND2x1_ASAP7_75t_R _32356_ (.A(_01932_),
    .B(_12234_),
    .Y(_12297_));
 OA21x2_ASAP7_75t_R _32357_ (.A1(_12234_),
    .A2(_12296_),
    .B(_12297_),
    .Y(_04282_));
 TAPCELL_ASAP7_75t_R PHY_127 ();
 INVx1_ASAP7_75t_R _32359_ (.A(_01893_),
    .Y(_12299_));
 AO22x1_ASAP7_75t_R _32360_ (.A1(_09569_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12299_),
    .Y(_12300_));
 AO21x1_ASAP7_75t_R _32361_ (.A1(net3541),
    .A2(_12231_),
    .B(_12300_),
    .Y(_12301_));
 NAND2x1_ASAP7_75t_R _32362_ (.A(_01931_),
    .B(_12234_),
    .Y(_12302_));
 OA21x2_ASAP7_75t_R _32363_ (.A1(_12234_),
    .A2(_12301_),
    .B(_12302_),
    .Y(_04283_));
 INVx1_ASAP7_75t_R _32364_ (.A(_01892_),
    .Y(_12303_));
 AO22x1_ASAP7_75t_R _32365_ (.A1(_09580_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12303_),
    .Y(_12304_));
 AO21x1_ASAP7_75t_R _32366_ (.A1(net3747),
    .A2(_12231_),
    .B(_12304_),
    .Y(_12305_));
 NAND2x1_ASAP7_75t_R _32367_ (.A(_01930_),
    .B(_12234_),
    .Y(_12306_));
 OA21x2_ASAP7_75t_R _32368_ (.A1(_12234_),
    .A2(_12305_),
    .B(_12306_),
    .Y(_04284_));
 INVx1_ASAP7_75t_R _32369_ (.A(_01891_),
    .Y(_12307_));
 AO22x1_ASAP7_75t_R _32370_ (.A1(_09587_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12307_),
    .Y(_12308_));
 AO21x1_ASAP7_75t_R _32371_ (.A1(net3604),
    .A2(_12231_),
    .B(_12308_),
    .Y(_12309_));
 NAND2x1_ASAP7_75t_R _32372_ (.A(_01929_),
    .B(_12234_),
    .Y(_12310_));
 OA21x2_ASAP7_75t_R _32373_ (.A1(_12234_),
    .A2(_12309_),
    .B(_12310_),
    .Y(_04285_));
 INVx1_ASAP7_75t_R _32374_ (.A(_01928_),
    .Y(_12311_));
 INVx1_ASAP7_75t_R _32375_ (.A(_01890_),
    .Y(_12312_));
 AO221x1_ASAP7_75t_R _32376_ (.A1(_09595_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12312_),
    .C(_12234_),
    .Y(_12313_));
 AO21x1_ASAP7_75t_R _32377_ (.A1(net3660),
    .A2(_12231_),
    .B(_12313_),
    .Y(_12314_));
 OA21x2_ASAP7_75t_R _32378_ (.A1(_12311_),
    .A2(_12232_),
    .B(_12314_),
    .Y(_04286_));
 INVx1_ASAP7_75t_R _32379_ (.A(_01889_),
    .Y(_12315_));
 AOI22x1_ASAP7_75t_R _32380_ (.A1(_09603_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12315_),
    .Y(_12316_));
 OA211x2_ASAP7_75t_R _32381_ (.A1(net3571),
    .A2(_11423_),
    .B(_12232_),
    .C(_12316_),
    .Y(_12317_));
 AOI21x1_ASAP7_75t_R _32382_ (.A1(_01927_),
    .A2(_12234_),
    .B(_12317_),
    .Y(_04287_));
 INVx1_ASAP7_75t_R _32383_ (.A(_01888_),
    .Y(_12318_));
 AO22x1_ASAP7_75t_R _32384_ (.A1(_09610_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12318_),
    .Y(_12319_));
 AO21x1_ASAP7_75t_R _32385_ (.A1(net3711),
    .A2(_12231_),
    .B(_12319_),
    .Y(_12320_));
 NAND2x1_ASAP7_75t_R _32386_ (.A(_01926_),
    .B(_12234_),
    .Y(_12321_));
 OA21x2_ASAP7_75t_R _32387_ (.A1(_12234_),
    .A2(_12320_),
    .B(_12321_),
    .Y(_04288_));
 INVx1_ASAP7_75t_R _32388_ (.A(_01887_),
    .Y(_12322_));
 AOI22x1_ASAP7_75t_R _32389_ (.A1(_09618_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12322_),
    .Y(_12323_));
 OA211x2_ASAP7_75t_R _32390_ (.A1(net3682),
    .A2(_11423_),
    .B(_12232_),
    .C(_12323_),
    .Y(_12324_));
 AOI21x1_ASAP7_75t_R _32391_ (.A1(_01925_),
    .A2(_12234_),
    .B(_12324_),
    .Y(_04289_));
 INVx1_ASAP7_75t_R _32392_ (.A(_01924_),
    .Y(_12325_));
 INVx1_ASAP7_75t_R _32393_ (.A(_01886_),
    .Y(_12326_));
 AO221x1_ASAP7_75t_R _32394_ (.A1(_09626_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12326_),
    .C(_12234_),
    .Y(_12327_));
 AO21x1_ASAP7_75t_R _32395_ (.A1(_09623_),
    .A2(_12231_),
    .B(_12327_),
    .Y(_12328_));
 OA21x2_ASAP7_75t_R _32396_ (.A1(_12325_),
    .A2(_12232_),
    .B(_12328_),
    .Y(_04290_));
 INVx1_ASAP7_75t_R _32397_ (.A(_01885_),
    .Y(_12329_));
 AO22x1_ASAP7_75t_R _32398_ (.A1(_09633_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12329_),
    .Y(_12330_));
 AO21x1_ASAP7_75t_R _32399_ (.A1(_09631_),
    .A2(_12231_),
    .B(_12330_),
    .Y(_12331_));
 NAND2x1_ASAP7_75t_R _32400_ (.A(_01923_),
    .B(_12234_),
    .Y(_12332_));
 OA21x2_ASAP7_75t_R _32401_ (.A1(_12234_),
    .A2(_12331_),
    .B(_12332_),
    .Y(_04291_));
 INVx1_ASAP7_75t_R _32402_ (.A(_01884_),
    .Y(_12333_));
 AOI22x1_ASAP7_75t_R _32403_ (.A1(_09640_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12333_),
    .Y(_12334_));
 OA211x2_ASAP7_75t_R _32404_ (.A1(net3599),
    .A2(_11423_),
    .B(_12232_),
    .C(_12334_),
    .Y(_12335_));
 AOI21x1_ASAP7_75t_R _32405_ (.A1(_01922_),
    .A2(_12234_),
    .B(_12335_),
    .Y(_04292_));
 OAI22x1_ASAP7_75t_R _32406_ (.A1(_09649_),
    .A2(_11408_),
    .B1(_11414_),
    .B2(_01883_),
    .Y(_12336_));
 AO21x1_ASAP7_75t_R _32407_ (.A1(_09647_),
    .A2(_12231_),
    .B(_12336_),
    .Y(_12337_));
 NAND2x1_ASAP7_75t_R _32408_ (.A(_01921_),
    .B(_12234_),
    .Y(_12338_));
 OA21x2_ASAP7_75t_R _32409_ (.A1(_12234_),
    .A2(_12337_),
    .B(_12338_),
    .Y(_04293_));
 INVx1_ASAP7_75t_R _32410_ (.A(_01882_),
    .Y(_12339_));
 AO22x1_ASAP7_75t_R _32411_ (.A1(_09656_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12339_),
    .Y(_12340_));
 AO21x1_ASAP7_75t_R _32412_ (.A1(net3639),
    .A2(_12231_),
    .B(_12340_),
    .Y(_12341_));
 NAND2x1_ASAP7_75t_R _32413_ (.A(_01920_),
    .B(_12234_),
    .Y(_12342_));
 OA21x2_ASAP7_75t_R _32414_ (.A1(_12234_),
    .A2(_12341_),
    .B(_12342_),
    .Y(_04294_));
 INVx1_ASAP7_75t_R _32415_ (.A(_01881_),
    .Y(_12343_));
 AOI22x1_ASAP7_75t_R _32416_ (.A1(_09664_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12343_),
    .Y(_12344_));
 OA211x2_ASAP7_75t_R _32417_ (.A1(_09661_),
    .A2(_11423_),
    .B(_12232_),
    .C(_12344_),
    .Y(_12345_));
 AOI21x1_ASAP7_75t_R _32418_ (.A1(_01919_),
    .A2(_12234_),
    .B(_12345_),
    .Y(_04295_));
 INVx1_ASAP7_75t_R _32419_ (.A(_01880_),
    .Y(_12346_));
 AO22x1_ASAP7_75t_R _32420_ (.A1(_09671_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12346_),
    .Y(_12347_));
 AO21x1_ASAP7_75t_R _32421_ (.A1(net3594),
    .A2(_12231_),
    .B(_12347_),
    .Y(_12348_));
 NAND2x1_ASAP7_75t_R _32422_ (.A(_01918_),
    .B(_12234_),
    .Y(_12349_));
 OA21x2_ASAP7_75t_R _32423_ (.A1(_12234_),
    .A2(_12348_),
    .B(_12349_),
    .Y(_04296_));
 INVx1_ASAP7_75t_R _32424_ (.A(_01879_),
    .Y(_12350_));
 AO22x1_ASAP7_75t_R _32425_ (.A1(_09678_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12350_),
    .Y(_12351_));
 AO21x1_ASAP7_75t_R _32426_ (.A1(_09676_),
    .A2(_12231_),
    .B(_12351_),
    .Y(_12352_));
 NAND2x1_ASAP7_75t_R _32427_ (.A(_01917_),
    .B(_12234_),
    .Y(_12353_));
 OA21x2_ASAP7_75t_R _32428_ (.A1(_12234_),
    .A2(_12352_),
    .B(_12353_),
    .Y(_04297_));
 INVx1_ASAP7_75t_R _32429_ (.A(_01878_),
    .Y(_12354_));
 AO22x1_ASAP7_75t_R _32430_ (.A1(_09686_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12354_),
    .Y(_12355_));
 AO21x1_ASAP7_75t_R _32431_ (.A1(_09683_),
    .A2(_12231_),
    .B(_12355_),
    .Y(_12356_));
 NAND2x1_ASAP7_75t_R _32432_ (.A(_01916_),
    .B(_12234_),
    .Y(_12357_));
 OA21x2_ASAP7_75t_R _32433_ (.A1(_12234_),
    .A2(_12356_),
    .B(_12357_),
    .Y(_04298_));
 INVx1_ASAP7_75t_R _32434_ (.A(_01915_),
    .Y(_12358_));
 INVx1_ASAP7_75t_R _32435_ (.A(_01877_),
    .Y(_12359_));
 AO221x1_ASAP7_75t_R _32436_ (.A1(_09694_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_12359_),
    .C(_12234_),
    .Y(_12360_));
 AO21x1_ASAP7_75t_R _32437_ (.A1(_09691_),
    .A2(_12231_),
    .B(_12360_),
    .Y(_12361_));
 OA21x2_ASAP7_75t_R _32438_ (.A1(_12358_),
    .A2(_12232_),
    .B(_12361_),
    .Y(_04299_));
 NOR2x1_ASAP7_75t_R _32439_ (.A(_09698_),
    .B(_11423_),
    .Y(_12362_));
 AO221x1_ASAP7_75t_R _32440_ (.A1(_09701_),
    .A2(_11675_),
    .B1(_12240_),
    .B2(_01876_),
    .C(_12234_),
    .Y(_12363_));
 OAI22x1_ASAP7_75t_R _32441_ (.A1(_01914_),
    .A2(_12232_),
    .B1(_12362_),
    .B2(_12363_),
    .Y(_04300_));
 AO21x2_ASAP7_75t_R _32442_ (.A1(_06965_),
    .A2(_11327_),
    .B(_11423_),
    .Y(_12364_));
 INVx4_ASAP7_75t_R _32443_ (.A(_12364_),
    .Y(_12365_));
 AND5x1_ASAP7_75t_R _32444_ (.A(_01740_),
    .B(_01741_),
    .C(_06612_),
    .D(_14813_),
    .E(_06372_),
    .Y(_12366_));
 AND2x2_ASAP7_75t_R _32445_ (.A(net375),
    .B(_05732_),
    .Y(_12367_));
 AO21x1_ASAP7_75t_R _32446_ (.A1(net323),
    .A2(_06210_),
    .B(_12367_),
    .Y(_12368_));
 AND5x1_ASAP7_75t_R _32447_ (.A(net2277),
    .B(_01312_),
    .C(_01721_),
    .D(_12366_),
    .E(_12368_),
    .Y(_12369_));
 NOR2x1_ASAP7_75t_R _32448_ (.A(_06211_),
    .B(_12369_),
    .Y(_12370_));
 AO21x1_ASAP7_75t_R _32449_ (.A1(_11902_),
    .A2(_12370_),
    .B(_06319_),
    .Y(_12371_));
 AO21x1_ASAP7_75t_R _32450_ (.A1(net3390),
    .A2(_12371_),
    .B(_11408_),
    .Y(_12372_));
 OA21x2_ASAP7_75t_R _32451_ (.A1(_02104_),
    .A2(_11414_),
    .B(_12372_),
    .Y(_12373_));
 OA211x2_ASAP7_75t_R _32452_ (.A1(net3517),
    .A2(_11423_),
    .B(_12364_),
    .C(_12373_),
    .Y(_12374_));
 AOI21x1_ASAP7_75t_R _32453_ (.A1(_01913_),
    .A2(_12365_),
    .B(net3518),
    .Y(_04301_));
 AO21x1_ASAP7_75t_R _32454_ (.A1(net2277),
    .A2(_12366_),
    .B(_01725_),
    .Y(_12375_));
 NAND2x1_ASAP7_75t_R _32455_ (.A(_01312_),
    .B(_12375_),
    .Y(_12376_));
 OA211x2_ASAP7_75t_R _32456_ (.A1(_12369_),
    .A2(_12376_),
    .B(_06205_),
    .C(_06385_),
    .Y(_12377_));
 OA211x2_ASAP7_75t_R _32457_ (.A1(net3509),
    .A2(_12377_),
    .B(_06932_),
    .C(_01311_),
    .Y(_12378_));
 AO21x1_ASAP7_75t_R _32458_ (.A1(_09452_),
    .A2(_11407_),
    .B(_12378_),
    .Y(_12379_));
 AND3x1_ASAP7_75t_R _32459_ (.A(_09452_),
    .B(_11406_),
    .C(_11414_),
    .Y(_12380_));
 AO21x1_ASAP7_75t_R _32460_ (.A1(_11683_),
    .A2(_12240_),
    .B(_12380_),
    .Y(_12381_));
 AO21x1_ASAP7_75t_R _32461_ (.A1(_11422_),
    .A2(_12379_),
    .B(_12381_),
    .Y(_12382_));
 NAND2x1_ASAP7_75t_R _32462_ (.A(_01912_),
    .B(_12365_),
    .Y(_12383_));
 OA21x2_ASAP7_75t_R _32463_ (.A1(_12365_),
    .A2(_12382_),
    .B(_12383_),
    .Y(_04302_));
 AO21x1_ASAP7_75t_R _32464_ (.A1(_02102_),
    .A2(_12240_),
    .B(_12242_),
    .Y(_12384_));
 OR4x1_ASAP7_75t_R _32465_ (.A(_06225_),
    .B(_01715_),
    .C(_01716_),
    .D(_14791_),
    .Y(_12385_));
 OA22x2_ASAP7_75t_R _32466_ (.A1(_06271_),
    .A2(net3502),
    .B1(_11902_),
    .B2(_12385_),
    .Y(_12386_));
 OA211x2_ASAP7_75t_R _32467_ (.A1(_11407_),
    .A2(_12386_),
    .B(_12245_),
    .C(_11422_),
    .Y(_12387_));
 OR3x1_ASAP7_75t_R _32468_ (.A(_12365_),
    .B(_12384_),
    .C(_12387_),
    .Y(_12388_));
 OAI21x1_ASAP7_75t_R _32469_ (.A1(_01911_),
    .A2(_12364_),
    .B(_12388_),
    .Y(_04303_));
 NAND2x1_ASAP7_75t_R _32470_ (.A(_13390_),
    .B(_06385_),
    .Y(_12389_));
 OA211x2_ASAP7_75t_R _32471_ (.A1(_06889_),
    .A2(_12389_),
    .B(_11675_),
    .C(_06350_),
    .Y(_12390_));
 AOI21x1_ASAP7_75t_R _32472_ (.A1(_02101_),
    .A2(_12240_),
    .B(_12390_),
    .Y(_12391_));
 OA211x2_ASAP7_75t_R _32473_ (.A1(net3544),
    .A2(_11423_),
    .B(_12364_),
    .C(_12391_),
    .Y(_12392_));
 AO21x1_ASAP7_75t_R _32474_ (.A1(_11689_),
    .A2(_12365_),
    .B(_12392_),
    .Y(_04304_));
 OA21x2_ASAP7_75t_R _32475_ (.A1(_02100_),
    .A2(_11414_),
    .B(net3413),
    .Y(_12393_));
 OA211x2_ASAP7_75t_R _32476_ (.A1(net3378),
    .A2(_11423_),
    .B(_12364_),
    .C(net3414),
    .Y(_12394_));
 AOI21x1_ASAP7_75t_R _32477_ (.A1(_01909_),
    .A2(_12365_),
    .B(_12394_),
    .Y(_04305_));
 NAND2x1_ASAP7_75t_R _32478_ (.A(_09698_),
    .B(_12231_),
    .Y(_12395_));
 OA211x2_ASAP7_75t_R _32479_ (.A1(_02099_),
    .A2(_11414_),
    .B(_12364_),
    .C(net3211),
    .Y(_12396_));
 AOI22x1_ASAP7_75t_R _32480_ (.A1(_01908_),
    .A2(_12365_),
    .B1(_12395_),
    .B2(_12396_),
    .Y(_04306_));
 AND2x2_ASAP7_75t_R _32481_ (.A(_01945_),
    .B(_11675_),
    .Y(_12397_));
 AOI21x1_ASAP7_75t_R _32482_ (.A1(_01907_),
    .A2(_11408_),
    .B(_12397_),
    .Y(_04307_));
 AND2x2_ASAP7_75t_R _32483_ (.A(_01944_),
    .B(_11675_),
    .Y(_12398_));
 AOI21x1_ASAP7_75t_R _32484_ (.A1(_01906_),
    .A2(_11408_),
    .B(_12398_),
    .Y(_04308_));
 NAND2x1_ASAP7_75t_R _32485_ (.A(_01905_),
    .B(_11408_),
    .Y(_12399_));
 OA21x2_ASAP7_75t_R _32486_ (.A1(_07449_),
    .A2(_11408_),
    .B(_12399_),
    .Y(_04309_));
 NAND2x1_ASAP7_75t_R _32487_ (.A(_01904_),
    .B(_11408_),
    .Y(_12400_));
 OA21x2_ASAP7_75t_R _32488_ (.A1(_12248_),
    .A2(_11408_),
    .B(_12400_),
    .Y(_04310_));
 NAND2x1_ASAP7_75t_R _32489_ (.A(_01903_),
    .B(_11408_),
    .Y(_12401_));
 OA21x2_ASAP7_75t_R _32490_ (.A1(_12255_),
    .A2(_11408_),
    .B(_12401_),
    .Y(_04311_));
 NAND2x1_ASAP7_75t_R _32491_ (.A(_01940_),
    .B(_11675_),
    .Y(_12402_));
 OA21x2_ASAP7_75t_R _32492_ (.A1(_12261_),
    .A2(_11675_),
    .B(_12402_),
    .Y(_04312_));
 OR3x1_ASAP7_75t_R _32493_ (.A(_12265_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12403_));
 OA21x2_ASAP7_75t_R _32494_ (.A1(_12266_),
    .A2(_11675_),
    .B(_12403_),
    .Y(_04313_));
 NAND2x1_ASAP7_75t_R _32495_ (.A(_01938_),
    .B(_11675_),
    .Y(_12404_));
 OA21x2_ASAP7_75t_R _32496_ (.A1(_12270_),
    .A2(_11675_),
    .B(_12404_),
    .Y(_04314_));
 OR3x1_ASAP7_75t_R _32497_ (.A(_06381_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12405_));
 OA21x2_ASAP7_75t_R _32498_ (.A1(_12274_),
    .A2(_11675_),
    .B(_12405_),
    .Y(_04315_));
 NAND2x1_ASAP7_75t_R _32499_ (.A(_01936_),
    .B(_11675_),
    .Y(_12406_));
 OA21x2_ASAP7_75t_R _32500_ (.A1(_12277_),
    .A2(_11675_),
    .B(_12406_),
    .Y(_04316_));
 TAPCELL_ASAP7_75t_R PHY_126 ();
 NAND2x1_ASAP7_75t_R _32502_ (.A(_01935_),
    .B(_11675_),
    .Y(_12408_));
 OA21x2_ASAP7_75t_R _32503_ (.A1(_12282_),
    .A2(_11675_),
    .B(_12408_),
    .Y(_04317_));
 NAND2x1_ASAP7_75t_R _32504_ (.A(_01934_),
    .B(_11675_),
    .Y(_12409_));
 OA21x2_ASAP7_75t_R _32505_ (.A1(_12286_),
    .A2(_11675_),
    .B(_12409_),
    .Y(_04318_));
 OR3x1_ASAP7_75t_R _32506_ (.A(_12290_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12410_));
 OA21x2_ASAP7_75t_R _32507_ (.A1(_12291_),
    .A2(_11675_),
    .B(_12410_),
    .Y(_04319_));
 NAND2x1_ASAP7_75t_R _32508_ (.A(_01932_),
    .B(_11675_),
    .Y(_12411_));
 OA21x2_ASAP7_75t_R _32509_ (.A1(_12294_),
    .A2(_11675_),
    .B(_12411_),
    .Y(_04320_));
 TAPCELL_ASAP7_75t_R PHY_125 ();
 NAND2x1_ASAP7_75t_R _32511_ (.A(_01931_),
    .B(_11675_),
    .Y(_12413_));
 OA21x2_ASAP7_75t_R _32512_ (.A1(_12299_),
    .A2(_11675_),
    .B(_12413_),
    .Y(_04321_));
 NAND2x1_ASAP7_75t_R _32513_ (.A(_01930_),
    .B(_11675_),
    .Y(_12414_));
 OA21x2_ASAP7_75t_R _32514_ (.A1(_12303_),
    .A2(_11675_),
    .B(_12414_),
    .Y(_04322_));
 NAND2x1_ASAP7_75t_R _32515_ (.A(_01929_),
    .B(_11675_),
    .Y(_12415_));
 OA21x2_ASAP7_75t_R _32516_ (.A1(_12307_),
    .A2(_11675_),
    .B(_12415_),
    .Y(_04323_));
 OR3x1_ASAP7_75t_R _32517_ (.A(_12311_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12416_));
 OA21x2_ASAP7_75t_R _32518_ (.A1(_12312_),
    .A2(_11675_),
    .B(_12416_),
    .Y(_04324_));
 NAND2x1_ASAP7_75t_R _32519_ (.A(_01927_),
    .B(_11675_),
    .Y(_12417_));
 OA21x2_ASAP7_75t_R _32520_ (.A1(_12315_),
    .A2(_11675_),
    .B(_12417_),
    .Y(_04325_));
 NAND2x1_ASAP7_75t_R _32521_ (.A(_01926_),
    .B(_11675_),
    .Y(_12418_));
 OA21x2_ASAP7_75t_R _32522_ (.A1(_12318_),
    .A2(_11675_),
    .B(_12418_),
    .Y(_04326_));
 NAND2x1_ASAP7_75t_R _32523_ (.A(_01925_),
    .B(_11675_),
    .Y(_12419_));
 OA21x2_ASAP7_75t_R _32524_ (.A1(_12322_),
    .A2(_11675_),
    .B(_12419_),
    .Y(_04327_));
 OR3x1_ASAP7_75t_R _32525_ (.A(_12325_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12420_));
 OA21x2_ASAP7_75t_R _32526_ (.A1(_12326_),
    .A2(_11675_),
    .B(_12420_),
    .Y(_04328_));
 NAND2x1_ASAP7_75t_R _32527_ (.A(_01923_),
    .B(_11675_),
    .Y(_12421_));
 OA21x2_ASAP7_75t_R _32528_ (.A1(_12329_),
    .A2(_11675_),
    .B(_12421_),
    .Y(_04329_));
 NAND2x1_ASAP7_75t_R _32529_ (.A(_01922_),
    .B(_11675_),
    .Y(_12422_));
 OA21x2_ASAP7_75t_R _32530_ (.A1(_12333_),
    .A2(_11675_),
    .B(_12422_),
    .Y(_04330_));
 AND2x2_ASAP7_75t_R _32531_ (.A(_01921_),
    .B(_11675_),
    .Y(_12423_));
 AOI21x1_ASAP7_75t_R _32532_ (.A1(_01883_),
    .A2(_11408_),
    .B(_12423_),
    .Y(_04331_));
 NAND2x1_ASAP7_75t_R _32533_ (.A(_01920_),
    .B(_11675_),
    .Y(_12424_));
 OA21x2_ASAP7_75t_R _32534_ (.A1(_12339_),
    .A2(_11675_),
    .B(_12424_),
    .Y(_04332_));
 NAND2x1_ASAP7_75t_R _32535_ (.A(_01919_),
    .B(_11675_),
    .Y(_12425_));
 OA21x2_ASAP7_75t_R _32536_ (.A1(_12343_),
    .A2(_11675_),
    .B(_12425_),
    .Y(_04333_));
 NAND2x1_ASAP7_75t_R _32537_ (.A(_01918_),
    .B(_11675_),
    .Y(_12426_));
 OA21x2_ASAP7_75t_R _32538_ (.A1(_12346_),
    .A2(_11675_),
    .B(_12426_),
    .Y(_04334_));
 NAND2x1_ASAP7_75t_R _32539_ (.A(_01917_),
    .B(_11675_),
    .Y(_12427_));
 OA21x2_ASAP7_75t_R _32540_ (.A1(_12350_),
    .A2(_11675_),
    .B(_12427_),
    .Y(_04335_));
 NAND2x1_ASAP7_75t_R _32541_ (.A(_01916_),
    .B(_11675_),
    .Y(_12428_));
 OA21x2_ASAP7_75t_R _32542_ (.A1(_12354_),
    .A2(_11675_),
    .B(_12428_),
    .Y(_04336_));
 OR3x1_ASAP7_75t_R _32543_ (.A(_12358_),
    .B(_11406_),
    .C(_11407_),
    .Y(_12429_));
 OA21x2_ASAP7_75t_R _32544_ (.A1(_12359_),
    .A2(_11675_),
    .B(_12429_),
    .Y(_04337_));
 AND2x2_ASAP7_75t_R _32545_ (.A(_01914_),
    .B(_11675_),
    .Y(_12430_));
 AOI21x1_ASAP7_75t_R _32546_ (.A1(_01876_),
    .A2(_11408_),
    .B(_12430_),
    .Y(_04338_));
 AND4x2_ASAP7_75t_R _32547_ (.A(net302),
    .B(_14358_),
    .C(_05693_),
    .D(_11081_),
    .Y(_12431_));
 NAND2x1_ASAP7_75t_R _32548_ (.A(_12431_),
    .B(_11096_),
    .Y(_12432_));
 AO21x1_ASAP7_75t_R _32549_ (.A1(_12431_),
    .A2(_11096_),
    .B(_11103_),
    .Y(_12433_));
 OA21x2_ASAP7_75t_R _32550_ (.A1(_11262_),
    .A2(_12432_),
    .B(_12433_),
    .Y(_04339_));
 NAND2x1_ASAP7_75t_R _32551_ (.A(_01315_),
    .B(_12432_),
    .Y(_12434_));
 OA21x2_ASAP7_75t_R _32552_ (.A1(_11159_),
    .A2(_12432_),
    .B(_12434_),
    .Y(_04340_));
 NAND2x1_ASAP7_75t_R _32553_ (.A(_01727_),
    .B(_05777_),
    .Y(_12435_));
 OA21x2_ASAP7_75t_R _32554_ (.A1(_13775_),
    .A2(_05777_),
    .B(_12435_),
    .Y(_04343_));
 NAND2x1_ASAP7_75t_R _32555_ (.A(_00284_),
    .B(_05777_),
    .Y(_12436_));
 OA21x2_ASAP7_75t_R _32556_ (.A1(_05776_),
    .A2(_05777_),
    .B(_12436_),
    .Y(_04344_));
 NAND2x1_ASAP7_75t_R _32557_ (.A(_01728_),
    .B(_05777_),
    .Y(_12437_));
 OA21x2_ASAP7_75t_R _32558_ (.A1(_05782_),
    .A2(_05777_),
    .B(_12437_),
    .Y(_04345_));
 AND3x4_ASAP7_75t_R _32559_ (.A(net3055),
    .B(_01316_),
    .C(_01609_),
    .Y(_12438_));
 NAND2x2_ASAP7_75t_R _32560_ (.A(_09313_),
    .B(_12438_),
    .Y(_12439_));
 TAPCELL_ASAP7_75t_R PHY_124 ();
 TAPCELL_ASAP7_75t_R PHY_123 ();
 NAND2x1_ASAP7_75t_R _32563_ (.A(_01871_),
    .B(_12439_),
    .Y(_12442_));
 OA21x2_ASAP7_75t_R _32564_ (.A1(net3817),
    .A2(_12439_),
    .B(_12442_),
    .Y(_04346_));
 TAPCELL_ASAP7_75t_R PHY_122 ();
 TAPCELL_ASAP7_75t_R PHY_121 ();
 AO21x1_ASAP7_75t_R _32567_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07258_),
    .Y(_12445_));
 OA21x2_ASAP7_75t_R _32568_ (.A1(net3871),
    .A2(_12439_),
    .B(_12445_),
    .Y(_04347_));
 AO21x1_ASAP7_75t_R _32569_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07466_),
    .Y(_12446_));
 OA21x2_ASAP7_75t_R _32570_ (.A1(net3823),
    .A2(_12439_),
    .B(_12446_),
    .Y(_04348_));
 NAND2x1_ASAP7_75t_R _32571_ (.A(_01868_),
    .B(_12439_),
    .Y(_12447_));
 OA21x2_ASAP7_75t_R _32572_ (.A1(net3877),
    .A2(_12439_),
    .B(_12447_),
    .Y(_04349_));
 AO21x1_ASAP7_75t_R _32573_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07602_),
    .Y(_12448_));
 OA21x2_ASAP7_75t_R _32574_ (.A1(net3805),
    .A2(_12439_),
    .B(_12448_),
    .Y(_04350_));
 AO21x1_ASAP7_75t_R _32575_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07657_),
    .Y(_12449_));
 OA21x2_ASAP7_75t_R _32576_ (.A1(net3919),
    .A2(_12439_),
    .B(_12449_),
    .Y(_04351_));
 NAND2x1_ASAP7_75t_R _32577_ (.A(_01865_),
    .B(_12439_),
    .Y(_12450_));
 OA21x2_ASAP7_75t_R _32578_ (.A1(net3829),
    .A2(_12439_),
    .B(_12450_),
    .Y(_04352_));
 AO21x1_ASAP7_75t_R _32579_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07754_),
    .Y(_12451_));
 OA21x2_ASAP7_75t_R _32580_ (.A1(net3889),
    .A2(_12439_),
    .B(_12451_),
    .Y(_04353_));
 AO21x1_ASAP7_75t_R _32581_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07035_),
    .Y(_12452_));
 OA21x2_ASAP7_75t_R _32582_ (.A1(net3859),
    .A2(_12439_),
    .B(_12452_),
    .Y(_04354_));
 AO21x1_ASAP7_75t_R _32583_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07257_),
    .Y(_12453_));
 OA21x2_ASAP7_75t_R _32584_ (.A1(net3895),
    .A2(_12439_),
    .B(_12453_),
    .Y(_04355_));
 TAPCELL_ASAP7_75t_R PHY_120 ();
 AO21x1_ASAP7_75t_R _32586_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07465_),
    .Y(_12455_));
 OA21x2_ASAP7_75t_R _32587_ (.A1(net3847),
    .A2(_12439_),
    .B(_12455_),
    .Y(_04356_));
 AO21x1_ASAP7_75t_R _32588_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07545_),
    .Y(_12456_));
 OA21x2_ASAP7_75t_R _32589_ (.A1(net3901),
    .A2(_12439_),
    .B(_12456_),
    .Y(_04357_));
 AO21x1_ASAP7_75t_R _32590_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07601_),
    .Y(_12457_));
 OA21x2_ASAP7_75t_R _32591_ (.A1(net3927),
    .A2(_12439_),
    .B(_12457_),
    .Y(_04358_));
 AO21x1_ASAP7_75t_R _32592_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07656_),
    .Y(_12458_));
 OA21x2_ASAP7_75t_R _32593_ (.A1(net3853),
    .A2(_12439_),
    .B(_12458_),
    .Y(_04359_));
 AO21x1_ASAP7_75t_R _32594_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07666_),
    .Y(_12459_));
 OA21x2_ASAP7_75t_R _32595_ (.A1(net3883),
    .A2(_12439_),
    .B(_12459_),
    .Y(_04360_));
 AO21x1_ASAP7_75t_R _32596_ (.A1(_09313_),
    .A2(_12438_),
    .B(_07753_),
    .Y(_12460_));
 OA21x2_ASAP7_75t_R _32597_ (.A1(net3935),
    .A2(_12439_),
    .B(_12460_),
    .Y(_04361_));
 NAND2x1_ASAP7_75t_R _32598_ (.A(_01855_),
    .B(_12439_),
    .Y(_12461_));
 OA21x2_ASAP7_75t_R _32599_ (.A1(net3944),
    .A2(_12439_),
    .B(_12461_),
    .Y(_04362_));
 NAND2x1_ASAP7_75t_R _32600_ (.A(_01854_),
    .B(_12439_),
    .Y(_12462_));
 OA21x2_ASAP7_75t_R _32601_ (.A1(net3835),
    .A2(_12439_),
    .B(_12462_),
    .Y(_04363_));
 NAND2x1_ASAP7_75t_R _32602_ (.A(_01853_),
    .B(_12439_),
    .Y(_12463_));
 OA21x2_ASAP7_75t_R _32603_ (.A1(net3799),
    .A2(_12439_),
    .B(_12463_),
    .Y(_04364_));
 NAND2x1_ASAP7_75t_R _32604_ (.A(_01852_),
    .B(_12439_),
    .Y(_12464_));
 OA21x2_ASAP7_75t_R _32605_ (.A1(net3841),
    .A2(_12439_),
    .B(_12464_),
    .Y(_04365_));
 NAND2x1_ASAP7_75t_R _32606_ (.A(_01851_),
    .B(_12439_),
    .Y(_12465_));
 OA21x2_ASAP7_75t_R _32607_ (.A1(net3910),
    .A2(_12439_),
    .B(_12465_),
    .Y(_04366_));
 AO21x1_ASAP7_75t_R _32608_ (.A1(_09313_),
    .A2(_12438_),
    .B(_08021_),
    .Y(_12466_));
 OA21x2_ASAP7_75t_R _32609_ (.A1(net3778),
    .A2(_12439_),
    .B(_12466_),
    .Y(_04367_));
 NAND2x1_ASAP7_75t_R _32610_ (.A(_01849_),
    .B(_12439_),
    .Y(_12467_));
 OA21x2_ASAP7_75t_R _32611_ (.A1(net3811),
    .A2(_12439_),
    .B(_12467_),
    .Y(_04368_));
 AO21x1_ASAP7_75t_R _32612_ (.A1(_09313_),
    .A2(_12438_),
    .B(_08402_),
    .Y(_12468_));
 OA21x2_ASAP7_75t_R _32613_ (.A1(net3865),
    .A2(_12439_),
    .B(_12468_),
    .Y(_04369_));
 AND3x1_ASAP7_75t_R _32614_ (.A(_00240_),
    .B(_00239_),
    .C(_06727_),
    .Y(_12469_));
 OR3x1_ASAP7_75t_R _32615_ (.A(_00240_),
    .B(_06734_),
    .C(_06678_),
    .Y(_12470_));
 INVx1_ASAP7_75t_R _32616_ (.A(_12470_),
    .Y(_12471_));
 AND3x1_ASAP7_75t_R _32617_ (.A(_06618_),
    .B(_06723_),
    .C(_12471_),
    .Y(_12472_));
 AO21x2_ASAP7_75t_R _32618_ (.A1(_06724_),
    .A2(_12469_),
    .B(_12472_),
    .Y(_12473_));
 TAPCELL_ASAP7_75t_R PHY_119 ();
 NAND2x2_ASAP7_75t_R _32620_ (.A(_00240_),
    .B(_06727_),
    .Y(_12475_));
 OA21x2_ASAP7_75t_R _32621_ (.A1(_00240_),
    .A2(_06678_),
    .B(_00239_),
    .Y(_12476_));
 AND3x1_ASAP7_75t_R _32622_ (.A(_06618_),
    .B(_06723_),
    .C(_12476_),
    .Y(_12477_));
 AO21x2_ASAP7_75t_R _32623_ (.A1(_06724_),
    .A2(_12475_),
    .B(_12477_),
    .Y(_12478_));
 TAPCELL_ASAP7_75t_R PHY_118 ();
 INVx1_ASAP7_75t_R _32625_ (.A(_01846_),
    .Y(_12480_));
 AOI21x1_ASAP7_75t_R _32626_ (.A1(_06724_),
    .A2(_12475_),
    .B(_00239_),
    .Y(_12481_));
 TAPCELL_ASAP7_75t_R PHY_117 ();
 INVx1_ASAP7_75t_R _32628_ (.A(_01813_),
    .Y(_12483_));
 AO222x2_ASAP7_75t_R _32629_ (.A1(net3002),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12480_),
    .C1(_12481_),
    .C2(_12483_),
    .Y(_04371_));
 INVx1_ASAP7_75t_R _32630_ (.A(_01845_),
    .Y(_12484_));
 INVx1_ASAP7_75t_R _32631_ (.A(_01812_),
    .Y(_12485_));
 AO222x2_ASAP7_75t_R _32632_ (.A1(net3022),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12484_),
    .C1(_12481_),
    .C2(_12485_),
    .Y(_04372_));
 INVx1_ASAP7_75t_R _32633_ (.A(_01844_),
    .Y(_12486_));
 INVx1_ASAP7_75t_R _32634_ (.A(_01811_),
    .Y(_12487_));
 AO222x2_ASAP7_75t_R _32635_ (.A1(net2846),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12486_),
    .C1(net253),
    .C2(_12487_),
    .Y(_04373_));
 INVx1_ASAP7_75t_R _32636_ (.A(_01843_),
    .Y(_12488_));
 INVx1_ASAP7_75t_R _32637_ (.A(_01810_),
    .Y(_12489_));
 AO222x2_ASAP7_75t_R _32638_ (.A1(net2961),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12488_),
    .C1(net253),
    .C2(_12489_),
    .Y(_04374_));
 INVx1_ASAP7_75t_R _32639_ (.A(_01842_),
    .Y(_12490_));
 INVx1_ASAP7_75t_R _32640_ (.A(_01809_),
    .Y(_12491_));
 AO222x2_ASAP7_75t_R _32641_ (.A1(net3122),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12490_),
    .C1(_12481_),
    .C2(_12491_),
    .Y(_04375_));
 INVx1_ASAP7_75t_R _32642_ (.A(_01841_),
    .Y(_12492_));
 INVx1_ASAP7_75t_R _32643_ (.A(_01808_),
    .Y(_12493_));
 AO222x2_ASAP7_75t_R _32644_ (.A1(net2886),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12492_),
    .C1(net253),
    .C2(_12493_),
    .Y(_04376_));
 INVx1_ASAP7_75t_R _32645_ (.A(_01840_),
    .Y(_12494_));
 INVx1_ASAP7_75t_R _32646_ (.A(_01807_),
    .Y(_12495_));
 AO222x2_ASAP7_75t_R _32647_ (.A1(net3077),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12494_),
    .C1(net253),
    .C2(_12495_),
    .Y(_04377_));
 INVx1_ASAP7_75t_R _32648_ (.A(_01839_),
    .Y(_12496_));
 INVx1_ASAP7_75t_R _32649_ (.A(_01806_),
    .Y(_12497_));
 AO222x2_ASAP7_75t_R _32650_ (.A1(net2870),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12496_),
    .C1(net253),
    .C2(_12497_),
    .Y(_04378_));
 INVx1_ASAP7_75t_R _32651_ (.A(_01838_),
    .Y(_12498_));
 INVx1_ASAP7_75t_R _32652_ (.A(_01805_),
    .Y(_12499_));
 AO222x2_ASAP7_75t_R _32653_ (.A1(net2986),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12498_),
    .C1(_12481_),
    .C2(_12499_),
    .Y(_04379_));
 TAPCELL_ASAP7_75t_R PHY_116 ();
 INVx1_ASAP7_75t_R _32655_ (.A(_01837_),
    .Y(_12501_));
 INVx1_ASAP7_75t_R _32656_ (.A(_01804_),
    .Y(_12502_));
 AO222x2_ASAP7_75t_R _32657_ (.A1(net2797),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12501_),
    .C1(net253),
    .C2(_12502_),
    .Y(_04380_));
 TAPCELL_ASAP7_75t_R PHY_115 ();
 INVx1_ASAP7_75t_R _32659_ (.A(_01836_),
    .Y(_12504_));
 TAPCELL_ASAP7_75t_R PHY_114 ();
 INVx1_ASAP7_75t_R _32661_ (.A(_01803_),
    .Y(_12506_));
 AO222x2_ASAP7_75t_R _32662_ (.A1(net2953),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12504_),
    .C1(net253),
    .C2(_12506_),
    .Y(_04381_));
 INVx1_ASAP7_75t_R _32663_ (.A(_01835_),
    .Y(_12507_));
 INVx1_ASAP7_75t_R _32664_ (.A(_01802_),
    .Y(_12508_));
 AO222x2_ASAP7_75t_R _32665_ (.A1(net2838),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12507_),
    .C1(net253),
    .C2(_12508_),
    .Y(_04382_));
 INVx1_ASAP7_75t_R _32666_ (.A(_01834_),
    .Y(_12509_));
 INVx1_ASAP7_75t_R _32667_ (.A(_01801_),
    .Y(_12510_));
 AO222x2_ASAP7_75t_R _32668_ (.A1(net2789),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12509_),
    .C1(net253),
    .C2(_12510_),
    .Y(_04383_));
 INVx1_ASAP7_75t_R _32669_ (.A(_01833_),
    .Y(_12511_));
 INVx1_ASAP7_75t_R _32670_ (.A(_01800_),
    .Y(_12512_));
 AO222x2_ASAP7_75t_R _32671_ (.A1(net2822),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12511_),
    .C1(net253),
    .C2(_12512_),
    .Y(_04384_));
 INVx1_ASAP7_75t_R _32672_ (.A(_01832_),
    .Y(_12513_));
 INVx1_ASAP7_75t_R _32673_ (.A(_01799_),
    .Y(_12514_));
 AO222x2_ASAP7_75t_R _32674_ (.A1(net2830),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12513_),
    .C1(net253),
    .C2(_12514_),
    .Y(_04385_));
 INVx1_ASAP7_75t_R _32675_ (.A(_01831_),
    .Y(_12515_));
 INVx1_ASAP7_75t_R _32676_ (.A(_01798_),
    .Y(_12516_));
 AO222x2_ASAP7_75t_R _32677_ (.A1(net2768),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12515_),
    .C1(net253),
    .C2(_12516_),
    .Y(_04386_));
 INVx1_ASAP7_75t_R _32678_ (.A(_01830_),
    .Y(_12517_));
 INVx1_ASAP7_75t_R _32679_ (.A(_01797_),
    .Y(_12518_));
 AO222x2_ASAP7_75t_R _32680_ (.A1(net2994),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12517_),
    .C1(_12481_),
    .C2(_12518_),
    .Y(_04387_));
 INVx1_ASAP7_75t_R _32681_ (.A(_01829_),
    .Y(_12519_));
 INVx1_ASAP7_75t_R _32682_ (.A(_01796_),
    .Y(_12520_));
 AO222x2_ASAP7_75t_R _32683_ (.A1(net2902),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12519_),
    .C1(net253),
    .C2(_12520_),
    .Y(_04388_));
 INVx1_ASAP7_75t_R _32684_ (.A(_01828_),
    .Y(_12521_));
 INVx1_ASAP7_75t_R _32685_ (.A(_01795_),
    .Y(_12522_));
 AO222x2_ASAP7_75t_R _32686_ (.A1(net2894),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12521_),
    .C1(net253),
    .C2(_12522_),
    .Y(_04389_));
 TAPCELL_ASAP7_75t_R PHY_113 ();
 INVx1_ASAP7_75t_R _32688_ (.A(_01827_),
    .Y(_12524_));
 INVx1_ASAP7_75t_R _32689_ (.A(_01794_),
    .Y(_12525_));
 AO222x2_ASAP7_75t_R _32690_ (.A1(net3010),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12524_),
    .C1(_12481_),
    .C2(_12525_),
    .Y(_04390_));
 TAPCELL_ASAP7_75t_R PHY_112 ();
 INVx1_ASAP7_75t_R _32692_ (.A(_01826_),
    .Y(_12527_));
 TAPCELL_ASAP7_75t_R PHY_111 ();
 INVx1_ASAP7_75t_R _32694_ (.A(_01793_),
    .Y(_12529_));
 AO222x2_ASAP7_75t_R _32695_ (.A1(net3098),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12527_),
    .C1(net253),
    .C2(_12529_),
    .Y(_04391_));
 INVx1_ASAP7_75t_R _32696_ (.A(_01825_),
    .Y(_12530_));
 INVx1_ASAP7_75t_R _32697_ (.A(_01792_),
    .Y(_12531_));
 AO222x2_ASAP7_75t_R _32698_ (.A1(net2878),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12530_),
    .C1(net253),
    .C2(_12531_),
    .Y(_04392_));
 INVx1_ASAP7_75t_R _32699_ (.A(_01824_),
    .Y(_12532_));
 INVx1_ASAP7_75t_R _32700_ (.A(_01791_),
    .Y(_12533_));
 AO222x2_ASAP7_75t_R _32701_ (.A1(net3085),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12532_),
    .C1(net253),
    .C2(_12533_),
    .Y(_04393_));
 INVx1_ASAP7_75t_R _32702_ (.A(_01823_),
    .Y(_12534_));
 INVx1_ASAP7_75t_R _32703_ (.A(_01790_),
    .Y(_12535_));
 AO222x2_ASAP7_75t_R _32704_ (.A1(net2931),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12534_),
    .C1(net253),
    .C2(_12535_),
    .Y(_04394_));
 INVx1_ASAP7_75t_R _32705_ (.A(_01822_),
    .Y(_12536_));
 INVx1_ASAP7_75t_R _32706_ (.A(_01789_),
    .Y(_12537_));
 AO222x2_ASAP7_75t_R _32707_ (.A1(net3114),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12536_),
    .C1(net253),
    .C2(_12537_),
    .Y(_04395_));
 INVx1_ASAP7_75t_R _32708_ (.A(_01821_),
    .Y(_12538_));
 INVx1_ASAP7_75t_R _32709_ (.A(_01788_),
    .Y(_12539_));
 AO222x2_ASAP7_75t_R _32710_ (.A1(net2918),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12538_),
    .C1(net253),
    .C2(_12539_),
    .Y(_04396_));
 INVx1_ASAP7_75t_R _32711_ (.A(_01820_),
    .Y(_12540_));
 INVx1_ASAP7_75t_R _32712_ (.A(_01787_),
    .Y(_12541_));
 AO222x2_ASAP7_75t_R _32713_ (.A1(net2945),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12540_),
    .C1(net253),
    .C2(_12541_),
    .Y(_04397_));
 INVx1_ASAP7_75t_R _32714_ (.A(_01819_),
    .Y(_12542_));
 INVx1_ASAP7_75t_R _32715_ (.A(_01786_),
    .Y(_12543_));
 AO222x2_ASAP7_75t_R _32716_ (.A1(net2854),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12542_),
    .C1(net253),
    .C2(_12543_),
    .Y(_04398_));
 INVx1_ASAP7_75t_R _32717_ (.A(_01818_),
    .Y(_12544_));
 INVx1_ASAP7_75t_R _32718_ (.A(_01785_),
    .Y(_12545_));
 AO222x2_ASAP7_75t_R _32719_ (.A1(net2781),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12544_),
    .C1(net253),
    .C2(_12545_),
    .Y(_04399_));
 INVx1_ASAP7_75t_R _32720_ (.A(_01817_),
    .Y(_12546_));
 INVx1_ASAP7_75t_R _32721_ (.A(_01784_),
    .Y(_12547_));
 AO222x2_ASAP7_75t_R _32722_ (.A1(net2910),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12546_),
    .C1(net253),
    .C2(_12547_),
    .Y(_04400_));
 INVx1_ASAP7_75t_R _32723_ (.A(_01816_),
    .Y(_12548_));
 INVx1_ASAP7_75t_R _32724_ (.A(_01783_),
    .Y(_12549_));
 AO222x2_ASAP7_75t_R _32725_ (.A1(net2814),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12548_),
    .C1(net253),
    .C2(_12549_),
    .Y(_04401_));
 INVx1_ASAP7_75t_R _32726_ (.A(_01738_),
    .Y(_12550_));
 INVx1_ASAP7_75t_R _32727_ (.A(_01782_),
    .Y(_12551_));
 AO222x2_ASAP7_75t_R _32728_ (.A1(net2862),
    .A2(_12473_),
    .B1(_12478_),
    .B2(_12550_),
    .C1(net253),
    .C2(_12551_),
    .Y(_04402_));
 NAND2x1_ASAP7_75t_R _32729_ (.A(_00239_),
    .B(net2936),
    .Y(_12552_));
 NAND2x1_ASAP7_75t_R _32730_ (.A(_06734_),
    .B(_01781_),
    .Y(_12553_));
 AOI221x1_ASAP7_75t_R _32731_ (.A1(_06724_),
    .A2(_12475_),
    .B1(_12552_),
    .B2(_12553_),
    .C(_12477_),
    .Y(_12554_));
 AOI21x1_ASAP7_75t_R _32732_ (.A1(_01814_),
    .A2(_12478_),
    .B(_12554_),
    .Y(_04403_));
 AND3x1_ASAP7_75t_R _32733_ (.A(_06618_),
    .B(_06723_),
    .C(_06744_),
    .Y(_12555_));
 AO21x2_ASAP7_75t_R _32734_ (.A1(_06724_),
    .A2(_12471_),
    .B(_12555_),
    .Y(_12556_));
 TAPCELL_ASAP7_75t_R PHY_110 ();
 TAPCELL_ASAP7_75t_R PHY_109 ();
 OR2x2_ASAP7_75t_R _32737_ (.A(net2688),
    .B(_06729_),
    .Y(_12559_));
 TAPCELL_ASAP7_75t_R PHY_108 ();
 NAND2x1_ASAP7_75t_R _32739_ (.A(_06729_),
    .B(_01780_),
    .Y(_12561_));
 AND4x1_ASAP7_75t_R _32740_ (.A(_06734_),
    .B(_06618_),
    .C(_06727_),
    .D(_06723_),
    .Y(_12562_));
 AOI21x1_ASAP7_75t_R _32741_ (.A1(_06724_),
    .A2(_12471_),
    .B(_12562_),
    .Y(_12563_));
 NOR2x1_ASAP7_75t_R _32742_ (.A(_01813_),
    .B(_06730_),
    .Y(_12564_));
 AO32x1_ASAP7_75t_R _32743_ (.A1(_12556_),
    .A2(_12559_),
    .A3(_12561_),
    .B1(_12563_),
    .B2(_12564_),
    .Y(_04404_));
 INVx1_ASAP7_75t_R _32744_ (.A(net2696),
    .Y(_12565_));
 NAND2x1_ASAP7_75t_R _32745_ (.A(_12565_),
    .B(_01815_),
    .Y(_12566_));
 NAND2x1_ASAP7_75t_R _32746_ (.A(_06729_),
    .B(_01779_),
    .Y(_12567_));
 NOR2x1_ASAP7_75t_R _32747_ (.A(_01812_),
    .B(_06730_),
    .Y(_12568_));
 TAPCELL_ASAP7_75t_R PHY_107 ();
 AO32x1_ASAP7_75t_R _32749_ (.A1(_12556_),
    .A2(_12566_),
    .A3(_12567_),
    .B1(_12568_),
    .B2(_12563_),
    .Y(_04405_));
 INVx1_ASAP7_75t_R _32750_ (.A(net2580),
    .Y(_12570_));
 NAND2x1_ASAP7_75t_R _32751_ (.A(_12570_),
    .B(_01815_),
    .Y(_12571_));
 NAND2x1_ASAP7_75t_R _32752_ (.A(_06729_),
    .B(_01778_),
    .Y(_12572_));
 NOR2x1_ASAP7_75t_R _32753_ (.A(_01811_),
    .B(_06730_),
    .Y(_12573_));
 AO32x1_ASAP7_75t_R _32754_ (.A1(_12556_),
    .A2(_12571_),
    .A3(_12572_),
    .B1(_12573_),
    .B2(_12563_),
    .Y(_04406_));
 OR2x2_ASAP7_75t_R _32755_ (.A(net2670),
    .B(_06729_),
    .Y(_12574_));
 NAND2x1_ASAP7_75t_R _32756_ (.A(_06729_),
    .B(_01777_),
    .Y(_12575_));
 NOR2x1_ASAP7_75t_R _32757_ (.A(_01810_),
    .B(_06730_),
    .Y(_12576_));
 AO32x1_ASAP7_75t_R _32758_ (.A1(_12556_),
    .A2(_12574_),
    .A3(_12575_),
    .B1(_12576_),
    .B2(_12563_),
    .Y(_04407_));
 OR2x2_ASAP7_75t_R _32759_ (.A(net2801),
    .B(_06729_),
    .Y(_12577_));
 NAND2x1_ASAP7_75t_R _32760_ (.A(_06729_),
    .B(_01776_),
    .Y(_12578_));
 NOR2x1_ASAP7_75t_R _32761_ (.A(_01809_),
    .B(_06730_),
    .Y(_12579_));
 AO32x1_ASAP7_75t_R _32762_ (.A1(_12556_),
    .A2(_12577_),
    .A3(_12578_),
    .B1(_12579_),
    .B2(_12563_),
    .Y(_04408_));
 OR2x2_ASAP7_75t_R _32763_ (.A(net2603),
    .B(_06729_),
    .Y(_12580_));
 NAND2x1_ASAP7_75t_R _32764_ (.A(_06729_),
    .B(_01775_),
    .Y(_12581_));
 NOR2x1_ASAP7_75t_R _32765_ (.A(_01808_),
    .B(_06730_),
    .Y(_12582_));
 AO32x1_ASAP7_75t_R _32766_ (.A1(_12556_),
    .A2(_12580_),
    .A3(_12581_),
    .B1(_12582_),
    .B2(_12563_),
    .Y(_04409_));
 OR2x2_ASAP7_75t_R _32767_ (.A(net2614),
    .B(_06729_),
    .Y(_12583_));
 NAND2x1_ASAP7_75t_R _32768_ (.A(_06729_),
    .B(_01774_),
    .Y(_12584_));
 NOR2x1_ASAP7_75t_R _32769_ (.A(_01807_),
    .B(_06730_),
    .Y(_12585_));
 AO32x1_ASAP7_75t_R _32770_ (.A1(_12556_),
    .A2(_12583_),
    .A3(_12584_),
    .B1(_12585_),
    .B2(_12563_),
    .Y(_04410_));
 INVx1_ASAP7_75t_R _32771_ (.A(net2607),
    .Y(_12586_));
 NAND2x1_ASAP7_75t_R _32772_ (.A(_12586_),
    .B(_01815_),
    .Y(_12587_));
 NAND2x1_ASAP7_75t_R _32773_ (.A(_06729_),
    .B(_01773_),
    .Y(_12588_));
 NOR2x1_ASAP7_75t_R _32774_ (.A(_01806_),
    .B(_06730_),
    .Y(_12589_));
 AO32x1_ASAP7_75t_R _32775_ (.A1(_12556_),
    .A2(_12587_),
    .A3(_12588_),
    .B1(_12589_),
    .B2(_12563_),
    .Y(_04411_));
 OR2x2_ASAP7_75t_R _32776_ (.A(net2682),
    .B(_06729_),
    .Y(_12590_));
 NAND2x1_ASAP7_75t_R _32777_ (.A(_06729_),
    .B(_01772_),
    .Y(_12591_));
 NOR2x1_ASAP7_75t_R _32778_ (.A(_01805_),
    .B(_06730_),
    .Y(_12592_));
 AO32x1_ASAP7_75t_R _32779_ (.A1(_12556_),
    .A2(_12590_),
    .A3(_12591_),
    .B1(_12592_),
    .B2(_12563_),
    .Y(_04412_));
 INVx1_ASAP7_75t_R _32780_ (.A(net2591),
    .Y(_12593_));
 NAND2x1_ASAP7_75t_R _32781_ (.A(_12593_),
    .B(_01815_),
    .Y(_12594_));
 NAND2x1_ASAP7_75t_R _32782_ (.A(_06729_),
    .B(_01771_),
    .Y(_12595_));
 TAPCELL_ASAP7_75t_R PHY_106 ();
 NOR2x1_ASAP7_75t_R _32784_ (.A(_01804_),
    .B(_06730_),
    .Y(_12597_));
 AO32x1_ASAP7_75t_R _32785_ (.A1(_12556_),
    .A2(_12594_),
    .A3(_12595_),
    .B1(_12597_),
    .B2(_12563_),
    .Y(_04413_));
 TAPCELL_ASAP7_75t_R PHY_105 ();
 OR2x2_ASAP7_75t_R _32787_ (.A(net2658),
    .B(_06729_),
    .Y(_12599_));
 TAPCELL_ASAP7_75t_R PHY_104 ();
 NAND2x1_ASAP7_75t_R _32789_ (.A(_06729_),
    .B(_01770_),
    .Y(_12601_));
 NOR2x1_ASAP7_75t_R _32790_ (.A(_01803_),
    .B(_06730_),
    .Y(_12602_));
 AO32x1_ASAP7_75t_R _32791_ (.A1(_12556_),
    .A2(_12599_),
    .A3(_12601_),
    .B1(_12602_),
    .B2(_12563_),
    .Y(_04414_));
 TAPCELL_ASAP7_75t_R PHY_103 ();
 OR2x2_ASAP7_75t_R _32793_ (.A(net2584),
    .B(_06729_),
    .Y(_12604_));
 NAND2x1_ASAP7_75t_R _32794_ (.A(_06729_),
    .B(_01769_),
    .Y(_12605_));
 NOR2x1_ASAP7_75t_R _32795_ (.A(_01802_),
    .B(_06730_),
    .Y(_12606_));
 TAPCELL_ASAP7_75t_R PHY_102 ();
 AO32x1_ASAP7_75t_R _32797_ (.A1(_12556_),
    .A2(_12604_),
    .A3(_12605_),
    .B1(_12606_),
    .B2(_12563_),
    .Y(_04415_));
 OR2x2_ASAP7_75t_R _32798_ (.A(net2541),
    .B(_06729_),
    .Y(_12608_));
 NAND2x1_ASAP7_75t_R _32799_ (.A(_06729_),
    .B(_01768_),
    .Y(_12609_));
 NOR2x1_ASAP7_75t_R _32800_ (.A(_01801_),
    .B(_06730_),
    .Y(_12610_));
 AO32x1_ASAP7_75t_R _32801_ (.A1(_12556_),
    .A2(_12608_),
    .A3(_12609_),
    .B1(_12610_),
    .B2(_12563_),
    .Y(_04416_));
 OR2x2_ASAP7_75t_R _32802_ (.A(net2633),
    .B(_06729_),
    .Y(_12611_));
 NAND2x1_ASAP7_75t_R _32803_ (.A(_06729_),
    .B(_01767_),
    .Y(_12612_));
 NOR2x1_ASAP7_75t_R _32804_ (.A(_01800_),
    .B(_06730_),
    .Y(_12613_));
 AO32x1_ASAP7_75t_R _32805_ (.A1(_12556_),
    .A2(_12611_),
    .A3(_12612_),
    .B1(_12613_),
    .B2(_12563_),
    .Y(_04417_));
 OR2x2_ASAP7_75t_R _32806_ (.A(net2558),
    .B(_06729_),
    .Y(_12614_));
 NAND2x1_ASAP7_75t_R _32807_ (.A(_06729_),
    .B(_01766_),
    .Y(_12615_));
 NOR2x1_ASAP7_75t_R _32808_ (.A(_01799_),
    .B(_06730_),
    .Y(_12616_));
 AO32x1_ASAP7_75t_R _32809_ (.A1(_12556_),
    .A2(_12614_),
    .A3(_12615_),
    .B1(_12616_),
    .B2(_12563_),
    .Y(_04418_));
 OR2x2_ASAP7_75t_R _32810_ (.A(net2505),
    .B(_06729_),
    .Y(_12617_));
 NAND2x1_ASAP7_75t_R _32811_ (.A(_06729_),
    .B(_01765_),
    .Y(_12618_));
 NOR2x1_ASAP7_75t_R _32812_ (.A(_01798_),
    .B(_06730_),
    .Y(_12619_));
 AO32x1_ASAP7_75t_R _32813_ (.A1(_12556_),
    .A2(_12617_),
    .A3(_12618_),
    .B1(_12619_),
    .B2(_12563_),
    .Y(_04419_));
 NAND2x1_ASAP7_75t_R _32814_ (.A(_06584_),
    .B(_01815_),
    .Y(_12620_));
 NAND2x1_ASAP7_75t_R _32815_ (.A(_06729_),
    .B(_01764_),
    .Y(_12621_));
 NOR2x1_ASAP7_75t_R _32816_ (.A(_01797_),
    .B(_06730_),
    .Y(_12622_));
 AO32x1_ASAP7_75t_R _32817_ (.A1(_12556_),
    .A2(_12620_),
    .A3(_12621_),
    .B1(_12622_),
    .B2(_12563_),
    .Y(_04420_));
 OR2x2_ASAP7_75t_R _32818_ (.A(net2625),
    .B(_06729_),
    .Y(_12623_));
 NAND2x1_ASAP7_75t_R _32819_ (.A(_06729_),
    .B(_01763_),
    .Y(_12624_));
 NOR2x1_ASAP7_75t_R _32820_ (.A(_01796_),
    .B(_06730_),
    .Y(_12625_));
 AO32x1_ASAP7_75t_R _32821_ (.A1(_12556_),
    .A2(_12623_),
    .A3(_12624_),
    .B1(_12625_),
    .B2(_12563_),
    .Y(_04421_));
 OR2x2_ASAP7_75t_R _32822_ (.A(net2618),
    .B(_06729_),
    .Y(_12626_));
 NAND2x1_ASAP7_75t_R _32823_ (.A(_06729_),
    .B(_01762_),
    .Y(_12627_));
 NOR2x1_ASAP7_75t_R _32824_ (.A(_01795_),
    .B(_06730_),
    .Y(_12628_));
 AO32x1_ASAP7_75t_R _32825_ (.A1(_12556_),
    .A2(_12626_),
    .A3(_12627_),
    .B1(_12628_),
    .B2(_12563_),
    .Y(_04422_));
 OR2x2_ASAP7_75t_R _32826_ (.A(net2652),
    .B(_06729_),
    .Y(_12629_));
 NAND2x1_ASAP7_75t_R _32827_ (.A(_06729_),
    .B(_01761_),
    .Y(_12630_));
 TAPCELL_ASAP7_75t_R PHY_101 ();
 NOR2x1_ASAP7_75t_R _32829_ (.A(_01794_),
    .B(_06730_),
    .Y(_12632_));
 AO32x1_ASAP7_75t_R _32830_ (.A1(_12556_),
    .A2(_12629_),
    .A3(_12630_),
    .B1(_12632_),
    .B2(_12563_),
    .Y(_04423_));
 TAPCELL_ASAP7_75t_R PHY_100 ();
 OR2x2_ASAP7_75t_R _32832_ (.A(net2772),
    .B(_06729_),
    .Y(_12634_));
 TAPCELL_ASAP7_75t_R PHY_99 ();
 NAND2x1_ASAP7_75t_R _32834_ (.A(_06729_),
    .B(_01760_),
    .Y(_12636_));
 NOR2x1_ASAP7_75t_R _32835_ (.A(_01793_),
    .B(_06730_),
    .Y(_12637_));
 AO32x1_ASAP7_75t_R _32836_ (.A1(_12556_),
    .A2(_12634_),
    .A3(_12636_),
    .B1(_12637_),
    .B2(_12563_),
    .Y(_04424_));
 OR2x2_ASAP7_75t_R _32837_ (.A(net2599),
    .B(_06729_),
    .Y(_12638_));
 NAND2x1_ASAP7_75t_R _32838_ (.A(_06729_),
    .B(_01759_),
    .Y(_12639_));
 NOR2x1_ASAP7_75t_R _32839_ (.A(_01792_),
    .B(_06730_),
    .Y(_12640_));
 TAPCELL_ASAP7_75t_R PHY_98 ();
 AO32x1_ASAP7_75t_R _32841_ (.A1(_12556_),
    .A2(_12638_),
    .A3(_12639_),
    .B1(_12640_),
    .B2(_12563_),
    .Y(_04425_));
 TAPCELL_ASAP7_75t_R PHY_97 ();
 OR2x2_ASAP7_75t_R _32843_ (.A(net2629),
    .B(_06729_),
    .Y(_12643_));
 NAND2x1_ASAP7_75t_R _32844_ (.A(_06729_),
    .B(_01758_),
    .Y(_12644_));
 NOR2x1_ASAP7_75t_R _32845_ (.A(_01791_),
    .B(_06730_),
    .Y(_12645_));
 AO32x1_ASAP7_75t_R _32846_ (.A1(_12556_),
    .A2(_12643_),
    .A3(_12644_),
    .B1(_12645_),
    .B2(_12563_),
    .Y(_04426_));
 OR2x2_ASAP7_75t_R _32847_ (.A(net2641),
    .B(_06729_),
    .Y(_12646_));
 NAND2x1_ASAP7_75t_R _32848_ (.A(_06729_),
    .B(_01757_),
    .Y(_12647_));
 NOR2x1_ASAP7_75t_R _32849_ (.A(_01790_),
    .B(_06730_),
    .Y(_12648_));
 AO32x1_ASAP7_75t_R _32850_ (.A1(_12556_),
    .A2(_12646_),
    .A3(_12647_),
    .B1(_12648_),
    .B2(_12563_),
    .Y(_04427_));
 OR2x2_ASAP7_75t_R _32851_ (.A(net2666),
    .B(_06729_),
    .Y(_12649_));
 NAND2x1_ASAP7_75t_R _32852_ (.A(_06729_),
    .B(_01756_),
    .Y(_12650_));
 NOR2x1_ASAP7_75t_R _32853_ (.A(_01789_),
    .B(_06730_),
    .Y(_12651_));
 AO32x1_ASAP7_75t_R _32854_ (.A1(_12556_),
    .A2(_12649_),
    .A3(_12650_),
    .B1(_12651_),
    .B2(_12563_),
    .Y(_04428_));
 OR2x2_ASAP7_75t_R _32855_ (.A(net2648),
    .B(_06729_),
    .Y(_12652_));
 NAND2x1_ASAP7_75t_R _32856_ (.A(_06729_),
    .B(_01755_),
    .Y(_12653_));
 NOR2x1_ASAP7_75t_R _32857_ (.A(_01788_),
    .B(_06730_),
    .Y(_12654_));
 AO32x1_ASAP7_75t_R _32858_ (.A1(_12556_),
    .A2(_12652_),
    .A3(_12653_),
    .B1(_12654_),
    .B2(_12563_),
    .Y(_04429_));
 OR2x2_ASAP7_75t_R _32859_ (.A(net2662),
    .B(_06729_),
    .Y(_12655_));
 NAND2x1_ASAP7_75t_R _32860_ (.A(_06729_),
    .B(_01754_),
    .Y(_12656_));
 NOR2x1_ASAP7_75t_R _32861_ (.A(_01787_),
    .B(_06730_),
    .Y(_12657_));
 AO32x1_ASAP7_75t_R _32862_ (.A1(_12556_),
    .A2(_12655_),
    .A3(_12656_),
    .B1(_12657_),
    .B2(_12563_),
    .Y(_04430_));
 OR2x2_ASAP7_75t_R _32863_ (.A(net2595),
    .B(_06729_),
    .Y(_12658_));
 NAND2x1_ASAP7_75t_R _32864_ (.A(_06729_),
    .B(_01753_),
    .Y(_12659_));
 NOR2x1_ASAP7_75t_R _32865_ (.A(_01786_),
    .B(_06730_),
    .Y(_12660_));
 AO32x1_ASAP7_75t_R _32866_ (.A1(_12556_),
    .A2(_12658_),
    .A3(_12659_),
    .B1(_12660_),
    .B2(_12563_),
    .Y(_04431_));
 OR2x2_ASAP7_75t_R _32867_ (.A(net2524),
    .B(_06729_),
    .Y(_12661_));
 NAND2x1_ASAP7_75t_R _32868_ (.A(_06729_),
    .B(_01752_),
    .Y(_12662_));
 NOR2x1_ASAP7_75t_R _32869_ (.A(_01785_),
    .B(_06730_),
    .Y(_12663_));
 AO32x1_ASAP7_75t_R _32870_ (.A1(_12556_),
    .A2(_12661_),
    .A3(_12662_),
    .B1(_12663_),
    .B2(_12563_),
    .Y(_04432_));
 OR2x2_ASAP7_75t_R _32871_ (.A(net2637),
    .B(_06729_),
    .Y(_12664_));
 NAND2x1_ASAP7_75t_R _32872_ (.A(_06729_),
    .B(_01751_),
    .Y(_12665_));
 NOR2x1_ASAP7_75t_R _32873_ (.A(_01784_),
    .B(_06730_),
    .Y(_12666_));
 AO32x1_ASAP7_75t_R _32874_ (.A1(_12556_),
    .A2(_12664_),
    .A3(_12665_),
    .B1(_12666_),
    .B2(_12563_),
    .Y(_04433_));
 OR2x2_ASAP7_75t_R _32875_ (.A(net2548),
    .B(_06729_),
    .Y(_12667_));
 NAND2x1_ASAP7_75t_R _32876_ (.A(_06729_),
    .B(_01750_),
    .Y(_12668_));
 NOR2x1_ASAP7_75t_R _32877_ (.A(_01783_),
    .B(_06730_),
    .Y(_12669_));
 AO32x1_ASAP7_75t_R _32878_ (.A1(_12556_),
    .A2(_12667_),
    .A3(_12668_),
    .B1(_12669_),
    .B2(_12563_),
    .Y(_04434_));
 OR2x2_ASAP7_75t_R _32879_ (.A(net2537),
    .B(_06729_),
    .Y(_12670_));
 NAND2x1_ASAP7_75t_R _32880_ (.A(_06729_),
    .B(_01749_),
    .Y(_12671_));
 NOR2x1_ASAP7_75t_R _32881_ (.A(_01782_),
    .B(_06730_),
    .Y(_12672_));
 AO32x1_ASAP7_75t_R _32882_ (.A1(_12556_),
    .A2(_12670_),
    .A3(_12671_),
    .B1(_12672_),
    .B2(_12563_),
    .Y(_04435_));
 NAND2x1_ASAP7_75t_R _32883_ (.A(net2936),
    .B(_01815_),
    .Y(_12673_));
 NAND2x1_ASAP7_75t_R _32884_ (.A(_06729_),
    .B(_01748_),
    .Y(_12674_));
 NOR2x1_ASAP7_75t_R _32885_ (.A(_01781_),
    .B(_06730_),
    .Y(_12675_));
 AO32x1_ASAP7_75t_R _32886_ (.A1(_12556_),
    .A2(net2937),
    .A3(_12674_),
    .B1(_12675_),
    .B2(_12563_),
    .Y(_04436_));
 OR3x4_ASAP7_75t_R _32887_ (.A(_00239_),
    .B(_06729_),
    .C(_06678_),
    .Y(_12676_));
 TAPCELL_ASAP7_75t_R PHY_96 ();
 TAPCELL_ASAP7_75t_R PHY_95 ();
 TAPCELL_ASAP7_75t_R PHY_94 ();
 NAND2x1_ASAP7_75t_R _32891_ (.A(_01780_),
    .B(_12676_),
    .Y(_12680_));
 OA21x2_ASAP7_75t_R _32892_ (.A1(net2688),
    .A2(_12676_),
    .B(_12680_),
    .Y(_04437_));
 NAND2x1_ASAP7_75t_R _32893_ (.A(_01779_),
    .B(_12676_),
    .Y(_12681_));
 OA21x2_ASAP7_75t_R _32894_ (.A1(net2696),
    .A2(_12676_),
    .B(_12681_),
    .Y(_04438_));
 NAND2x1_ASAP7_75t_R _32895_ (.A(_01778_),
    .B(_12676_),
    .Y(_12682_));
 OA21x2_ASAP7_75t_R _32896_ (.A1(net2580),
    .A2(_12676_),
    .B(_12682_),
    .Y(_04439_));
 NAND2x1_ASAP7_75t_R _32897_ (.A(_01777_),
    .B(_12676_),
    .Y(_12683_));
 OA21x2_ASAP7_75t_R _32898_ (.A1(net2670),
    .A2(_12676_),
    .B(_12683_),
    .Y(_04440_));
 NAND2x1_ASAP7_75t_R _32899_ (.A(_01776_),
    .B(_12676_),
    .Y(_12684_));
 OA21x2_ASAP7_75t_R _32900_ (.A1(net2801),
    .A2(_12676_),
    .B(_12684_),
    .Y(_04441_));
 NAND2x1_ASAP7_75t_R _32901_ (.A(_01775_),
    .B(_12676_),
    .Y(_12685_));
 OA21x2_ASAP7_75t_R _32902_ (.A1(net2603),
    .A2(_12676_),
    .B(_12685_),
    .Y(_04442_));
 NAND2x1_ASAP7_75t_R _32903_ (.A(_01774_),
    .B(_12676_),
    .Y(_12686_));
 OA21x2_ASAP7_75t_R _32904_ (.A1(net2614),
    .A2(_12676_),
    .B(_12686_),
    .Y(_04443_));
 TAPCELL_ASAP7_75t_R PHY_93 ();
 NAND2x1_ASAP7_75t_R _32906_ (.A(_01773_),
    .B(_12676_),
    .Y(_12688_));
 OA21x2_ASAP7_75t_R _32907_ (.A1(net2607),
    .A2(_12676_),
    .B(_12688_),
    .Y(_04444_));
 NAND2x1_ASAP7_75t_R _32908_ (.A(_01772_),
    .B(_12676_),
    .Y(_12689_));
 OA21x2_ASAP7_75t_R _32909_ (.A1(net2682),
    .A2(_12676_),
    .B(_12689_),
    .Y(_04445_));
 NAND2x1_ASAP7_75t_R _32910_ (.A(_01771_),
    .B(_12676_),
    .Y(_12690_));
 OA21x2_ASAP7_75t_R _32911_ (.A1(net2591),
    .A2(_12676_),
    .B(_12690_),
    .Y(_04446_));
 TAPCELL_ASAP7_75t_R PHY_92 ();
 NAND2x1_ASAP7_75t_R _32913_ (.A(_01770_),
    .B(_12676_),
    .Y(_12692_));
 OA21x2_ASAP7_75t_R _32914_ (.A1(net2658),
    .A2(_12676_),
    .B(_12692_),
    .Y(_04447_));
 NAND2x1_ASAP7_75t_R _32915_ (.A(_01769_),
    .B(_12676_),
    .Y(_12693_));
 OA21x2_ASAP7_75t_R _32916_ (.A1(net2584),
    .A2(_12676_),
    .B(_12693_),
    .Y(_04448_));
 NAND2x1_ASAP7_75t_R _32917_ (.A(_01768_),
    .B(_12676_),
    .Y(_12694_));
 OA21x2_ASAP7_75t_R _32918_ (.A1(net2789),
    .A2(_12676_),
    .B(_12694_),
    .Y(_04449_));
 NAND2x1_ASAP7_75t_R _32919_ (.A(_01767_),
    .B(_12676_),
    .Y(_12695_));
 OA21x2_ASAP7_75t_R _32920_ (.A1(net2633),
    .A2(_12676_),
    .B(_12695_),
    .Y(_04450_));
 NAND2x1_ASAP7_75t_R _32921_ (.A(_01766_),
    .B(_12676_),
    .Y(_12696_));
 OA21x2_ASAP7_75t_R _32922_ (.A1(net2558),
    .A2(_12676_),
    .B(_12696_),
    .Y(_04451_));
 NAND2x1_ASAP7_75t_R _32923_ (.A(_01765_),
    .B(_12676_),
    .Y(_12697_));
 OA21x2_ASAP7_75t_R _32924_ (.A1(net2768),
    .A2(_12676_),
    .B(_12697_),
    .Y(_04452_));
 NAND2x1_ASAP7_75t_R _32925_ (.A(_01764_),
    .B(_12676_),
    .Y(_12698_));
 OA21x2_ASAP7_75t_R _32926_ (.A1(net2692),
    .A2(_12676_),
    .B(_12698_),
    .Y(_04453_));
 TAPCELL_ASAP7_75t_R PHY_91 ();
 NAND2x1_ASAP7_75t_R _32928_ (.A(_01763_),
    .B(_12676_),
    .Y(_12700_));
 OA21x2_ASAP7_75t_R _32929_ (.A1(net2625),
    .A2(_12676_),
    .B(_12700_),
    .Y(_04454_));
 NAND2x1_ASAP7_75t_R _32930_ (.A(_01762_),
    .B(_12676_),
    .Y(_12701_));
 OA21x2_ASAP7_75t_R _32931_ (.A1(net2618),
    .A2(_12676_),
    .B(_12701_),
    .Y(_04455_));
 NAND2x1_ASAP7_75t_R _32932_ (.A(_01761_),
    .B(_12676_),
    .Y(_12702_));
 OA21x2_ASAP7_75t_R _32933_ (.A1(net2652),
    .A2(_12676_),
    .B(_12702_),
    .Y(_04456_));
 TAPCELL_ASAP7_75t_R PHY_90 ();
 NAND2x1_ASAP7_75t_R _32935_ (.A(_01760_),
    .B(_12676_),
    .Y(_12704_));
 OA21x2_ASAP7_75t_R _32936_ (.A1(net2772),
    .A2(_12676_),
    .B(_12704_),
    .Y(_04457_));
 NAND2x1_ASAP7_75t_R _32937_ (.A(_01759_),
    .B(_12676_),
    .Y(_12705_));
 OA21x2_ASAP7_75t_R _32938_ (.A1(net2599),
    .A2(_12676_),
    .B(_12705_),
    .Y(_04458_));
 NAND2x1_ASAP7_75t_R _32939_ (.A(_01758_),
    .B(_12676_),
    .Y(_12706_));
 OA21x2_ASAP7_75t_R _32940_ (.A1(net2629),
    .A2(_12676_),
    .B(_12706_),
    .Y(_04459_));
 NAND2x1_ASAP7_75t_R _32941_ (.A(_01757_),
    .B(_12676_),
    .Y(_12707_));
 OA21x2_ASAP7_75t_R _32942_ (.A1(net2641),
    .A2(_12676_),
    .B(_12707_),
    .Y(_04460_));
 NAND2x1_ASAP7_75t_R _32943_ (.A(_01756_),
    .B(_12676_),
    .Y(_12708_));
 OA21x2_ASAP7_75t_R _32944_ (.A1(net2666),
    .A2(_12676_),
    .B(_12708_),
    .Y(_04461_));
 NAND2x1_ASAP7_75t_R _32945_ (.A(_01755_),
    .B(_12676_),
    .Y(_12709_));
 OA21x2_ASAP7_75t_R _32946_ (.A1(net2648),
    .A2(_12676_),
    .B(_12709_),
    .Y(_04462_));
 NAND2x1_ASAP7_75t_R _32947_ (.A(_01754_),
    .B(_12676_),
    .Y(_12710_));
 OA21x2_ASAP7_75t_R _32948_ (.A1(net2662),
    .A2(_12676_),
    .B(_12710_),
    .Y(_04463_));
 NAND2x1_ASAP7_75t_R _32949_ (.A(_01753_),
    .B(_12676_),
    .Y(_12711_));
 OA21x2_ASAP7_75t_R _32950_ (.A1(net2595),
    .A2(_12676_),
    .B(_12711_),
    .Y(_04464_));
 NAND2x1_ASAP7_75t_R _32951_ (.A(_01752_),
    .B(_12676_),
    .Y(_12712_));
 OA21x2_ASAP7_75t_R _32952_ (.A1(net2781),
    .A2(_12676_),
    .B(_12712_),
    .Y(_04465_));
 NAND2x1_ASAP7_75t_R _32953_ (.A(_01751_),
    .B(_12676_),
    .Y(_12713_));
 OA21x2_ASAP7_75t_R _32954_ (.A1(net2637),
    .A2(_12676_),
    .B(_12713_),
    .Y(_04466_));
 NAND2x1_ASAP7_75t_R _32955_ (.A(_01750_),
    .B(_12676_),
    .Y(_12714_));
 OA21x2_ASAP7_75t_R _32956_ (.A1(net2814),
    .A2(_12676_),
    .B(_12714_),
    .Y(_04467_));
 NAND2x1_ASAP7_75t_R _32957_ (.A(_01749_),
    .B(_12676_),
    .Y(_12715_));
 OA21x2_ASAP7_75t_R _32958_ (.A1(net2537),
    .A2(_12676_),
    .B(_12715_),
    .Y(_04468_));
 NAND2x1_ASAP7_75t_R _32959_ (.A(_01748_),
    .B(_12676_),
    .Y(_12716_));
 OA21x2_ASAP7_75t_R _32960_ (.A1(net2935),
    .A2(_12676_),
    .B(_12716_),
    .Y(_04469_));
 INVx1_ASAP7_75t_R _32961_ (.A(net3948),
    .Y(_12717_));
 NAND2x1_ASAP7_75t_R _32962_ (.A(_01747_),
    .B(net3950),
    .Y(_04470_));
 OAI21x1_ASAP7_75t_R _32963_ (.A1(_01311_),
    .A2(_06366_),
    .B(_06232_),
    .Y(_04503_));
 TAPCELL_ASAP7_75t_R PHY_89 ();
 TAPCELL_ASAP7_75t_R PHY_88 ();
 AND2x2_ASAP7_75t_R _32966_ (.A(net431),
    .B(net2688),
    .Y(_12720_));
 AO21x1_ASAP7_75t_R _32967_ (.A1(_06580_),
    .A2(net2692),
    .B(_12720_),
    .Y(_12721_));
 NAND2x1_ASAP7_75t_R _32968_ (.A(net431),
    .B(_01846_),
    .Y(_12722_));
 OA211x2_ASAP7_75t_R _32969_ (.A1(net431),
    .A2(_12517_),
    .B(_12722_),
    .C(_06589_),
    .Y(_12723_));
 AO21x2_ASAP7_75t_R _32970_ (.A1(_00240_),
    .A2(_12721_),
    .B(_12723_),
    .Y(_12724_));
 TAPCELL_ASAP7_75t_R PHY_87 ();
 TAPCELL_ASAP7_75t_R PHY_86 ();
 TAPCELL_ASAP7_75t_R PHY_85 ();
 NAND2x1_ASAP7_75t_R _32974_ (.A(_01723_),
    .B(net254),
    .Y(_12728_));
 OA21x2_ASAP7_75t_R _32975_ (.A1(net254),
    .A2(_12724_),
    .B(_12728_),
    .Y(_02597_));
 AND2x2_ASAP7_75t_R _32976_ (.A(net431),
    .B(net2696),
    .Y(_12729_));
 AO21x1_ASAP7_75t_R _32977_ (.A1(_06580_),
    .A2(net2625),
    .B(_12729_),
    .Y(_12730_));
 NAND2x1_ASAP7_75t_R _32978_ (.A(net431),
    .B(_01845_),
    .Y(_12731_));
 OA211x2_ASAP7_75t_R _32979_ (.A1(net431),
    .A2(_12519_),
    .B(_12731_),
    .C(_06589_),
    .Y(_12732_));
 AO21x2_ASAP7_75t_R _32980_ (.A1(_00240_),
    .A2(_12730_),
    .B(_12732_),
    .Y(_12733_));
 TAPCELL_ASAP7_75t_R PHY_84 ();
 TAPCELL_ASAP7_75t_R PHY_83 ();
 NAND2x1_ASAP7_75t_R _32983_ (.A(_00164_),
    .B(net254),
    .Y(_12736_));
 OA21x2_ASAP7_75t_R _32984_ (.A1(net254),
    .A2(_12733_),
    .B(_12736_),
    .Y(_02598_));
 TAPCELL_ASAP7_75t_R PHY_82 ();
 AND2x2_ASAP7_75t_R _32986_ (.A(net431),
    .B(net2580),
    .Y(_12738_));
 AO21x1_ASAP7_75t_R _32987_ (.A1(_06580_),
    .A2(net2618),
    .B(_12738_),
    .Y(_12739_));
 NAND2x1_ASAP7_75t_R _32988_ (.A(net431),
    .B(_01844_),
    .Y(_12740_));
 OA211x2_ASAP7_75t_R _32989_ (.A1(net431),
    .A2(_12521_),
    .B(_12740_),
    .C(_06589_),
    .Y(_12741_));
 AO21x2_ASAP7_75t_R _32990_ (.A1(_00240_),
    .A2(_12739_),
    .B(_12741_),
    .Y(_12742_));
 TAPCELL_ASAP7_75t_R PHY_81 ();
 NAND2x1_ASAP7_75t_R _32992_ (.A(_00166_),
    .B(net254),
    .Y(_12744_));
 OA21x2_ASAP7_75t_R _32993_ (.A1(net254),
    .A2(_12742_),
    .B(_12744_),
    .Y(_02599_));
 TAPCELL_ASAP7_75t_R PHY_80 ();
 AND2x2_ASAP7_75t_R _32995_ (.A(net431),
    .B(net2670),
    .Y(_12746_));
 AO21x1_ASAP7_75t_R _32996_ (.A1(_06580_),
    .A2(net2652),
    .B(_12746_),
    .Y(_12747_));
 NAND2x1_ASAP7_75t_R _32997_ (.A(net431),
    .B(_01843_),
    .Y(_12748_));
 OA211x2_ASAP7_75t_R _32998_ (.A1(net431),
    .A2(_12524_),
    .B(_12748_),
    .C(_06589_),
    .Y(_12749_));
 AO21x2_ASAP7_75t_R _32999_ (.A1(net428),
    .A2(_12747_),
    .B(_12749_),
    .Y(_12750_));
 TAPCELL_ASAP7_75t_R PHY_79 ();
 NAND2x1_ASAP7_75t_R _33001_ (.A(_00169_),
    .B(net254),
    .Y(_12752_));
 OA21x2_ASAP7_75t_R _33002_ (.A1(net254),
    .A2(_12750_),
    .B(_12752_),
    .Y(_02600_));
 AND2x2_ASAP7_75t_R _33003_ (.A(net431),
    .B(net2801),
    .Y(_12753_));
 AO21x1_ASAP7_75t_R _33004_ (.A1(_06580_),
    .A2(net2772),
    .B(_12753_),
    .Y(_12754_));
 NAND2x1_ASAP7_75t_R _33005_ (.A(net431),
    .B(_01842_),
    .Y(_12755_));
 OA211x2_ASAP7_75t_R _33006_ (.A1(net431),
    .A2(_12527_),
    .B(_12755_),
    .C(_06589_),
    .Y(_12756_));
 AO21x2_ASAP7_75t_R _33007_ (.A1(net428),
    .A2(_12754_),
    .B(_12756_),
    .Y(_12757_));
 TAPCELL_ASAP7_75t_R PHY_78 ();
 NAND2x1_ASAP7_75t_R _33009_ (.A(_00173_),
    .B(net254),
    .Y(_12759_));
 OA21x2_ASAP7_75t_R _33010_ (.A1(net254),
    .A2(_12757_),
    .B(_12759_),
    .Y(_02601_));
 AND2x2_ASAP7_75t_R _33011_ (.A(net430),
    .B(net2603),
    .Y(_12760_));
 AO21x1_ASAP7_75t_R _33012_ (.A1(_06580_),
    .A2(net2599),
    .B(_12760_),
    .Y(_12761_));
 NAND2x1_ASAP7_75t_R _33013_ (.A(net430),
    .B(_01841_),
    .Y(_12762_));
 OA211x2_ASAP7_75t_R _33014_ (.A1(net430),
    .A2(_12530_),
    .B(_12762_),
    .C(_06589_),
    .Y(_12763_));
 AO21x2_ASAP7_75t_R _33015_ (.A1(net428),
    .A2(_12761_),
    .B(_12763_),
    .Y(_12764_));
 TAPCELL_ASAP7_75t_R PHY_77 ();
 NAND2x1_ASAP7_75t_R _33017_ (.A(_00176_),
    .B(net254),
    .Y(_12766_));
 OA21x2_ASAP7_75t_R _33018_ (.A1(net254),
    .A2(_12764_),
    .B(_12766_),
    .Y(_02602_));
 AND2x2_ASAP7_75t_R _33019_ (.A(net430),
    .B(net2614),
    .Y(_12767_));
 AO21x1_ASAP7_75t_R _33020_ (.A1(_06580_),
    .A2(net2629),
    .B(_12767_),
    .Y(_12768_));
 NAND2x1_ASAP7_75t_R _33021_ (.A(net430),
    .B(_01840_),
    .Y(_12769_));
 OA211x2_ASAP7_75t_R _33022_ (.A1(net430),
    .A2(_12532_),
    .B(_12769_),
    .C(_06589_),
    .Y(_12770_));
 AO21x2_ASAP7_75t_R _33023_ (.A1(net428),
    .A2(_12768_),
    .B(_12770_),
    .Y(_12771_));
 TAPCELL_ASAP7_75t_R PHY_76 ();
 NAND2x1_ASAP7_75t_R _33025_ (.A(_00179_),
    .B(net254),
    .Y(_12773_));
 OA21x2_ASAP7_75t_R _33026_ (.A1(net254),
    .A2(_12771_),
    .B(_12773_),
    .Y(_02603_));
 TAPCELL_ASAP7_75t_R PHY_75 ();
 TAPCELL_ASAP7_75t_R PHY_74 ();
 AND2x2_ASAP7_75t_R _33029_ (.A(net431),
    .B(net2607),
    .Y(_12776_));
 AO21x1_ASAP7_75t_R _33030_ (.A1(_06580_),
    .A2(net2641),
    .B(_12776_),
    .Y(_12777_));
 NAND2x1_ASAP7_75t_R _33031_ (.A(net431),
    .B(_01839_),
    .Y(_12778_));
 OA211x2_ASAP7_75t_R _33032_ (.A1(net431),
    .A2(_12534_),
    .B(_12778_),
    .C(_06589_),
    .Y(_12779_));
 AO21x2_ASAP7_75t_R _33033_ (.A1(_00240_),
    .A2(_12777_),
    .B(_12779_),
    .Y(_12780_));
 TAPCELL_ASAP7_75t_R PHY_73 ();
 NAND2x1_ASAP7_75t_R _33035_ (.A(_00181_),
    .B(net254),
    .Y(_12782_));
 OA21x2_ASAP7_75t_R _33036_ (.A1(net254),
    .A2(_12780_),
    .B(_12782_),
    .Y(_02604_));
 AND2x2_ASAP7_75t_R _33037_ (.A(net431),
    .B(net2682),
    .Y(_12783_));
 AO21x1_ASAP7_75t_R _33038_ (.A1(_06580_),
    .A2(net2666),
    .B(_12783_),
    .Y(_12784_));
 NAND2x1_ASAP7_75t_R _33039_ (.A(net431),
    .B(_01838_),
    .Y(_12785_));
 OA211x2_ASAP7_75t_R _33040_ (.A1(net431),
    .A2(_12536_),
    .B(_12785_),
    .C(_06589_),
    .Y(_12786_));
 AO21x2_ASAP7_75t_R _33041_ (.A1(net428),
    .A2(_12784_),
    .B(_12786_),
    .Y(_12787_));
 TAPCELL_ASAP7_75t_R PHY_72 ();
 NAND2x1_ASAP7_75t_R _33043_ (.A(_00185_),
    .B(net254),
    .Y(_12789_));
 OA21x2_ASAP7_75t_R _33044_ (.A1(net254),
    .A2(_12787_),
    .B(_12789_),
    .Y(_02605_));
 AND2x2_ASAP7_75t_R _33045_ (.A(net431),
    .B(net2591),
    .Y(_12790_));
 AO21x1_ASAP7_75t_R _33046_ (.A1(_06580_),
    .A2(net2648),
    .B(_12790_),
    .Y(_12791_));
 NAND2x1_ASAP7_75t_R _33047_ (.A(net431),
    .B(_01837_),
    .Y(_12792_));
 OA211x2_ASAP7_75t_R _33048_ (.A1(net431),
    .A2(_12538_),
    .B(_12792_),
    .C(_06589_),
    .Y(_12793_));
 AO21x2_ASAP7_75t_R _33049_ (.A1(_00240_),
    .A2(_12791_),
    .B(_12793_),
    .Y(_12794_));
 NAND2x1_ASAP7_75t_R _33050_ (.A(_00188_),
    .B(net254),
    .Y(_12795_));
 OA21x2_ASAP7_75t_R _33051_ (.A1(net254),
    .A2(_12794_),
    .B(_12795_),
    .Y(_02606_));
 AND2x2_ASAP7_75t_R _33052_ (.A(net430),
    .B(net2658),
    .Y(_12796_));
 AO21x1_ASAP7_75t_R _33053_ (.A1(_06580_),
    .A2(net2662),
    .B(_12796_),
    .Y(_12797_));
 NAND2x1_ASAP7_75t_R _33054_ (.A(net430),
    .B(_01836_),
    .Y(_12798_));
 OA211x2_ASAP7_75t_R _33055_ (.A1(net430),
    .A2(_12540_),
    .B(_12798_),
    .C(_06589_),
    .Y(_12799_));
 AO21x2_ASAP7_75t_R _33056_ (.A1(net428),
    .A2(_12797_),
    .B(_12799_),
    .Y(_12800_));
 TAPCELL_ASAP7_75t_R PHY_71 ();
 NAND2x1_ASAP7_75t_R _33058_ (.A(_00192_),
    .B(net254),
    .Y(_12802_));
 OA21x2_ASAP7_75t_R _33059_ (.A1(net254),
    .A2(_12800_),
    .B(_12802_),
    .Y(_02607_));
 AND2x2_ASAP7_75t_R _33060_ (.A(net430),
    .B(net2584),
    .Y(_12803_));
 AO21x1_ASAP7_75t_R _33061_ (.A1(_06580_),
    .A2(net2595),
    .B(_12803_),
    .Y(_12804_));
 NAND2x1_ASAP7_75t_R _33062_ (.A(net430),
    .B(_01835_),
    .Y(_12805_));
 OA211x2_ASAP7_75t_R _33063_ (.A1(net430),
    .A2(_12542_),
    .B(_12805_),
    .C(_06589_),
    .Y(_12806_));
 AO21x2_ASAP7_75t_R _33064_ (.A1(net428),
    .A2(_12804_),
    .B(_12806_),
    .Y(_12807_));
 TAPCELL_ASAP7_75t_R PHY_70 ();
 NAND2x1_ASAP7_75t_R _33066_ (.A(_00195_),
    .B(net254),
    .Y(_12809_));
 OA21x2_ASAP7_75t_R _33067_ (.A1(net254),
    .A2(_12807_),
    .B(_12809_),
    .Y(_02608_));
 AND2x2_ASAP7_75t_R _33068_ (.A(net430),
    .B(net2541),
    .Y(_12810_));
 AO21x1_ASAP7_75t_R _33069_ (.A1(_06580_),
    .A2(net2524),
    .B(_12810_),
    .Y(_12811_));
 NAND2x1_ASAP7_75t_R _33070_ (.A(net430),
    .B(_01834_),
    .Y(_12812_));
 OA211x2_ASAP7_75t_R _33071_ (.A1(net430),
    .A2(_12544_),
    .B(_12812_),
    .C(_06589_),
    .Y(_12813_));
 AO21x2_ASAP7_75t_R _33072_ (.A1(net428),
    .A2(_12811_),
    .B(_12813_),
    .Y(_12814_));
 TAPCELL_ASAP7_75t_R PHY_69 ();
 TAPCELL_ASAP7_75t_R PHY_68 ();
 TAPCELL_ASAP7_75t_R PHY_67 ();
 NAND2x1_ASAP7_75t_R _33076_ (.A(_00198_),
    .B(net254),
    .Y(_12818_));
 OA21x2_ASAP7_75t_R _33077_ (.A1(net254),
    .A2(_12814_),
    .B(_12818_),
    .Y(_02609_));
 AND2x2_ASAP7_75t_R _33078_ (.A(net430),
    .B(net2633),
    .Y(_12819_));
 AO21x1_ASAP7_75t_R _33079_ (.A1(_06580_),
    .A2(net2637),
    .B(_12819_),
    .Y(_12820_));
 NAND2x1_ASAP7_75t_R _33080_ (.A(net431),
    .B(_01833_),
    .Y(_12821_));
 OA211x2_ASAP7_75t_R _33081_ (.A1(net431),
    .A2(_12546_),
    .B(_12821_),
    .C(_06589_),
    .Y(_12822_));
 AO21x2_ASAP7_75t_R _33082_ (.A1(_00240_),
    .A2(_12820_),
    .B(_12822_),
    .Y(_12823_));
 TAPCELL_ASAP7_75t_R PHY_66 ();
 TAPCELL_ASAP7_75t_R PHY_65 ();
 TAPCELL_ASAP7_75t_R PHY_64 ();
 NAND2x1_ASAP7_75t_R _33086_ (.A(_00200_),
    .B(net254),
    .Y(_12827_));
 OA21x2_ASAP7_75t_R _33087_ (.A1(net254),
    .A2(_12823_),
    .B(_12827_),
    .Y(_02610_));
 AND2x2_ASAP7_75t_R _33088_ (.A(net430),
    .B(net2558),
    .Y(_12828_));
 AO21x1_ASAP7_75t_R _33089_ (.A1(_06580_),
    .A2(net2548),
    .B(_12828_),
    .Y(_12829_));
 NAND2x1_ASAP7_75t_R _33090_ (.A(net430),
    .B(_01832_),
    .Y(_12830_));
 OA211x2_ASAP7_75t_R _33091_ (.A1(net430),
    .A2(_12548_),
    .B(_12830_),
    .C(_06589_),
    .Y(_12831_));
 AO21x2_ASAP7_75t_R _33092_ (.A1(net428),
    .A2(_12829_),
    .B(_12831_),
    .Y(_12832_));
 TAPCELL_ASAP7_75t_R PHY_63 ();
 TAPCELL_ASAP7_75t_R PHY_62 ();
 NAND2x1_ASAP7_75t_R _33095_ (.A(_00203_),
    .B(net254),
    .Y(_12835_));
 OA21x2_ASAP7_75t_R _33096_ (.A1(net254),
    .A2(_12832_),
    .B(_12835_),
    .Y(_02611_));
 AND2x2_ASAP7_75t_R _33097_ (.A(net2505),
    .B(net430),
    .Y(_12836_));
 AO21x1_ASAP7_75t_R _33098_ (.A1(net2537),
    .A2(_06580_),
    .B(_12836_),
    .Y(_12837_));
 NAND2x1_ASAP7_75t_R _33099_ (.A(net430),
    .B(_01831_),
    .Y(_12838_));
 OA211x2_ASAP7_75t_R _33100_ (.A1(net430),
    .A2(_12550_),
    .B(_12838_),
    .C(_06589_),
    .Y(_12839_));
 AO21x2_ASAP7_75t_R _33101_ (.A1(net428),
    .A2(_12837_),
    .B(_12839_),
    .Y(_12840_));
 TAPCELL_ASAP7_75t_R PHY_61 ();
 TAPCELL_ASAP7_75t_R PHY_60 ();
 NAND2x1_ASAP7_75t_R _33104_ (.A(_00205_),
    .B(net254),
    .Y(_12843_));
 OA21x2_ASAP7_75t_R _33105_ (.A1(net254),
    .A2(_12840_),
    .B(_12843_),
    .Y(_02612_));
 TAPCELL_ASAP7_75t_R PHY_59 ();
 AND2x4_ASAP7_75t_R _33107_ (.A(_12724_),
    .B(_12733_),
    .Y(_12845_));
 NAND2x1_ASAP7_75t_R _33108_ (.A(_06686_),
    .B(_12845_),
    .Y(_12846_));
 OA21x2_ASAP7_75t_R _33109_ (.A1(_05659_),
    .A2(_06686_),
    .B(_12846_),
    .Y(_02613_));
 INVx1_ASAP7_75t_R _33110_ (.A(_01814_),
    .Y(_12847_));
 OR3x1_ASAP7_75t_R _33111_ (.A(_00240_),
    .B(_06734_),
    .C(net2936),
    .Y(_12848_));
 OA21x2_ASAP7_75t_R _33112_ (.A1(_00239_),
    .A2(_01781_),
    .B(_12848_),
    .Y(_12849_));
 OR4x1_ASAP7_75t_R _33113_ (.A(_00662_),
    .B(_12847_),
    .C(net255),
    .D(_12849_),
    .Y(_12850_));
 OAI21x1_ASAP7_75t_R _33114_ (.A1(_01722_),
    .A2(_06686_),
    .B(_12850_),
    .Y(_02614_));
 OA21x2_ASAP7_75t_R _33115_ (.A1(net2936),
    .A2(_06588_),
    .B(_00239_),
    .Y(_12851_));
 OAI21x1_ASAP7_75t_R _33116_ (.A1(net431),
    .A2(_12851_),
    .B(_06593_),
    .Y(_12852_));
 NOR2x1_ASAP7_75t_R _33117_ (.A(_01781_),
    .B(_06676_),
    .Y(_12853_));
 OR4x1_ASAP7_75t_R _33118_ (.A(_00662_),
    .B(_00239_),
    .C(_12847_),
    .D(_12853_),
    .Y(_12854_));
 AND3x1_ASAP7_75t_R _33119_ (.A(_06686_),
    .B(_12852_),
    .C(_12854_),
    .Y(_12855_));
 AO21x1_ASAP7_75t_R _33120_ (.A1(_05744_),
    .A2(net255),
    .B(_12855_),
    .Y(_02615_));
 TAPCELL_ASAP7_75t_R PHY_58 ();
 TAPCELL_ASAP7_75t_R PHY_57 ();
 TAPCELL_ASAP7_75t_R PHY_56 ();
 AO21x1_ASAP7_75t_R _33124_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[1] ),
    .Y(_12859_));
 OA21x2_ASAP7_75t_R _33125_ (.A1(_06580_),
    .A2(net255),
    .B(_12859_),
    .Y(_02616_));
 AO21x1_ASAP7_75t_R _33126_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[2] ),
    .Y(_12860_));
 OA21x2_ASAP7_75t_R _33127_ (.A1(\cs_registers_i.pc_if_i[2] ),
    .A2(net255),
    .B(_12860_),
    .Y(_02617_));
 AO21x1_ASAP7_75t_R _33128_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[3] ),
    .Y(_12861_));
 OA21x2_ASAP7_75t_R _33129_ (.A1(\cs_registers_i.pc_if_i[3] ),
    .A2(net255),
    .B(_12861_),
    .Y(_02618_));
 NAND2x1_ASAP7_75t_R _33130_ (.A(_01605_),
    .B(_06686_),
    .Y(_12862_));
 OA21x2_ASAP7_75t_R _33131_ (.A1(_15051_),
    .A2(_06686_),
    .B(_12862_),
    .Y(_02619_));
 AO21x1_ASAP7_75t_R _33132_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[5] ),
    .Y(_12863_));
 OA21x2_ASAP7_75t_R _33133_ (.A1(\cs_registers_i.pc_if_i[5] ),
    .A2(net255),
    .B(_12863_),
    .Y(_02620_));
 NAND2x1_ASAP7_75t_R _33134_ (.A(_01603_),
    .B(_06686_),
    .Y(_12864_));
 OA21x2_ASAP7_75t_R _33135_ (.A1(_15169_),
    .A2(_06686_),
    .B(_12864_),
    .Y(_02621_));
 AO21x1_ASAP7_75t_R _33136_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[7] ),
    .Y(_12865_));
 OA21x2_ASAP7_75t_R _33137_ (.A1(\cs_registers_i.pc_if_i[7] ),
    .A2(net255),
    .B(_12865_),
    .Y(_02622_));
 TAPCELL_ASAP7_75t_R PHY_55 ();
 TAPCELL_ASAP7_75t_R PHY_54 ();
 TAPCELL_ASAP7_75t_R PHY_53 ();
 AND3x1_ASAP7_75t_R _33141_ (.A(_01601_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12869_));
 AOI21x1_ASAP7_75t_R _33142_ (.A1(_00186_),
    .A2(net255),
    .B(_12869_),
    .Y(_02623_));
 TAPCELL_ASAP7_75t_R PHY_52 ();
 AO21x1_ASAP7_75t_R _33144_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[9] ),
    .Y(_12871_));
 OA21x2_ASAP7_75t_R _33145_ (.A1(\cs_registers_i.pc_if_i[9] ),
    .A2(net255),
    .B(_12871_),
    .Y(_02624_));
 NAND2x1_ASAP7_75t_R _33146_ (.A(_01599_),
    .B(_06686_),
    .Y(_12872_));
 OA21x2_ASAP7_75t_R _33147_ (.A1(_15398_),
    .A2(_06686_),
    .B(_12872_),
    .Y(_02625_));
 AO21x1_ASAP7_75t_R _33148_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[11] ),
    .Y(_12873_));
 OA21x2_ASAP7_75t_R _33149_ (.A1(\cs_registers_i.pc_if_i[11] ),
    .A2(net255),
    .B(_12873_),
    .Y(_02626_));
 AND3x1_ASAP7_75t_R _33150_ (.A(_01597_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12874_));
 AOI21x1_ASAP7_75t_R _33151_ (.A1(_00199_),
    .A2(net255),
    .B(_12874_),
    .Y(_02627_));
 AO21x1_ASAP7_75t_R _33152_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[13] ),
    .Y(_12875_));
 OA21x2_ASAP7_75t_R _33153_ (.A1(\cs_registers_i.pc_if_i[13] ),
    .A2(net255),
    .B(_12875_),
    .Y(_02628_));
 NAND2x1_ASAP7_75t_R _33154_ (.A(_01595_),
    .B(_06686_),
    .Y(_12876_));
 OA21x2_ASAP7_75t_R _33155_ (.A1(_15775_),
    .A2(_06686_),
    .B(_12876_),
    .Y(_02629_));
 AO21x1_ASAP7_75t_R _33156_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[15] ),
    .Y(_12877_));
 OA21x2_ASAP7_75t_R _33157_ (.A1(\cs_registers_i.pc_if_i[15] ),
    .A2(net255),
    .B(_12877_),
    .Y(_02630_));
 AND3x1_ASAP7_75t_R _33158_ (.A(_01593_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12878_));
 AOI21x1_ASAP7_75t_R _33159_ (.A1(_00208_),
    .A2(net255),
    .B(_12878_),
    .Y(_02631_));
 AO21x1_ASAP7_75t_R _33160_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[17] ),
    .Y(_12879_));
 OA21x2_ASAP7_75t_R _33161_ (.A1(\cs_registers_i.pc_if_i[17] ),
    .A2(net255),
    .B(_12879_),
    .Y(_02632_));
 AND3x1_ASAP7_75t_R _33162_ (.A(_01591_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12880_));
 AOI21x1_ASAP7_75t_R _33163_ (.A1(_00211_),
    .A2(net255),
    .B(_12880_),
    .Y(_02633_));
 TAPCELL_ASAP7_75t_R PHY_51 ();
 TAPCELL_ASAP7_75t_R PHY_50 ();
 AO21x1_ASAP7_75t_R _33166_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[19] ),
    .Y(_12883_));
 OA21x2_ASAP7_75t_R _33167_ (.A1(\cs_registers_i.pc_if_i[19] ),
    .A2(net255),
    .B(_12883_),
    .Y(_02634_));
 AND3x1_ASAP7_75t_R _33168_ (.A(_01589_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12884_));
 AOI21x1_ASAP7_75t_R _33169_ (.A1(_00214_),
    .A2(net255),
    .B(_12884_),
    .Y(_02635_));
 AO21x1_ASAP7_75t_R _33170_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[21] ),
    .Y(_12885_));
 OA21x2_ASAP7_75t_R _33171_ (.A1(\cs_registers_i.pc_if_i[21] ),
    .A2(net255),
    .B(_12885_),
    .Y(_02636_));
 AND3x1_ASAP7_75t_R _33172_ (.A(_01587_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12886_));
 AOI21x1_ASAP7_75t_R _33173_ (.A1(_00217_),
    .A2(net255),
    .B(_12886_),
    .Y(_02637_));
 AO21x1_ASAP7_75t_R _33174_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[23] ),
    .Y(_12887_));
 OA21x2_ASAP7_75t_R _33175_ (.A1(\cs_registers_i.pc_if_i[23] ),
    .A2(net255),
    .B(_12887_),
    .Y(_02638_));
 AND3x1_ASAP7_75t_R _33176_ (.A(_01585_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12888_));
 AOI21x1_ASAP7_75t_R _33177_ (.A1(_00220_),
    .A2(net255),
    .B(_12888_),
    .Y(_02639_));
 AO21x1_ASAP7_75t_R _33178_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[25] ),
    .Y(_12889_));
 OA21x2_ASAP7_75t_R _33179_ (.A1(\cs_registers_i.pc_if_i[25] ),
    .A2(net255),
    .B(_12889_),
    .Y(_02640_));
 AND3x1_ASAP7_75t_R _33180_ (.A(_01583_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12890_));
 AOI21x1_ASAP7_75t_R _33181_ (.A1(_00223_),
    .A2(net255),
    .B(_12890_),
    .Y(_02641_));
 AO21x1_ASAP7_75t_R _33182_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[27] ),
    .Y(_12891_));
 OA21x2_ASAP7_75t_R _33183_ (.A1(\cs_registers_i.pc_if_i[27] ),
    .A2(net255),
    .B(_12891_),
    .Y(_02642_));
 AND3x1_ASAP7_75t_R _33184_ (.A(_01581_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12892_));
 AOI21x1_ASAP7_75t_R _33185_ (.A1(_00226_),
    .A2(net255),
    .B(_12892_),
    .Y(_02643_));
 AO21x1_ASAP7_75t_R _33186_ (.A1(_06618_),
    .A2(_06685_),
    .B(\cs_registers_i.pc_id_i[29] ),
    .Y(_12893_));
 OA21x2_ASAP7_75t_R _33187_ (.A1(\cs_registers_i.pc_if_i[29] ),
    .A2(net255),
    .B(_12893_),
    .Y(_02644_));
 NAND2x1_ASAP7_75t_R _33188_ (.A(_01579_),
    .B(_06686_),
    .Y(_12894_));
 OA21x2_ASAP7_75t_R _33189_ (.A1(_05401_),
    .A2(_06686_),
    .B(_12894_),
    .Y(_02645_));
 AND3x1_ASAP7_75t_R _33190_ (.A(_01578_),
    .B(_06618_),
    .C(_06685_),
    .Y(_12895_));
 AOI21x1_ASAP7_75t_R _33191_ (.A1(_00230_),
    .A2(net255),
    .B(_12895_),
    .Y(_02646_));
 INVx1_ASAP7_75t_R _33192_ (.A(_09452_),
    .Y(_12896_));
 AND2x2_ASAP7_75t_R _33193_ (.A(_05693_),
    .B(_11141_),
    .Y(_12897_));
 AND4x2_ASAP7_75t_R _33194_ (.A(_11087_),
    .B(_12896_),
    .C(net3517),
    .D(_12897_),
    .Y(_12898_));
 AO21x1_ASAP7_75t_R _33195_ (.A1(_01577_),
    .A2(_11894_),
    .B(_06935_),
    .Y(_12899_));
 OAI22x1_ASAP7_75t_R _33196_ (.A1(_02140_),
    .A2(_06932_),
    .B1(_12898_),
    .B2(_12899_),
    .Y(_02863_));
 AO21x1_ASAP7_75t_R _33197_ (.A1(_01576_),
    .A2(_11894_),
    .B(_06935_),
    .Y(_12900_));
 OAI22x1_ASAP7_75t_R _33198_ (.A1(_17810_),
    .A2(_06932_),
    .B1(_12898_),
    .B2(_12900_),
    .Y(_02864_));
 NAND2x1_ASAP7_75t_R _33199_ (.A(_01875_),
    .B(_14845_),
    .Y(_12901_));
 OA21x2_ASAP7_75t_R _33200_ (.A1(_14788_),
    .A2(_14845_),
    .B(_12901_),
    .Y(_04341_));
 AND3x1_ASAP7_75t_R _33201_ (.A(_00279_),
    .B(_01875_),
    .C(_14843_),
    .Y(_12902_));
 AOI21x1_ASAP7_75t_R _33202_ (.A1(_01874_),
    .A2(_14845_),
    .B(_12902_),
    .Y(_04342_));
 AOI21x1_ASAP7_75t_R _33203_ (.A1(net428),
    .A2(_12811_),
    .B(_12813_),
    .Y(_12903_));
 AOI21x1_ASAP7_75t_R _33204_ (.A1(net428),
    .A2(_12837_),
    .B(_12839_),
    .Y(_12904_));
 OR3x4_ASAP7_75t_R _33205_ (.A(_12823_),
    .B(_12832_),
    .C(_12904_),
    .Y(_12905_));
 AOI21x1_ASAP7_75t_R _33206_ (.A1(net428),
    .A2(_12797_),
    .B(_12799_),
    .Y(_12906_));
 AND2x2_ASAP7_75t_R _33207_ (.A(_12906_),
    .B(_12807_),
    .Y(_12907_));
 NOR3x1_ASAP7_75t_R _33208_ (.A(_12903_),
    .B(_12905_),
    .C(_12907_),
    .Y(_12908_));
 OR2x2_ASAP7_75t_R _33209_ (.A(_12764_),
    .B(_12771_),
    .Y(_12909_));
 OR3x4_ASAP7_75t_R _33210_ (.A(_12742_),
    .B(_12750_),
    .C(_12909_),
    .Y(_12910_));
 NOR2x2_ASAP7_75t_R _33211_ (.A(_12757_),
    .B(_12910_),
    .Y(_12911_));
 AND3x2_ASAP7_75t_R _33212_ (.A(_12823_),
    .B(_12832_),
    .C(_12904_),
    .Y(_12912_));
 AND3x1_ASAP7_75t_R _33213_ (.A(_12903_),
    .B(_12911_),
    .C(_12912_),
    .Y(_12913_));
 AOI21x1_ASAP7_75t_R _33214_ (.A1(_00240_),
    .A2(_12730_),
    .B(_12732_),
    .Y(_12914_));
 AND2x6_ASAP7_75t_R _33215_ (.A(_12724_),
    .B(_12914_),
    .Y(_12915_));
 TAPCELL_ASAP7_75t_R PHY_49 ();
 TAPCELL_ASAP7_75t_R PHY_48 ();
 OA21x2_ASAP7_75t_R _33218_ (.A1(_12908_),
    .A2(_12913_),
    .B(_12915_),
    .Y(_12918_));
 AOI21x1_ASAP7_75t_R _33219_ (.A1(net428),
    .A2(_12829_),
    .B(_12831_),
    .Y(_12919_));
 TAPCELL_ASAP7_75t_R PHY_47 ();
 AND2x2_ASAP7_75t_R _33221_ (.A(_12919_),
    .B(_12840_),
    .Y(_12921_));
 NOR2x2_ASAP7_75t_R _33222_ (.A(_12823_),
    .B(_12921_),
    .Y(_12922_));
 OR4x1_ASAP7_75t_R _33223_ (.A(_12780_),
    .B(_12794_),
    .C(_12800_),
    .D(_12807_),
    .Y(_12923_));
 OR2x2_ASAP7_75t_R _33224_ (.A(_12787_),
    .B(_12923_),
    .Y(_12924_));
 OR4x1_ASAP7_75t_R _33225_ (.A(_12814_),
    .B(_12832_),
    .C(_12909_),
    .D(_12924_),
    .Y(_12925_));
 AOI21x1_ASAP7_75t_R _33226_ (.A1(_00240_),
    .A2(_12721_),
    .B(_12723_),
    .Y(_12926_));
 AND2x6_ASAP7_75t_R _33227_ (.A(_12926_),
    .B(_12914_),
    .Y(_12927_));
 INVx1_ASAP7_75t_R _33228_ (.A(_12927_),
    .Y(_12928_));
 AOI21x1_ASAP7_75t_R _33229_ (.A1(_12922_),
    .A2(_12925_),
    .B(_12928_),
    .Y(_12929_));
 OR3x4_ASAP7_75t_R _33230_ (.A(_12823_),
    .B(_12832_),
    .C(_12840_),
    .Y(_12930_));
 TAPCELL_ASAP7_75t_R PHY_46 ();
 AND2x6_ASAP7_75t_R _33232_ (.A(_12926_),
    .B(_12733_),
    .Y(_12932_));
 TAPCELL_ASAP7_75t_R PHY_45 ();
 OR2x2_ASAP7_75t_R _33234_ (.A(_12757_),
    .B(_12910_),
    .Y(_12934_));
 OR3x1_ASAP7_75t_R _33235_ (.A(_12814_),
    .B(_12832_),
    .C(_12934_),
    .Y(_12935_));
 AOI21x1_ASAP7_75t_R _33236_ (.A1(_12840_),
    .A2(_12935_),
    .B(_12924_),
    .Y(_12936_));
 TAPCELL_ASAP7_75t_R PHY_44 ();
 AND2x2_ASAP7_75t_R _33238_ (.A(_12919_),
    .B(_12904_),
    .Y(_12938_));
 OR3x1_ASAP7_75t_R _33239_ (.A(_12823_),
    .B(_12936_),
    .C(_12938_),
    .Y(_12939_));
 OA211x2_ASAP7_75t_R _33240_ (.A1(_12814_),
    .A2(_12930_),
    .B(_12932_),
    .C(_12939_),
    .Y(_12940_));
 OR4x1_ASAP7_75t_R _33241_ (.A(net254),
    .B(_12918_),
    .C(_12929_),
    .D(_12940_),
    .Y(_12941_));
 OA21x2_ASAP7_75t_R _33242_ (.A1(_14837_),
    .A2(_06686_),
    .B(_12941_),
    .Y(_04370_));
 TAPCELL_ASAP7_75t_R PHY_43 ();
 AND3x1_ASAP7_75t_R _33244_ (.A(_12914_),
    .B(_12919_),
    .C(_12840_),
    .Y(_12943_));
 TAPCELL_ASAP7_75t_R PHY_42 ();
 OA211x2_ASAP7_75t_R _33246_ (.A1(_12823_),
    .A2(_12943_),
    .B(_06686_),
    .C(_12926_),
    .Y(_12945_));
 AOI21x1_ASAP7_75t_R _33247_ (.A1(_01746_),
    .A2(net254),
    .B(_12945_),
    .Y(_04471_));
 TAPCELL_ASAP7_75t_R PHY_41 ();
 AOI21x1_ASAP7_75t_R _33249_ (.A1(_00240_),
    .A2(_12820_),
    .B(_12822_),
    .Y(_12947_));
 AND3x4_ASAP7_75t_R _33250_ (.A(_12947_),
    .B(_12919_),
    .C(_12840_),
    .Y(_12948_));
 TAPCELL_ASAP7_75t_R PHY_40 ();
 AND2x6_ASAP7_75t_R _33252_ (.A(_12800_),
    .B(_12807_),
    .Y(_12950_));
 AND3x4_ASAP7_75t_R _33253_ (.A(_12814_),
    .B(_12948_),
    .C(_12950_),
    .Y(_12951_));
 AO21x2_ASAP7_75t_R _33254_ (.A1(_12919_),
    .A2(_12840_),
    .B(_12823_),
    .Y(_12952_));
 AND2x2_ASAP7_75t_R _33255_ (.A(_12926_),
    .B(_12952_),
    .Y(_12953_));
 AO21x1_ASAP7_75t_R _33256_ (.A1(_12724_),
    .A2(_12951_),
    .B(_12953_),
    .Y(_12954_));
 AND3x1_ASAP7_75t_R _33257_ (.A(_06686_),
    .B(_12914_),
    .C(_12954_),
    .Y(_12955_));
 AOI21x1_ASAP7_75t_R _33258_ (.A1(_00163_),
    .A2(net254),
    .B(_12955_),
    .Y(_04472_));
 INVx1_ASAP7_75t_R _33259_ (.A(_12923_),
    .Y(_12956_));
 NAND2x2_ASAP7_75t_R _33260_ (.A(_12787_),
    .B(_12956_),
    .Y(_12957_));
 AND2x4_ASAP7_75t_R _33261_ (.A(_12823_),
    .B(_12919_),
    .Y(_12958_));
 AO21x2_ASAP7_75t_R _33262_ (.A1(_12912_),
    .A2(_12957_),
    .B(_12958_),
    .Y(_12959_));
 AO21x1_ASAP7_75t_R _33263_ (.A1(_12742_),
    .A2(_12951_),
    .B(_12959_),
    .Y(_12960_));
 TAPCELL_ASAP7_75t_R PHY_39 ();
 AND2x2_ASAP7_75t_R _33265_ (.A(_12948_),
    .B(_12911_),
    .Y(_12962_));
 NOR2x1_ASAP7_75t_R _33266_ (.A(_12903_),
    .B(_12924_),
    .Y(_12963_));
 INVx1_ASAP7_75t_R _33267_ (.A(_12963_),
    .Y(_12964_));
 TAPCELL_ASAP7_75t_R PHY_38 ();
 NAND2x2_ASAP7_75t_R _33269_ (.A(_12926_),
    .B(_12947_),
    .Y(_12966_));
 AO22x2_ASAP7_75t_R _33270_ (.A1(_12927_),
    .A2(_12952_),
    .B1(_12966_),
    .B2(_12733_),
    .Y(_12967_));
 AO32x1_ASAP7_75t_R _33271_ (.A1(_12932_),
    .A2(_12962_),
    .A3(_12964_),
    .B1(_12967_),
    .B2(_12742_),
    .Y(_12968_));
 AO21x1_ASAP7_75t_R _33272_ (.A1(_12915_),
    .A2(_12960_),
    .B(_12968_),
    .Y(_12969_));
 AO21x1_ASAP7_75t_R _33273_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13496_),
    .Y(_12970_));
 OA21x2_ASAP7_75t_R _33274_ (.A1(net254),
    .A2(_12969_),
    .B(_12970_),
    .Y(_04473_));
 AND4x1_ASAP7_75t_R _33275_ (.A(_12814_),
    .B(_12915_),
    .C(_12921_),
    .D(_12950_),
    .Y(_12971_));
 OR2x2_ASAP7_75t_R _33276_ (.A(_12967_),
    .B(_12971_),
    .Y(_12972_));
 AO221x1_ASAP7_75t_R _33277_ (.A1(_12915_),
    .A2(_12958_),
    .B1(_12972_),
    .B2(_12750_),
    .C(net254),
    .Y(_12973_));
 OA21x2_ASAP7_75t_R _33278_ (.A1(_13480_),
    .A2(_06686_),
    .B(_12973_),
    .Y(_04474_));
 TAPCELL_ASAP7_75t_R PHY_37 ();
 NAND2x2_ASAP7_75t_R _33280_ (.A(_12814_),
    .B(_12950_),
    .Y(_12975_));
 OR3x1_ASAP7_75t_R _33281_ (.A(_12757_),
    .B(_12904_),
    .C(_12975_),
    .Y(_12976_));
 AND2x4_ASAP7_75t_R _33282_ (.A(_12832_),
    .B(_12840_),
    .Y(_12977_));
 OR2x2_ASAP7_75t_R _33283_ (.A(_12958_),
    .B(_12977_),
    .Y(_12978_));
 INVx1_ASAP7_75t_R _33284_ (.A(_12978_),
    .Y(_12979_));
 AND3x4_ASAP7_75t_R _33285_ (.A(_12947_),
    .B(_12919_),
    .C(_12904_),
    .Y(_12980_));
 TAPCELL_ASAP7_75t_R PHY_36 ();
 AO21x1_ASAP7_75t_R _33287_ (.A1(_12927_),
    .A2(_12980_),
    .B(_12757_),
    .Y(_12982_));
 NAND2x1_ASAP7_75t_R _33288_ (.A(_12947_),
    .B(_12832_),
    .Y(_12983_));
 AO21x1_ASAP7_75t_R _33289_ (.A1(_12927_),
    .A2(_12983_),
    .B(_12845_),
    .Y(_12984_));
 AO32x1_ASAP7_75t_R _33290_ (.A1(_12915_),
    .A2(_12976_),
    .A3(_12979_),
    .B1(_12982_),
    .B2(_12984_),
    .Y(_12985_));
 TAPCELL_ASAP7_75t_R PHY_35 ();
 OR3x1_ASAP7_75t_R _33292_ (.A(_12904_),
    .B(_12910_),
    .C(_12963_),
    .Y(_12987_));
 AO21x1_ASAP7_75t_R _33293_ (.A1(_12947_),
    .A2(_12987_),
    .B(_12757_),
    .Y(_12988_));
 AND3x1_ASAP7_75t_R _33294_ (.A(_12932_),
    .B(_12983_),
    .C(_12988_),
    .Y(_12989_));
 OR3x1_ASAP7_75t_R _33295_ (.A(net254),
    .B(_12985_),
    .C(_12989_),
    .Y(_12990_));
 OA21x2_ASAP7_75t_R _33296_ (.A1(_13460_),
    .A2(_06686_),
    .B(_12990_),
    .Y(_04475_));
 TAPCELL_ASAP7_75t_R PHY_34 ();
 AND2x4_ASAP7_75t_R _33298_ (.A(_12912_),
    .B(_12957_),
    .Y(_12992_));
 OA211x2_ASAP7_75t_R _33299_ (.A1(_12764_),
    .A2(_12903_),
    .B(_12948_),
    .C(_12950_),
    .Y(_12993_));
 OR3x1_ASAP7_75t_R _33300_ (.A(_12992_),
    .B(_12978_),
    .C(_12993_),
    .Y(_12994_));
 NAND2x2_ASAP7_75t_R _33301_ (.A(_12947_),
    .B(_12904_),
    .Y(_12995_));
 AO22x1_ASAP7_75t_R _33302_ (.A1(_12764_),
    .A2(_12845_),
    .B1(_12995_),
    .B2(_12926_),
    .Y(_12996_));
 NAND2x1_ASAP7_75t_R _33303_ (.A(_12914_),
    .B(_12919_),
    .Y(_12997_));
 AO21x1_ASAP7_75t_R _33304_ (.A1(_12947_),
    .A2(_12997_),
    .B(_12764_),
    .Y(_12998_));
 AO221x1_ASAP7_75t_R _33305_ (.A1(_12915_),
    .A2(_12994_),
    .B1(_12996_),
    .B2(_12998_),
    .C(net254),
    .Y(_12999_));
 OA21x2_ASAP7_75t_R _33306_ (.A1(_13456_),
    .A2(_06686_),
    .B(_12999_),
    .Y(_04476_));
 AO21x1_ASAP7_75t_R _33307_ (.A1(_12771_),
    .A2(_12823_),
    .B(_12962_),
    .Y(_13000_));
 NAND2x1_ASAP7_75t_R _33308_ (.A(_12724_),
    .B(_12914_),
    .Y(_13001_));
 AO21x1_ASAP7_75t_R _33309_ (.A1(_12914_),
    .A2(_12952_),
    .B(_12724_),
    .Y(_13002_));
 OA211x2_ASAP7_75t_R _33310_ (.A1(_13001_),
    .A2(_12951_),
    .B(_13002_),
    .C(_12771_),
    .Y(_13003_));
 AO221x1_ASAP7_75t_R _33311_ (.A1(_12915_),
    .A2(_12978_),
    .B1(_13000_),
    .B2(_12932_),
    .C(_13003_),
    .Y(_13004_));
 AO21x1_ASAP7_75t_R _33312_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13479_),
    .Y(_13005_));
 OA21x2_ASAP7_75t_R _33313_ (.A1(net254),
    .A2(_13004_),
    .B(_13005_),
    .Y(_04477_));
 AO21x1_ASAP7_75t_R _33314_ (.A1(_12926_),
    .A2(_12948_),
    .B(_12780_),
    .Y(_13006_));
 AND3x1_ASAP7_75t_R _33315_ (.A(_12814_),
    .B(_12911_),
    .C(_12924_),
    .Y(_13007_));
 AO21x1_ASAP7_75t_R _33316_ (.A1(_12780_),
    .A2(_12934_),
    .B(_13007_),
    .Y(_13008_));
 OR3x1_ASAP7_75t_R _33317_ (.A(_12724_),
    .B(_12823_),
    .C(_12904_),
    .Y(_13009_));
 AO21x1_ASAP7_75t_R _33318_ (.A1(_12919_),
    .A2(_13008_),
    .B(_13009_),
    .Y(_13010_));
 AND3x1_ASAP7_75t_R _33319_ (.A(_12733_),
    .B(_13006_),
    .C(_13010_),
    .Y(_13011_));
 TAPCELL_ASAP7_75t_R PHY_33 ();
 AO32x1_ASAP7_75t_R _33321_ (.A1(_12742_),
    .A2(_12947_),
    .A3(_12904_),
    .B1(_12952_),
    .B2(_12780_),
    .Y(_13013_));
 AND2x2_ASAP7_75t_R _33322_ (.A(_12947_),
    .B(_12919_),
    .Y(_13014_));
 OA21x2_ASAP7_75t_R _33323_ (.A1(_12904_),
    .A2(_13014_),
    .B(_12780_),
    .Y(_13015_));
 AO221x1_ASAP7_75t_R _33324_ (.A1(_12823_),
    .A2(_12938_),
    .B1(_12977_),
    .B2(_12814_),
    .C(_13015_),
    .Y(_13016_));
 AO22x1_ASAP7_75t_R _33325_ (.A1(_12927_),
    .A2(_13013_),
    .B1(_13016_),
    .B2(_12915_),
    .Y(_13017_));
 OR3x1_ASAP7_75t_R _33326_ (.A(net254),
    .B(_13011_),
    .C(_13017_),
    .Y(_13018_));
 OA21x2_ASAP7_75t_R _33327_ (.A1(_13890_),
    .A2(_06686_),
    .B(_13018_),
    .Y(_04478_));
 AO32x1_ASAP7_75t_R _33328_ (.A1(_12750_),
    .A2(_12832_),
    .A3(_12840_),
    .B1(_13014_),
    .B2(_12787_),
    .Y(_13019_));
 AO32x1_ASAP7_75t_R _33329_ (.A1(_12750_),
    .A2(_12947_),
    .A3(_12904_),
    .B1(_12952_),
    .B2(_12787_),
    .Y(_13020_));
 AO32x1_ASAP7_75t_R _33330_ (.A1(_12915_),
    .A2(_12930_),
    .A3(_13019_),
    .B1(_13020_),
    .B2(_12927_),
    .Y(_13021_));
 NAND2x1_ASAP7_75t_R _33331_ (.A(_12823_),
    .B(_12919_),
    .Y(_13022_));
 AO21x1_ASAP7_75t_R _33332_ (.A1(_12904_),
    .A2(_13022_),
    .B(_12733_),
    .Y(_13023_));
 NAND2x1_ASAP7_75t_R _33333_ (.A(_12947_),
    .B(_12840_),
    .Y(_13024_));
 AO21x1_ASAP7_75t_R _33334_ (.A1(_12948_),
    .A2(_12934_),
    .B(_13024_),
    .Y(_13025_));
 AO21x1_ASAP7_75t_R _33335_ (.A1(_12733_),
    .A2(_13025_),
    .B(_12724_),
    .Y(_13026_));
 AND3x1_ASAP7_75t_R _33336_ (.A(_12787_),
    .B(_13023_),
    .C(_13026_),
    .Y(_13027_));
 OR3x1_ASAP7_75t_R _33337_ (.A(_09319_),
    .B(_13021_),
    .C(_13027_),
    .Y(_13028_));
 OA21x2_ASAP7_75t_R _33338_ (.A1(_05658_),
    .A2(_06686_),
    .B(_13028_),
    .Y(_04479_));
 INVx1_ASAP7_75t_R _33339_ (.A(_13014_),
    .Y(_13029_));
 OR3x1_ASAP7_75t_R _33340_ (.A(_12724_),
    .B(_13029_),
    .C(_12910_),
    .Y(_13030_));
 OA21x2_ASAP7_75t_R _33341_ (.A1(_12733_),
    .A2(_12919_),
    .B(_13030_),
    .Y(_13031_));
 OR3x1_ASAP7_75t_R _33342_ (.A(_12757_),
    .B(_12904_),
    .C(_13031_),
    .Y(_13032_));
 AO21x1_ASAP7_75t_R _33343_ (.A1(_12724_),
    .A2(_13022_),
    .B(_12733_),
    .Y(_13033_));
 AO21x1_ASAP7_75t_R _33344_ (.A1(_12914_),
    .A2(_12977_),
    .B(_12794_),
    .Y(_13034_));
 AND3x1_ASAP7_75t_R _33345_ (.A(_13032_),
    .B(_13033_),
    .C(_13034_),
    .Y(_13035_));
 OR2x2_ASAP7_75t_R _33346_ (.A(_12757_),
    .B(_12840_),
    .Y(_13036_));
 OR3x1_ASAP7_75t_R _33347_ (.A(_12771_),
    .B(_12919_),
    .C(_12904_),
    .Y(_13037_));
 AO21x1_ASAP7_75t_R _33348_ (.A1(_13036_),
    .A2(_13037_),
    .B(_12823_),
    .Y(_13038_));
 OA211x2_ASAP7_75t_R _33349_ (.A1(_12794_),
    .A2(_12922_),
    .B(_13038_),
    .C(_12927_),
    .Y(_13039_));
 OR3x1_ASAP7_75t_R _33350_ (.A(net254),
    .B(_13035_),
    .C(_13039_),
    .Y(_13040_));
 OA21x2_ASAP7_75t_R _33351_ (.A1(_14176_),
    .A2(_06686_),
    .B(_13040_),
    .Y(_04480_));
 OR3x1_ASAP7_75t_R _33352_ (.A(_12757_),
    .B(_12905_),
    .C(_12910_),
    .Y(_13041_));
 OA21x2_ASAP7_75t_R _33353_ (.A1(_12733_),
    .A2(_13022_),
    .B(_12724_),
    .Y(_13042_));
 AO21x1_ASAP7_75t_R _33354_ (.A1(_12733_),
    .A2(_13041_),
    .B(_13042_),
    .Y(_13043_));
 AND2x2_ASAP7_75t_R _33355_ (.A(_12947_),
    .B(_12904_),
    .Y(_13044_));
 OR3x1_ASAP7_75t_R _33356_ (.A(_12724_),
    .B(_12800_),
    .C(_13044_),
    .Y(_13045_));
 OA21x2_ASAP7_75t_R _33357_ (.A1(_12926_),
    .A2(_12948_),
    .B(_13045_),
    .Y(_13046_));
 AO221x1_ASAP7_75t_R _33358_ (.A1(_12800_),
    .A2(_13043_),
    .B1(_13046_),
    .B2(_12914_),
    .C(net254),
    .Y(_13047_));
 OA21x2_ASAP7_75t_R _33359_ (.A1(_14182_),
    .A2(_06686_),
    .B(_13047_),
    .Y(_04481_));
 AO21x1_ASAP7_75t_R _33360_ (.A1(_12807_),
    .A2(_12980_),
    .B(_12951_),
    .Y(_13048_));
 AND3x1_ASAP7_75t_R _33361_ (.A(_12926_),
    .B(_12807_),
    .C(_12995_),
    .Y(_13049_));
 AO21x1_ASAP7_75t_R _33362_ (.A1(_12724_),
    .A2(_13048_),
    .B(_13049_),
    .Y(_13050_));
 AO22x1_ASAP7_75t_R _33363_ (.A1(_12733_),
    .A2(_13041_),
    .B1(_12997_),
    .B2(_12724_),
    .Y(_13051_));
 AO221x1_ASAP7_75t_R _33364_ (.A1(_12914_),
    .A2(_13050_),
    .B1(_13051_),
    .B2(_12807_),
    .C(net254),
    .Y(_13052_));
 OA21x2_ASAP7_75t_R _33365_ (.A1(_14293_),
    .A2(_06686_),
    .B(_13052_),
    .Y(_04482_));
 AO21x1_ASAP7_75t_R _33366_ (.A1(_12814_),
    .A2(_12919_),
    .B(_12977_),
    .Y(_13053_));
 NAND2x1_ASAP7_75t_R _33367_ (.A(_12800_),
    .B(_12807_),
    .Y(_13054_));
 AO21x1_ASAP7_75t_R _33368_ (.A1(_12764_),
    .A2(_12771_),
    .B(_12814_),
    .Y(_13055_));
 OR2x2_ASAP7_75t_R _33369_ (.A(_13054_),
    .B(_13055_),
    .Y(_13056_));
 AO221x1_ASAP7_75t_R _33370_ (.A1(_12823_),
    .A2(_13053_),
    .B1(_13056_),
    .B2(_12948_),
    .C(_12733_),
    .Y(_13057_));
 AO21x1_ASAP7_75t_R _33371_ (.A1(_12742_),
    .A2(_12992_),
    .B(_13057_),
    .Y(_13058_));
 OA21x2_ASAP7_75t_R _33372_ (.A1(_12914_),
    .A2(_12814_),
    .B(_12724_),
    .Y(_13059_));
 INVx1_ASAP7_75t_R _33373_ (.A(_12966_),
    .Y(_13060_));
 AND2x2_ASAP7_75t_R _33374_ (.A(_12814_),
    .B(_12823_),
    .Y(_13061_));
 AO21x1_ASAP7_75t_R _33375_ (.A1(_12938_),
    .A2(_13060_),
    .B(_13061_),
    .Y(_13062_));
 OA211x2_ASAP7_75t_R _33376_ (.A1(_12823_),
    .A2(_12943_),
    .B(_12926_),
    .C(_12814_),
    .Y(_13063_));
 AO221x1_ASAP7_75t_R _33377_ (.A1(_13058_),
    .A2(_13059_),
    .B1(_13062_),
    .B2(_12733_),
    .C(_13063_),
    .Y(_13064_));
 AO21x1_ASAP7_75t_R _33378_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13483_),
    .Y(_13065_));
 OA21x2_ASAP7_75t_R _33379_ (.A1(net254),
    .A2(_13064_),
    .B(_13065_),
    .Y(_04483_));
 AO21x1_ASAP7_75t_R _33380_ (.A1(_12919_),
    .A2(_13061_),
    .B(_12733_),
    .Y(_13066_));
 AO21x1_ASAP7_75t_R _33381_ (.A1(_12771_),
    .A2(_12903_),
    .B(_13061_),
    .Y(_13067_));
 OA211x2_ASAP7_75t_R _33382_ (.A1(_12906_),
    .A2(_13067_),
    .B(_12948_),
    .C(_12807_),
    .Y(_13068_));
 AOI211x1_ASAP7_75t_R _33383_ (.A1(_12750_),
    .A2(_12992_),
    .B(_13066_),
    .C(_13068_),
    .Y(_13069_));
 AND2x2_ASAP7_75t_R _33384_ (.A(_12733_),
    .B(_12947_),
    .Y(_13070_));
 OR3x1_ASAP7_75t_R _33385_ (.A(_12926_),
    .B(_13069_),
    .C(_13070_),
    .Y(_13071_));
 OA211x2_ASAP7_75t_R _33386_ (.A1(_12724_),
    .A2(_13014_),
    .B(_13071_),
    .C(_06686_),
    .Y(_13072_));
 AOI21x1_ASAP7_75t_R _33387_ (.A1(_00282_),
    .A2(net254),
    .B(_13072_),
    .Y(_04484_));
 AO21x1_ASAP7_75t_R _33388_ (.A1(_12903_),
    .A2(_12909_),
    .B(_13054_),
    .Y(_13073_));
 AO221x1_ASAP7_75t_R _33389_ (.A1(_12757_),
    .A2(_12992_),
    .B1(_13073_),
    .B2(_12948_),
    .C(_13066_),
    .Y(_13074_));
 OA211x2_ASAP7_75t_R _33390_ (.A1(_12914_),
    .A2(_12832_),
    .B(_13074_),
    .C(_12724_),
    .Y(_13075_));
 AND3x1_ASAP7_75t_R _33391_ (.A(_12926_),
    .B(_12823_),
    .C(_12832_),
    .Y(_13076_));
 OR3x1_ASAP7_75t_R _33392_ (.A(net254),
    .B(_13075_),
    .C(_13076_),
    .Y(_13077_));
 OA21x2_ASAP7_75t_R _33393_ (.A1(_13570_),
    .A2(_06686_),
    .B(_13077_),
    .Y(_04485_));
 AND2x2_ASAP7_75t_R _33394_ (.A(_12947_),
    .B(_12832_),
    .Y(_13078_));
 AO32x1_ASAP7_75t_R _33395_ (.A1(_12780_),
    .A2(_12927_),
    .A3(_13078_),
    .B1(_12984_),
    .B2(_12840_),
    .Y(_13079_));
 AO21x1_ASAP7_75t_R _33396_ (.A1(_12948_),
    .A2(_12950_),
    .B(_12958_),
    .Y(_13080_));
 AND3x1_ASAP7_75t_R _33397_ (.A(_12764_),
    .B(_12771_),
    .C(_12903_),
    .Y(_13081_));
 AOI21x1_ASAP7_75t_R _33398_ (.A1(_12950_),
    .A2(_13055_),
    .B(_12905_),
    .Y(_13082_));
 OR3x1_ASAP7_75t_R _33399_ (.A(_12980_),
    .B(_12977_),
    .C(_13082_),
    .Y(_13083_));
 AO21x1_ASAP7_75t_R _33400_ (.A1(_12948_),
    .A2(_13081_),
    .B(_13083_),
    .Y(_13084_));
 AO222x2_ASAP7_75t_R _33401_ (.A1(_12764_),
    .A2(_12992_),
    .B1(_13080_),
    .B2(_12814_),
    .C1(_13084_),
    .C2(_12780_),
    .Y(_13085_));
 OA21x2_ASAP7_75t_R _33402_ (.A1(_12814_),
    .A2(_12911_),
    .B(_12948_),
    .Y(_13086_));
 OA21x2_ASAP7_75t_R _33403_ (.A1(_12980_),
    .A2(_13086_),
    .B(_12780_),
    .Y(_13087_));
 AO21x1_ASAP7_75t_R _33404_ (.A1(_12823_),
    .A2(_12840_),
    .B(_13087_),
    .Y(_13088_));
 AO22x1_ASAP7_75t_R _33405_ (.A1(_12915_),
    .A2(_13085_),
    .B1(_13088_),
    .B2(_12932_),
    .Y(_13089_));
 OR3x1_ASAP7_75t_R _33406_ (.A(net254),
    .B(_13079_),
    .C(_13089_),
    .Y(_13090_));
 OA21x2_ASAP7_75t_R _33407_ (.A1(_13649_),
    .A2(_06686_),
    .B(_13090_),
    .Y(_04486_));
 OR3x1_ASAP7_75t_R _33408_ (.A(_12814_),
    .B(_12905_),
    .C(_12911_),
    .Y(_13091_));
 AO21x1_ASAP7_75t_R _33409_ (.A1(_12787_),
    .A2(_13091_),
    .B(_13029_),
    .Y(_13092_));
 AND2x2_ASAP7_75t_R _33410_ (.A(_00240_),
    .B(net2692),
    .Y(_13093_));
 AO21x1_ASAP7_75t_R _33411_ (.A1(_06589_),
    .A2(_12517_),
    .B(_13093_),
    .Y(_13094_));
 NAND2x1_ASAP7_75t_R _33412_ (.A(_06734_),
    .B(_01813_),
    .Y(_13095_));
 OA211x2_ASAP7_75t_R _33413_ (.A1(net2688),
    .A2(_06734_),
    .B(_13095_),
    .C(_06580_),
    .Y(_13096_));
 AOI21x1_ASAP7_75t_R _33414_ (.A1(net431),
    .A2(_13094_),
    .B(_13096_),
    .Y(_13097_));
 INVx1_ASAP7_75t_R _33415_ (.A(_13097_),
    .Y(_13098_));
 OA21x2_ASAP7_75t_R _33416_ (.A1(_12787_),
    .A2(_12983_),
    .B(_12914_),
    .Y(_13099_));
 OA21x2_ASAP7_75t_R _33417_ (.A1(_12922_),
    .A2(_13098_),
    .B(_13099_),
    .Y(_13100_));
 AO21x1_ASAP7_75t_R _33418_ (.A1(_13070_),
    .A2(_13092_),
    .B(_13100_),
    .Y(_13101_));
 NAND2x1_ASAP7_75t_R _33419_ (.A(_12733_),
    .B(_13097_),
    .Y(_13102_));
 OR3x2_ASAP7_75t_R _33420_ (.A(_12764_),
    .B(_12771_),
    .C(_12814_),
    .Y(_13103_));
 AO32x1_ASAP7_75t_R _33421_ (.A1(_12814_),
    .A2(_12950_),
    .A3(_13098_),
    .B1(_13081_),
    .B2(_12787_),
    .Y(_13104_));
 AND3x1_ASAP7_75t_R _33422_ (.A(_12948_),
    .B(_13103_),
    .C(_13104_),
    .Y(_13105_));
 INVx1_ASAP7_75t_R _33423_ (.A(_12957_),
    .Y(_13106_));
 OA21x2_ASAP7_75t_R _33424_ (.A1(_12771_),
    .A2(_13106_),
    .B(_12912_),
    .Y(_13107_));
 OR3x1_ASAP7_75t_R _33425_ (.A(_13066_),
    .B(_13105_),
    .C(_13107_),
    .Y(_13108_));
 AO21x1_ASAP7_75t_R _33426_ (.A1(_12787_),
    .A2(_13083_),
    .B(_13108_),
    .Y(_13109_));
 AO22x1_ASAP7_75t_R _33427_ (.A1(_12733_),
    .A2(_13092_),
    .B1(_13109_),
    .B2(_12724_),
    .Y(_13110_));
 AO221x1_ASAP7_75t_R _33428_ (.A1(_12926_),
    .A2(_13101_),
    .B1(_13102_),
    .B2(_13110_),
    .C(net254),
    .Y(_13111_));
 OA21x2_ASAP7_75t_R _33429_ (.A1(_13675_),
    .A2(_06686_),
    .B(_13111_),
    .Y(_04487_));
 NAND2x1_ASAP7_75t_R _33430_ (.A(_12565_),
    .B(_00239_),
    .Y(_13112_));
 OA21x2_ASAP7_75t_R _33431_ (.A1(_00239_),
    .A2(_12485_),
    .B(_13112_),
    .Y(_13113_));
 NAND2x1_ASAP7_75t_R _33432_ (.A(_06589_),
    .B(_01829_),
    .Y(_13114_));
 OA211x2_ASAP7_75t_R _33433_ (.A1(_06589_),
    .A2(net2625),
    .B(_13114_),
    .C(net431),
    .Y(_13115_));
 AO21x1_ASAP7_75t_R _33434_ (.A1(_06580_),
    .A2(_13113_),
    .B(_13115_),
    .Y(_13116_));
 AO32x1_ASAP7_75t_R _33435_ (.A1(_12794_),
    .A2(_12947_),
    .A3(_12832_),
    .B1(_12952_),
    .B2(_13116_),
    .Y(_13117_));
 AO22x1_ASAP7_75t_R _33436_ (.A1(_12845_),
    .A2(_13116_),
    .B1(_13117_),
    .B2(_12927_),
    .Y(_13118_));
 AO221x1_ASAP7_75t_R _33437_ (.A1(_12794_),
    .A2(_13086_),
    .B1(_13116_),
    .B2(_12823_),
    .C(_12980_),
    .Y(_13119_));
 AND2x2_ASAP7_75t_R _33438_ (.A(_12932_),
    .B(_13119_),
    .Y(_13120_));
 AO22x1_ASAP7_75t_R _33439_ (.A1(_12814_),
    .A2(_12959_),
    .B1(_13116_),
    .B2(_12951_),
    .Y(_13121_));
 OA21x2_ASAP7_75t_R _33440_ (.A1(_13120_),
    .A2(_13121_),
    .B(_12930_),
    .Y(_13122_));
 OA21x2_ASAP7_75t_R _33441_ (.A1(_13084_),
    .A2(_13121_),
    .B(_12915_),
    .Y(_13123_));
 OA22x2_ASAP7_75t_R _33442_ (.A1(_12794_),
    .A2(_13122_),
    .B1(_13123_),
    .B2(_13120_),
    .Y(_13124_));
 OR3x1_ASAP7_75t_R _33443_ (.A(_09319_),
    .B(_13118_),
    .C(_13124_),
    .Y(_13125_));
 OA21x2_ASAP7_75t_R _33444_ (.A1(_13630_),
    .A2(_06686_),
    .B(_13125_),
    .Y(_04488_));
 NAND2x1_ASAP7_75t_R _33445_ (.A(_12570_),
    .B(_00239_),
    .Y(_13126_));
 OA21x2_ASAP7_75t_R _33446_ (.A1(_00239_),
    .A2(_12487_),
    .B(_13126_),
    .Y(_13127_));
 NAND2x1_ASAP7_75t_R _33447_ (.A(_06589_),
    .B(_01828_),
    .Y(_13128_));
 OA211x2_ASAP7_75t_R _33448_ (.A1(_06589_),
    .A2(net2618),
    .B(_13128_),
    .C(net431),
    .Y(_13129_));
 AO21x2_ASAP7_75t_R _33449_ (.A1(_06580_),
    .A2(_13127_),
    .B(_13129_),
    .Y(_13130_));
 AO21x1_ASAP7_75t_R _33450_ (.A1(_12995_),
    .A2(_13130_),
    .B(_13078_),
    .Y(_13131_));
 AO221x1_ASAP7_75t_R _33451_ (.A1(_12800_),
    .A2(_13086_),
    .B1(_13130_),
    .B2(_12823_),
    .C(_12980_),
    .Y(_13132_));
 OR3x1_ASAP7_75t_R _33452_ (.A(_12904_),
    .B(_12975_),
    .C(_13130_),
    .Y(_13133_));
 AO221x1_ASAP7_75t_R _33453_ (.A1(_12814_),
    .A2(_12959_),
    .B1(_13133_),
    .B2(_13014_),
    .C(_12977_),
    .Y(_13134_));
 AO22x1_ASAP7_75t_R _33454_ (.A1(_12932_),
    .A2(_13132_),
    .B1(_13134_),
    .B2(_12915_),
    .Y(_13135_));
 OA21x2_ASAP7_75t_R _33455_ (.A1(_12800_),
    .A2(_12930_),
    .B(_13135_),
    .Y(_13136_));
 AO21x1_ASAP7_75t_R _33456_ (.A1(_12733_),
    .A2(_13130_),
    .B(_13136_),
    .Y(_13137_));
 AO222x2_ASAP7_75t_R _33457_ (.A1(_12927_),
    .A2(_13131_),
    .B1(_13136_),
    .B2(_12733_),
    .C1(_12724_),
    .C2(_13137_),
    .Y(_13138_));
 AO21x1_ASAP7_75t_R _33458_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13636_),
    .Y(_13139_));
 OA21x2_ASAP7_75t_R _33459_ (.A1(net254),
    .A2(_13138_),
    .B(_13139_),
    .Y(_04489_));
 TAPCELL_ASAP7_75t_R PHY_32 ();
 AND2x2_ASAP7_75t_R _33461_ (.A(net428),
    .B(net2652),
    .Y(_13141_));
 AO21x1_ASAP7_75t_R _33462_ (.A1(_06589_),
    .A2(_12524_),
    .B(_13141_),
    .Y(_13142_));
 TAPCELL_ASAP7_75t_R PHY_31 ();
 NAND2x1_ASAP7_75t_R _33464_ (.A(_06734_),
    .B(_01810_),
    .Y(_13144_));
 OA211x2_ASAP7_75t_R _33465_ (.A1(net2670),
    .A2(_06734_),
    .B(_13144_),
    .C(_06580_),
    .Y(_13145_));
 AO21x1_ASAP7_75t_R _33466_ (.A1(net431),
    .A2(_13142_),
    .B(_13145_),
    .Y(_13146_));
 AO21x1_ASAP7_75t_R _33467_ (.A1(_12927_),
    .A2(_12952_),
    .B(_12845_),
    .Y(_13147_));
 AO221x1_ASAP7_75t_R _33468_ (.A1(_12807_),
    .A2(_13086_),
    .B1(_13146_),
    .B2(_12823_),
    .C(_12980_),
    .Y(_13148_));
 AO21x1_ASAP7_75t_R _33469_ (.A1(_12814_),
    .A2(_12959_),
    .B(_12980_),
    .Y(_13149_));
 AO21x1_ASAP7_75t_R _33470_ (.A1(_12951_),
    .A2(_13146_),
    .B(_13149_),
    .Y(_13150_));
 AO22x1_ASAP7_75t_R _33471_ (.A1(_12932_),
    .A2(_13148_),
    .B1(_13150_),
    .B2(_12915_),
    .Y(_13151_));
 OR2x2_ASAP7_75t_R _33472_ (.A(_12807_),
    .B(_12930_),
    .Y(_13152_));
 AO221x1_ASAP7_75t_R _33473_ (.A1(_13146_),
    .A2(_13147_),
    .B1(_13151_),
    .B2(_13152_),
    .C(_09319_),
    .Y(_13153_));
 OA21x2_ASAP7_75t_R _33474_ (.A1(_13626_),
    .A2(_06686_),
    .B(_13153_),
    .Y(_04490_));
 AO21x1_ASAP7_75t_R _33475_ (.A1(_12911_),
    .A2(_12963_),
    .B(_12904_),
    .Y(_13154_));
 AO22x1_ASAP7_75t_R _33476_ (.A1(_12742_),
    .A2(_12840_),
    .B1(_13154_),
    .B2(_12919_),
    .Y(_13155_));
 AND2x2_ASAP7_75t_R _33477_ (.A(net428),
    .B(net2772),
    .Y(_13156_));
 AO21x1_ASAP7_75t_R _33478_ (.A1(_06589_),
    .A2(_12527_),
    .B(_13156_),
    .Y(_13157_));
 NAND2x1_ASAP7_75t_R _33479_ (.A(_06734_),
    .B(_01809_),
    .Y(_13158_));
 OA211x2_ASAP7_75t_R _33480_ (.A1(net2801),
    .A2(_06734_),
    .B(_13158_),
    .C(_06580_),
    .Y(_13159_));
 AO21x1_ASAP7_75t_R _33481_ (.A1(net431),
    .A2(_13157_),
    .B(_13159_),
    .Y(_13160_));
 AND2x2_ASAP7_75t_R _33482_ (.A(_12823_),
    .B(_13160_),
    .Y(_13161_));
 AO21x1_ASAP7_75t_R _33483_ (.A1(_12947_),
    .A2(_13155_),
    .B(_13161_),
    .Y(_13162_));
 AND3x2_ASAP7_75t_R _33484_ (.A(_12947_),
    .B(_12832_),
    .C(_12904_),
    .Y(_13163_));
 AO21x1_ASAP7_75t_R _33485_ (.A1(_12948_),
    .A2(_12975_),
    .B(_13163_),
    .Y(_13164_));
 AO221x1_ASAP7_75t_R _33486_ (.A1(_12951_),
    .A2(_13160_),
    .B1(_13164_),
    .B2(_12742_),
    .C(_13149_),
    .Y(_13165_));
 AO22x1_ASAP7_75t_R _33487_ (.A1(_12932_),
    .A2(_13162_),
    .B1(_13165_),
    .B2(_12915_),
    .Y(_13166_));
 OA21x2_ASAP7_75t_R _33488_ (.A1(_12742_),
    .A2(_12930_),
    .B(_13166_),
    .Y(_13167_));
 AO22x1_ASAP7_75t_R _33489_ (.A1(_12742_),
    .A2(_13078_),
    .B1(_13160_),
    .B2(_12919_),
    .Y(_13168_));
 AO21x1_ASAP7_75t_R _33490_ (.A1(_12840_),
    .A2(_13168_),
    .B(_13161_),
    .Y(_13169_));
 AO22x1_ASAP7_75t_R _33491_ (.A1(_12845_),
    .A2(_13160_),
    .B1(_13169_),
    .B2(_12927_),
    .Y(_13170_));
 OR3x1_ASAP7_75t_R _33492_ (.A(_09319_),
    .B(_13167_),
    .C(_13170_),
    .Y(_13171_));
 OA21x2_ASAP7_75t_R _33493_ (.A1(_13376_),
    .A2(_06686_),
    .B(_13171_),
    .Y(_04491_));
 AND2x2_ASAP7_75t_R _33494_ (.A(net428),
    .B(net2599),
    .Y(_13172_));
 AO21x1_ASAP7_75t_R _33495_ (.A1(_06589_),
    .A2(_12530_),
    .B(_13172_),
    .Y(_13173_));
 NAND2x1_ASAP7_75t_R _33496_ (.A(_06734_),
    .B(_01808_),
    .Y(_13174_));
 OA211x2_ASAP7_75t_R _33497_ (.A1(net2603),
    .A2(_06734_),
    .B(_13174_),
    .C(_06580_),
    .Y(_13175_));
 AO21x1_ASAP7_75t_R _33498_ (.A1(net430),
    .A2(_13173_),
    .B(_13175_),
    .Y(_13176_));
 OA211x2_ASAP7_75t_R _33499_ (.A1(_12943_),
    .A2(_12966_),
    .B(_13176_),
    .C(_13001_),
    .Y(_13177_));
 AO21x1_ASAP7_75t_R _33500_ (.A1(_12948_),
    .A2(_13081_),
    .B(_13163_),
    .Y(_13178_));
 AND3x1_ASAP7_75t_R _33501_ (.A(_12814_),
    .B(_12912_),
    .C(_12957_),
    .Y(_13179_));
 AO221x1_ASAP7_75t_R _33502_ (.A1(_12951_),
    .A2(_13176_),
    .B1(_13178_),
    .B2(_12750_),
    .C(_13179_),
    .Y(_13180_));
 AO21x1_ASAP7_75t_R _33503_ (.A1(_12733_),
    .A2(_12919_),
    .B(_12977_),
    .Y(_13181_));
 AO21x1_ASAP7_75t_R _33504_ (.A1(_12919_),
    .A2(_12905_),
    .B(_13082_),
    .Y(_13182_));
 AO32x1_ASAP7_75t_R _33505_ (.A1(_12926_),
    .A2(_12947_),
    .A3(_13181_),
    .B1(_13182_),
    .B2(_12915_),
    .Y(_13183_));
 AO32x1_ASAP7_75t_R _33506_ (.A1(_12915_),
    .A2(_12930_),
    .A3(_13180_),
    .B1(_13183_),
    .B2(_12750_),
    .Y(_13184_));
 OR3x1_ASAP7_75t_R _33507_ (.A(_09319_),
    .B(_13177_),
    .C(_13184_),
    .Y(_13185_));
 OA21x2_ASAP7_75t_R _33508_ (.A1(net2278),
    .A2(_06686_),
    .B(_13185_),
    .Y(_04492_));
 AND2x2_ASAP7_75t_R _33509_ (.A(net428),
    .B(net2629),
    .Y(_13186_));
 AO21x1_ASAP7_75t_R _33510_ (.A1(_06589_),
    .A2(_12532_),
    .B(_13186_),
    .Y(_13187_));
 NAND2x1_ASAP7_75t_R _33511_ (.A(_06734_),
    .B(_01807_),
    .Y(_13188_));
 OA211x2_ASAP7_75t_R _33512_ (.A1(net2614),
    .A2(_06734_),
    .B(_13188_),
    .C(_06580_),
    .Y(_13189_));
 AO21x2_ASAP7_75t_R _33513_ (.A1(net430),
    .A2(_13187_),
    .B(_13189_),
    .Y(_13190_));
 OR3x1_ASAP7_75t_R _33514_ (.A(_12757_),
    .B(_12919_),
    .C(_12904_),
    .Y(_13191_));
 OA21x2_ASAP7_75t_R _33515_ (.A1(_12771_),
    .A2(_12840_),
    .B(_13191_),
    .Y(_13192_));
 OA21x2_ASAP7_75t_R _33516_ (.A1(_12823_),
    .A2(_13192_),
    .B(_13190_),
    .Y(_13193_));
 AO21x1_ASAP7_75t_R _33517_ (.A1(_12922_),
    .A2(_13192_),
    .B(_13193_),
    .Y(_13194_));
 AO22x1_ASAP7_75t_R _33518_ (.A1(_12845_),
    .A2(_13190_),
    .B1(_13194_),
    .B2(_12927_),
    .Y(_13195_));
 OR3x1_ASAP7_75t_R _33519_ (.A(_12757_),
    .B(_12823_),
    .C(_12938_),
    .Y(_13196_));
 OA211x2_ASAP7_75t_R _33520_ (.A1(_12947_),
    .A2(_13190_),
    .B(_13196_),
    .C(_12932_),
    .Y(_13197_));
 OR3x1_ASAP7_75t_R _33521_ (.A(_12958_),
    .B(_13044_),
    .C(_13082_),
    .Y(_13198_));
 AO32x1_ASAP7_75t_R _33522_ (.A1(_12814_),
    .A2(_12950_),
    .A3(_13190_),
    .B1(_13081_),
    .B2(_12757_),
    .Y(_13199_));
 AO221x1_ASAP7_75t_R _33523_ (.A1(_12757_),
    .A2(_13198_),
    .B1(_13199_),
    .B2(_12948_),
    .C(_12980_),
    .Y(_13200_));
 OA21x2_ASAP7_75t_R _33524_ (.A1(_13179_),
    .A2(_13200_),
    .B(_12915_),
    .Y(_13201_));
 OA22x2_ASAP7_75t_R _33525_ (.A1(_12757_),
    .A2(_12930_),
    .B1(_13197_),
    .B2(_13201_),
    .Y(_13202_));
 OR3x1_ASAP7_75t_R _33526_ (.A(_09319_),
    .B(_13195_),
    .C(_13202_),
    .Y(_13203_));
 OA21x2_ASAP7_75t_R _33527_ (.A1(_13350_),
    .A2(_06686_),
    .B(_13203_),
    .Y(_04493_));
 AND4x1_ASAP7_75t_R _33528_ (.A(_12724_),
    .B(_12914_),
    .C(_12919_),
    .D(_13024_),
    .Y(_13204_));
 AO21x1_ASAP7_75t_R _33529_ (.A1(_12926_),
    .A2(_13070_),
    .B(_13204_),
    .Y(_13205_));
 OR2x2_ASAP7_75t_R _33530_ (.A(_12764_),
    .B(_12832_),
    .Y(_13206_));
 OA21x2_ASAP7_75t_R _33531_ (.A1(_12800_),
    .A2(_12919_),
    .B(_13206_),
    .Y(_13207_));
 OA21x2_ASAP7_75t_R _33532_ (.A1(_12995_),
    .A2(_13207_),
    .B(_12927_),
    .Y(_13208_));
 NAND2x1_ASAP7_75t_R _33533_ (.A(_12586_),
    .B(_00239_),
    .Y(_13209_));
 OA21x2_ASAP7_75t_R _33534_ (.A1(_00239_),
    .A2(_12497_),
    .B(_13209_),
    .Y(_13210_));
 NAND2x1_ASAP7_75t_R _33535_ (.A(_06589_),
    .B(_01823_),
    .Y(_13211_));
 OA211x2_ASAP7_75t_R _33536_ (.A1(_06589_),
    .A2(net2641),
    .B(_13211_),
    .C(net431),
    .Y(_13212_));
 AO21x1_ASAP7_75t_R _33537_ (.A1(_06580_),
    .A2(_13210_),
    .B(_13212_),
    .Y(_13213_));
 AO21x1_ASAP7_75t_R _33538_ (.A1(_12922_),
    .A2(_13208_),
    .B(_13213_),
    .Y(_13214_));
 AO21x1_ASAP7_75t_R _33539_ (.A1(_12733_),
    .A2(_12966_),
    .B(_13208_),
    .Y(_13215_));
 OA21x2_ASAP7_75t_R _33540_ (.A1(_12975_),
    .A2(_13213_),
    .B(_12948_),
    .Y(_13216_));
 OA21x2_ASAP7_75t_R _33541_ (.A1(_13163_),
    .A2(_13216_),
    .B(_12764_),
    .Y(_13217_));
 AO221x1_ASAP7_75t_R _33542_ (.A1(_12814_),
    .A2(_12992_),
    .B1(_13216_),
    .B2(_12950_),
    .C(_13217_),
    .Y(_13218_));
 AND2x2_ASAP7_75t_R _33543_ (.A(_12915_),
    .B(_12930_),
    .Y(_13219_));
 AO222x2_ASAP7_75t_R _33544_ (.A1(_12764_),
    .A2(_13205_),
    .B1(_13214_),
    .B2(_13215_),
    .C1(_13218_),
    .C2(_13219_),
    .Y(_13220_));
 AO21x1_ASAP7_75t_R _33545_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13373_),
    .Y(_13221_));
 OA21x2_ASAP7_75t_R _33546_ (.A1(net254),
    .A2(_13220_),
    .B(_13221_),
    .Y(_04494_));
 AND2x2_ASAP7_75t_R _33547_ (.A(net428),
    .B(net2666),
    .Y(_13222_));
 AO21x1_ASAP7_75t_R _33548_ (.A1(_06589_),
    .A2(_12536_),
    .B(_13222_),
    .Y(_13223_));
 NAND2x1_ASAP7_75t_R _33549_ (.A(_06734_),
    .B(_01805_),
    .Y(_13224_));
 OA211x2_ASAP7_75t_R _33550_ (.A1(net2682),
    .A2(_06734_),
    .B(_13224_),
    .C(_06580_),
    .Y(_13225_));
 AO21x1_ASAP7_75t_R _33551_ (.A1(net431),
    .A2(_13223_),
    .B(_13225_),
    .Y(_13226_));
 AO32x1_ASAP7_75t_R _33552_ (.A1(_12807_),
    .A2(_12947_),
    .A3(_12904_),
    .B1(_12952_),
    .B2(_13226_),
    .Y(_13227_));
 AO22x1_ASAP7_75t_R _33553_ (.A1(_12845_),
    .A2(_13226_),
    .B1(_13227_),
    .B2(_12927_),
    .Y(_13228_));
 AND3x2_ASAP7_75t_R _33554_ (.A(_12787_),
    .B(_12912_),
    .C(_12956_),
    .Y(_13229_));
 OA21x2_ASAP7_75t_R _33555_ (.A1(_13044_),
    .A2(_13229_),
    .B(_12771_),
    .Y(_13230_));
 AO21x1_ASAP7_75t_R _33556_ (.A1(_12771_),
    .A2(_13054_),
    .B(_13024_),
    .Y(_13231_));
 OA211x2_ASAP7_75t_R _33557_ (.A1(_12807_),
    .A2(_12947_),
    .B(_12919_),
    .C(_13231_),
    .Y(_13232_));
 AO21x1_ASAP7_75t_R _33558_ (.A1(_12951_),
    .A2(_13226_),
    .B(_13232_),
    .Y(_13233_));
 OR3x1_ASAP7_75t_R _33559_ (.A(_13179_),
    .B(_13230_),
    .C(_13233_),
    .Y(_13234_));
 OR3x1_ASAP7_75t_R _33560_ (.A(_12771_),
    .B(_12823_),
    .C(_12938_),
    .Y(_13235_));
 OA211x2_ASAP7_75t_R _33561_ (.A1(_12947_),
    .A2(_13226_),
    .B(_13235_),
    .C(_12932_),
    .Y(_13236_));
 AO21x1_ASAP7_75t_R _33562_ (.A1(_12915_),
    .A2(_13234_),
    .B(_13236_),
    .Y(_13237_));
 OA21x2_ASAP7_75t_R _33563_ (.A1(_12771_),
    .A2(_12930_),
    .B(_13237_),
    .Y(_13238_));
 OR3x1_ASAP7_75t_R _33564_ (.A(_09319_),
    .B(_13228_),
    .C(_13238_),
    .Y(_13239_));
 OA21x2_ASAP7_75t_R _33565_ (.A1(_13355_),
    .A2(_06686_),
    .B(_13239_),
    .Y(_04495_));
 OA21x2_ASAP7_75t_R _33566_ (.A1(_12814_),
    .A2(_12930_),
    .B(_12915_),
    .Y(_13240_));
 OA21x2_ASAP7_75t_R _33567_ (.A1(_12978_),
    .A2(_13229_),
    .B(_12742_),
    .Y(_13241_));
 AND2x2_ASAP7_75t_R _33568_ (.A(_12593_),
    .B(_00239_),
    .Y(_13242_));
 AO21x1_ASAP7_75t_R _33569_ (.A1(_06734_),
    .A2(_01804_),
    .B(_13242_),
    .Y(_13243_));
 NAND2x1_ASAP7_75t_R _33570_ (.A(_00240_),
    .B(net2648),
    .Y(_13244_));
 OR2x2_ASAP7_75t_R _33571_ (.A(_00240_),
    .B(_01821_),
    .Y(_13245_));
 AO21x1_ASAP7_75t_R _33572_ (.A1(_13244_),
    .A2(_13245_),
    .B(_06580_),
    .Y(_13246_));
 OA21x2_ASAP7_75t_R _33573_ (.A1(_00662_),
    .A2(_13243_),
    .B(_13246_),
    .Y(_13247_));
 INVx1_ASAP7_75t_R _33574_ (.A(_13247_),
    .Y(_13248_));
 AND3x2_ASAP7_75t_R _33575_ (.A(_12807_),
    .B(_12814_),
    .C(_12948_),
    .Y(_13249_));
 OA21x2_ASAP7_75t_R _33576_ (.A1(_12906_),
    .A2(_13248_),
    .B(_13249_),
    .Y(_13250_));
 OA21x2_ASAP7_75t_R _33577_ (.A1(_12992_),
    .A2(_13163_),
    .B(_12814_),
    .Y(_13251_));
 OR4x1_ASAP7_75t_R _33578_ (.A(_12980_),
    .B(_13241_),
    .C(_13250_),
    .D(_13251_),
    .Y(_13252_));
 AND2x2_ASAP7_75t_R _33579_ (.A(_12952_),
    .B(_13248_),
    .Y(_13253_));
 AO21x1_ASAP7_75t_R _33580_ (.A1(_12814_),
    .A2(_12922_),
    .B(_13253_),
    .Y(_13254_));
 AND3x1_ASAP7_75t_R _33581_ (.A(_12814_),
    .B(_12947_),
    .C(_12832_),
    .Y(_13255_));
 AO32x1_ASAP7_75t_R _33582_ (.A1(_12733_),
    .A2(_12966_),
    .A3(_13248_),
    .B1(_13255_),
    .B2(_12932_),
    .Y(_13256_));
 AO221x1_ASAP7_75t_R _33583_ (.A1(_13240_),
    .A2(_13252_),
    .B1(_13254_),
    .B2(_12927_),
    .C(_13256_),
    .Y(_13257_));
 AO21x1_ASAP7_75t_R _33584_ (.A1(_06618_),
    .A2(_06685_),
    .B(_13528_),
    .Y(_13258_));
 OA21x2_ASAP7_75t_R _33585_ (.A1(net254),
    .A2(_13257_),
    .B(_13258_),
    .Y(_04496_));
 OR3x1_ASAP7_75t_R _33586_ (.A(_12780_),
    .B(_12832_),
    .C(_12840_),
    .Y(_13259_));
 OA211x2_ASAP7_75t_R _33587_ (.A1(_12764_),
    .A2(_12919_),
    .B(_13259_),
    .C(_12914_),
    .Y(_13260_));
 AND2x2_ASAP7_75t_R _33588_ (.A(net428),
    .B(net2662),
    .Y(_13261_));
 AO21x1_ASAP7_75t_R _33589_ (.A1(_06589_),
    .A2(_12540_),
    .B(_13261_),
    .Y(_13262_));
 NAND2x1_ASAP7_75t_R _33590_ (.A(_06734_),
    .B(_01803_),
    .Y(_13263_));
 OA211x2_ASAP7_75t_R _33591_ (.A1(net2658),
    .A2(_06734_),
    .B(_13263_),
    .C(_06580_),
    .Y(_13264_));
 AO21x1_ASAP7_75t_R _33592_ (.A1(net430),
    .A2(_13262_),
    .B(_13264_),
    .Y(_13265_));
 AO21x1_ASAP7_75t_R _33593_ (.A1(_12914_),
    .A2(_12922_),
    .B(_13265_),
    .Y(_13266_));
 OA211x2_ASAP7_75t_R _33594_ (.A1(_12966_),
    .A2(_13260_),
    .B(_13266_),
    .C(_13001_),
    .Y(_13267_));
 OA21x2_ASAP7_75t_R _33595_ (.A1(_12906_),
    .A2(_13265_),
    .B(_13249_),
    .Y(_13268_));
 AO21x1_ASAP7_75t_R _33596_ (.A1(_12780_),
    .A2(_12958_),
    .B(_13268_),
    .Y(_13269_));
 OA21x2_ASAP7_75t_R _33597_ (.A1(_12977_),
    .A2(_13229_),
    .B(_12764_),
    .Y(_13270_));
 OA21x2_ASAP7_75t_R _33598_ (.A1(_13269_),
    .A2(_13270_),
    .B(_13219_),
    .Y(_13271_));
 AND2x2_ASAP7_75t_R _33599_ (.A(_12742_),
    .B(_12904_),
    .Y(_13272_));
 AO21x1_ASAP7_75t_R _33600_ (.A1(_12780_),
    .A2(_12840_),
    .B(_13272_),
    .Y(_13273_));
 AND3x1_ASAP7_75t_R _33601_ (.A(_12932_),
    .B(_13078_),
    .C(_13273_),
    .Y(_13274_));
 OA211x2_ASAP7_75t_R _33602_ (.A1(_12992_),
    .A2(_13044_),
    .B(_12814_),
    .C(_12915_),
    .Y(_13275_));
 OR5x2_ASAP7_75t_R _33603_ (.A(_09319_),
    .B(_13267_),
    .C(_13271_),
    .D(_13274_),
    .E(_13275_),
    .Y(_13276_));
 OA21x2_ASAP7_75t_R _33604_ (.A1(_14362_),
    .A2(_06686_),
    .B(_13276_),
    .Y(_04497_));
 AND2x2_ASAP7_75t_R _33605_ (.A(net428),
    .B(net2595),
    .Y(_13277_));
 AO21x1_ASAP7_75t_R _33606_ (.A1(_06589_),
    .A2(_12542_),
    .B(_13277_),
    .Y(_13278_));
 NAND2x1_ASAP7_75t_R _33607_ (.A(_06734_),
    .B(_01802_),
    .Y(_13279_));
 OA211x2_ASAP7_75t_R _33608_ (.A1(net2584),
    .A2(_06734_),
    .B(_13279_),
    .C(_06580_),
    .Y(_13280_));
 AO21x2_ASAP7_75t_R _33609_ (.A1(net430),
    .A2(_13278_),
    .B(_13280_),
    .Y(_13281_));
 AO221x1_ASAP7_75t_R _33610_ (.A1(_12787_),
    .A2(_12980_),
    .B1(_13281_),
    .B2(_12952_),
    .C(_12928_),
    .Y(_13282_));
 OA21x2_ASAP7_75t_R _33611_ (.A1(_12906_),
    .A2(_13281_),
    .B(_13249_),
    .Y(_13283_));
 AO221x1_ASAP7_75t_R _33612_ (.A1(_12771_),
    .A2(_12978_),
    .B1(_13229_),
    .B2(_12750_),
    .C(_13283_),
    .Y(_13284_));
 AND2x2_ASAP7_75t_R _33613_ (.A(_12750_),
    .B(_12904_),
    .Y(_13285_));
 AO21x1_ASAP7_75t_R _33614_ (.A1(_12787_),
    .A2(_12840_),
    .B(_13285_),
    .Y(_13286_));
 AO221x1_ASAP7_75t_R _33615_ (.A1(_12823_),
    .A2(_13281_),
    .B1(_13286_),
    .B2(_13078_),
    .C(_12914_),
    .Y(_13287_));
 AO221x1_ASAP7_75t_R _33616_ (.A1(_12845_),
    .A2(_13281_),
    .B1(_13287_),
    .B2(_12926_),
    .C(_13275_),
    .Y(_13288_));
 AO21x1_ASAP7_75t_R _33617_ (.A1(_13219_),
    .A2(_13284_),
    .B(_13288_),
    .Y(_13289_));
 AND3x1_ASAP7_75t_R _33618_ (.A(_06686_),
    .B(_13282_),
    .C(_13289_),
    .Y(_13290_));
 AO21x1_ASAP7_75t_R _33619_ (.A1(_14423_),
    .A2(net254),
    .B(_13290_),
    .Y(_04498_));
 AND2x2_ASAP7_75t_R _33620_ (.A(net428),
    .B(net2524),
    .Y(_13291_));
 AO21x1_ASAP7_75t_R _33621_ (.A1(_06589_),
    .A2(_12544_),
    .B(_13291_),
    .Y(_13292_));
 NAND2x1_ASAP7_75t_R _33622_ (.A(_06734_),
    .B(_01801_),
    .Y(_13293_));
 OA211x2_ASAP7_75t_R _33623_ (.A1(net2541),
    .A2(_06734_),
    .B(_13293_),
    .C(_06580_),
    .Y(_13294_));
 AO21x1_ASAP7_75t_R _33624_ (.A1(net430),
    .A2(_13292_),
    .B(_13294_),
    .Y(_13295_));
 AO32x1_ASAP7_75t_R _33625_ (.A1(_12794_),
    .A2(_12927_),
    .A3(_12980_),
    .B1(_12967_),
    .B2(_13295_),
    .Y(_13296_));
 AO21x1_ASAP7_75t_R _33626_ (.A1(_12794_),
    .A2(_12823_),
    .B(_13044_),
    .Y(_13297_));
 OA21x2_ASAP7_75t_R _33627_ (.A1(_12906_),
    .A2(_13295_),
    .B(_13249_),
    .Y(_13298_));
 AO21x1_ASAP7_75t_R _33628_ (.A1(_12757_),
    .A2(_13229_),
    .B(_13298_),
    .Y(_13299_));
 AO221x1_ASAP7_75t_R _33629_ (.A1(_12814_),
    .A2(_12977_),
    .B1(_13297_),
    .B2(_12919_),
    .C(_13299_),
    .Y(_13300_));
 OA21x2_ASAP7_75t_R _33630_ (.A1(_13251_),
    .A2(_13300_),
    .B(_13240_),
    .Y(_13301_));
 OR3x2_ASAP7_75t_R _33631_ (.A(_09319_),
    .B(_13296_),
    .C(_13301_),
    .Y(_13302_));
 OA21x2_ASAP7_75t_R _33632_ (.A1(_14801_),
    .A2(_06686_),
    .B(_13302_),
    .Y(_04499_));
 AND2x2_ASAP7_75t_R _33633_ (.A(net428),
    .B(net2637),
    .Y(_13303_));
 AO21x1_ASAP7_75t_R _33634_ (.A1(_06589_),
    .A2(_12546_),
    .B(_13303_),
    .Y(_13304_));
 NAND2x1_ASAP7_75t_R _33635_ (.A(_06734_),
    .B(_01800_),
    .Y(_13305_));
 OA211x2_ASAP7_75t_R _33636_ (.A1(net2633),
    .A2(_06734_),
    .B(_13305_),
    .C(_06580_),
    .Y(_13306_));
 AOI21x1_ASAP7_75t_R _33637_ (.A1(net430),
    .A2(_13304_),
    .B(_13306_),
    .Y(_13307_));
 NAND2x1_ASAP7_75t_R _33638_ (.A(_12800_),
    .B(_13307_),
    .Y(_13308_));
 AO21x1_ASAP7_75t_R _33639_ (.A1(_12814_),
    .A2(_12832_),
    .B(_12980_),
    .Y(_13309_));
 AO221x1_ASAP7_75t_R _33640_ (.A1(_12800_),
    .A2(_12958_),
    .B1(_13249_),
    .B2(_13308_),
    .C(_13309_),
    .Y(_13310_));
 INVx1_ASAP7_75t_R _33641_ (.A(_13307_),
    .Y(_13311_));
 AO32x1_ASAP7_75t_R _33642_ (.A1(_12800_),
    .A2(_12927_),
    .A3(_12980_),
    .B1(_12967_),
    .B2(_13311_),
    .Y(_13312_));
 AO21x1_ASAP7_75t_R _33643_ (.A1(_13240_),
    .A2(_13310_),
    .B(_13312_),
    .Y(_13313_));
 OR2x2_ASAP7_75t_R _33644_ (.A(net254),
    .B(_13313_),
    .Y(_13314_));
 OA21x2_ASAP7_75t_R _33645_ (.A1(_14546_),
    .A2(_06686_),
    .B(_13314_),
    .Y(_04500_));
 AND2x2_ASAP7_75t_R _33646_ (.A(net428),
    .B(net2548),
    .Y(_13315_));
 AO21x1_ASAP7_75t_R _33647_ (.A1(_06589_),
    .A2(_12548_),
    .B(_13315_),
    .Y(_13316_));
 NAND2x1_ASAP7_75t_R _33648_ (.A(_06734_),
    .B(_01799_),
    .Y(_13317_));
 OA211x2_ASAP7_75t_R _33649_ (.A1(net2558),
    .A2(_06734_),
    .B(_13317_),
    .C(_06580_),
    .Y(_13318_));
 AOI21x1_ASAP7_75t_R _33650_ (.A1(net430),
    .A2(_13316_),
    .B(_13318_),
    .Y(_13319_));
 INVx1_ASAP7_75t_R _33651_ (.A(_13319_),
    .Y(_13320_));
 AO21x1_ASAP7_75t_R _33652_ (.A1(_12800_),
    .A2(_13320_),
    .B(_12907_),
    .Y(_13321_));
 AOI21x1_ASAP7_75t_R _33653_ (.A1(_12807_),
    .A2(_13103_),
    .B(_12906_),
    .Y(_13322_));
 AO21x1_ASAP7_75t_R _33654_ (.A1(_12814_),
    .A2(_13321_),
    .B(_13322_),
    .Y(_13323_));
 AO221x1_ASAP7_75t_R _33655_ (.A1(_12787_),
    .A2(_12958_),
    .B1(_13323_),
    .B2(_12948_),
    .C(_13309_),
    .Y(_13324_));
 AO221x2_ASAP7_75t_R _33656_ (.A1(_12967_),
    .A2(_13320_),
    .B1(_13324_),
    .B2(_13240_),
    .C(_09319_),
    .Y(_13325_));
 OA21x2_ASAP7_75t_R _33657_ (.A1(_13595_),
    .A2(_06686_),
    .B(_13325_),
    .Y(_04501_));
 NAND2x1_ASAP7_75t_R _33658_ (.A(_06734_),
    .B(_01798_),
    .Y(_13326_));
 OA211x2_ASAP7_75t_R _33659_ (.A1(net2505),
    .A2(_06734_),
    .B(_13326_),
    .C(_06580_),
    .Y(_13327_));
 NAND2x1_ASAP7_75t_R _33660_ (.A(_06589_),
    .B(_01738_),
    .Y(_13328_));
 OA211x2_ASAP7_75t_R _33661_ (.A1(_06589_),
    .A2(net2537),
    .B(net430),
    .C(_13328_),
    .Y(_13329_));
 NOR2x1_ASAP7_75t_R _33662_ (.A(_13327_),
    .B(_13329_),
    .Y(_13330_));
 INVx1_ASAP7_75t_R _33663_ (.A(_13330_),
    .Y(_13331_));
 OA21x2_ASAP7_75t_R _33664_ (.A1(_12906_),
    .A2(_13331_),
    .B(_13249_),
    .Y(_13332_));
 OR3x1_ASAP7_75t_R _33665_ (.A(_13061_),
    .B(_13309_),
    .C(_13332_),
    .Y(_13333_));
 AO221x1_ASAP7_75t_R _33666_ (.A1(_12967_),
    .A2(_13331_),
    .B1(_13333_),
    .B2(_13240_),
    .C(_09319_),
    .Y(_13334_));
 OA21x2_ASAP7_75t_R _33667_ (.A1(_14704_),
    .A2(_06686_),
    .B(_13334_),
    .Y(_04502_));
 INVx1_ASAP7_75t_R _33668_ (.A(_18089_),
    .Y(_17297_));
 INVx1_ASAP7_75t_R _33669_ (.A(_17981_),
    .Y(_17038_));
 INVx1_ASAP7_75t_R _33670_ (.A(_18005_),
    .Y(_17053_));
 INVx1_ASAP7_75t_R _33671_ (.A(_17985_),
    .Y(_17054_));
 INVx1_ASAP7_75t_R _33672_ (.A(_18004_),
    .Y(_17040_));
 INVx1_ASAP7_75t_R _33673_ (.A(_18023_),
    .Y(_17100_));
 INVx1_ASAP7_75t_R _33674_ (.A(_18003_),
    .Y(_17101_));
 INVx1_ASAP7_75t_R _33675_ (.A(_18001_),
    .Y(_17047_));
 INVx1_ASAP7_75t_R _33676_ (.A(_17984_),
    .Y(_17048_));
 INVx1_ASAP7_75t_R _33677_ (.A(_17982_),
    .Y(_16997_));
 INVx1_ASAP7_75t_R _33678_ (.A(_18000_),
    .Y(_17037_));
 INVx1_ASAP7_75t_R _33679_ (.A(_18048_),
    .Y(_17217_));
 INVx1_ASAP7_75t_R _33680_ (.A(_18076_),
    .Y(_17216_));
 INVx1_ASAP7_75t_R _33681_ (.A(_17948_),
    .Y(_16965_));
 INVx1_ASAP7_75t_R _33682_ (.A(_17966_),
    .Y(_16964_));
 INVx1_ASAP7_75t_R _33683_ (.A(_18038_),
    .Y(_17194_));
 INVx1_ASAP7_75t_R _33684_ (.A(_18070_),
    .Y(_17193_));
 INVx1_ASAP7_75t_R _33685_ (.A(_18039_),
    .Y(_17197_));
 INVx1_ASAP7_75t_R _33686_ (.A(_18066_),
    .Y(_17196_));
 INVx1_ASAP7_75t_R _33687_ (.A(_01362_),
    .Y(_17842_));
 INVx1_ASAP7_75t_R _33688_ (.A(_18043_),
    .Y(_17208_));
 INVx1_ASAP7_75t_R _33689_ (.A(_18072_),
    .Y(_17207_));
 INVx1_ASAP7_75t_R _33690_ (.A(_18022_),
    .Y(_17151_));
 INVx1_ASAP7_75t_R _33691_ (.A(_18044_),
    .Y(_17150_));
 INVx1_ASAP7_75t_R _33692_ (.A(_17949_),
    .Y(_16932_));
 INVx1_ASAP7_75t_R _33693_ (.A(_18045_),
    .Y(_17209_));
 INVx1_ASAP7_75t_R _33694_ (.A(_18046_),
    .Y(_17212_));
 INVx1_ASAP7_75t_R _33695_ (.A(_18075_),
    .Y(_17211_));
 INVx1_ASAP7_75t_R _33696_ (.A(_18006_),
    .Y(_17102_));
 INVx1_ASAP7_75t_R _33697_ (.A(_17999_),
    .Y(_17033_));
 INVx1_ASAP7_75t_R _33698_ (.A(_01367_),
    .Y(_17852_));
 INVx1_ASAP7_75t_R _33699_ (.A(_18218_),
    .Y(_17507_));
 INVx1_ASAP7_75t_R _33700_ (.A(_18200_),
    .Y(_17508_));
 INVx1_ASAP7_75t_R _33701_ (.A(_18195_),
    .Y(_17459_));
 INVx1_ASAP7_75t_R _33702_ (.A(_01428_),
    .Y(_17915_));
 INVx1_ASAP7_75t_R _33703_ (.A(_00010_),
    .Y(_17962_));
 INVx1_ASAP7_75t_R _33704_ (.A(_17986_),
    .Y(_17011_));
 INVx1_ASAP7_75t_R _33705_ (.A(_17968_),
    .Y(_17012_));
 INVx1_ASAP7_75t_R _33706_ (.A(_00066_),
    .Y(_17724_));
 INVx1_ASAP7_75t_R _33707_ (.A(_18174_),
    .Y(_17460_));
 INVx1_ASAP7_75t_R _33708_ (.A(_18160_),
    .Y(_17380_));
 INVx1_ASAP7_75t_R _33709_ (.A(_18135_),
    .Y(_17381_));
 INVx1_ASAP7_75t_R _33710_ (.A(_02297_),
    .Y(_17836_));
 INVx1_ASAP7_75t_R _33711_ (.A(_02298_),
    .Y(_17838_));
 INVx1_ASAP7_75t_R _33712_ (.A(_01361_),
    .Y(_17839_));
 INVx1_ASAP7_75t_R _33713_ (.A(_18157_),
    .Y(_17375_));
 INVx1_ASAP7_75t_R _33714_ (.A(_18133_),
    .Y(_17376_));
 INVx1_ASAP7_75t_R _33715_ (.A(_01435_),
    .Y(_16941_));
 INVx1_ASAP7_75t_R _33716_ (.A(_18027_),
    .Y(_17162_));
 INVx1_ASAP7_75t_R _33717_ (.A(_18049_),
    .Y(_17161_));
 INVx1_ASAP7_75t_R _33718_ (.A(_18024_),
    .Y(_17153_));
 INVx1_ASAP7_75t_R _33719_ (.A(_18052_),
    .Y(_17152_));
 INVx1_ASAP7_75t_R _33720_ (.A(_18025_),
    .Y(_17157_));
 INVx1_ASAP7_75t_R _33721_ (.A(_18047_),
    .Y(_17156_));
 INVx1_ASAP7_75t_R _33722_ (.A(_18029_),
    .Y(_17172_));
 INVx1_ASAP7_75t_R _33723_ (.A(_18055_),
    .Y(_17171_));
 INVx1_ASAP7_75t_R _33724_ (.A(net2233),
    .Y(_17174_));
 INVx1_ASAP7_75t_R _33725_ (.A(_18053_),
    .Y(_17222_));
 INVx1_ASAP7_75t_R _33726_ (.A(_18081_),
    .Y(_17221_));
 INVx1_ASAP7_75t_R _33727_ (.A(_18054_),
    .Y(_17224_));
 INVx1_ASAP7_75t_R _33728_ (.A(_18080_),
    .Y(_17223_));
 INVx1_ASAP7_75t_R _33729_ (.A(_02340_),
    .Y(_17139_));
 INVx1_ASAP7_75t_R _33730_ (.A(_00022_),
    .Y(_17088_));
 INVx1_ASAP7_75t_R _33731_ (.A(_00021_),
    .Y(_17081_));
 INVx1_ASAP7_75t_R _33732_ (.A(_17939_),
    .Y(_16918_));
 INVx1_ASAP7_75t_R _33733_ (.A(_18199_),
    .Y(_17464_));
 INVx1_ASAP7_75t_R _33734_ (.A(_18176_),
    .Y(_17465_));
 INVx1_ASAP7_75t_R _33735_ (.A(_01363_),
    .Y(_17843_));
 INVx1_ASAP7_75t_R _33736_ (.A(_02296_),
    .Y(_17834_));
 INVx1_ASAP7_75t_R _33737_ (.A(_01359_),
    .Y(_17835_));
 INVx1_ASAP7_75t_R _33738_ (.A(_18161_),
    .Y(_17431_));
 INVx1_ASAP7_75t_R _33739_ (.A(_18185_),
    .Y(_17430_));
 INVx1_ASAP7_75t_R _33740_ (.A(_02295_),
    .Y(_17831_));
 INVx1_ASAP7_75t_R _33741_ (.A(_01358_),
    .Y(_17832_));
 INVx1_ASAP7_75t_R _33742_ (.A(_18201_),
    .Y(_17471_));
 INVx1_ASAP7_75t_R _33743_ (.A(_18180_),
    .Y(_17472_));
 INVx1_ASAP7_75t_R _33744_ (.A(_18179_),
    .Y(_17421_));
 INVx1_ASAP7_75t_R _33745_ (.A(_18155_),
    .Y(_17422_));
 INVx1_ASAP7_75t_R _33746_ (.A(_02333_),
    .Y(_17024_));
 INVx1_ASAP7_75t_R _33747_ (.A(_18131_),
    .Y(_17324_));
 INVx1_ASAP7_75t_R _33748_ (.A(_18107_),
    .Y(_17325_));
 INVx1_ASAP7_75t_R _33749_ (.A(_02351_),
    .Y(_17487_));
 INVx1_ASAP7_75t_R _33750_ (.A(_00048_),
    .Y(_17447_));
 INVx1_ASAP7_75t_R _33751_ (.A(_18132_),
    .Y(_17374_));
 INVx1_ASAP7_75t_R _33752_ (.A(_18158_),
    .Y(_17373_));
 INVx1_ASAP7_75t_R _33753_ (.A(_18154_),
    .Y(_17368_));
 INVx1_ASAP7_75t_R _33754_ (.A(_18130_),
    .Y(_17369_));
 INVx1_ASAP7_75t_R _33755_ (.A(_01365_),
    .Y(_17846_));
 INVx1_ASAP7_75t_R _33756_ (.A(_02300_),
    .Y(_16778_));
 INVx1_ASAP7_75t_R _33757_ (.A(_17557_),
    .Y(_17516_));
 INVx2_ASAP7_75t_R _33758_ (.A(_17519_),
    .Y(_17517_));
 INVx1_ASAP7_75t_R _33759_ (.A(_02294_),
    .Y(_17828_));
 INVx1_ASAP7_75t_R _33760_ (.A(_18175_),
    .Y(_17416_));
 INVx1_ASAP7_75t_R _33761_ (.A(_18153_),
    .Y(_17417_));
 INVx1_ASAP7_75t_R _33762_ (.A(_18215_),
    .Y(_17502_));
 INVx1_ASAP7_75t_R _33763_ (.A(_18197_),
    .Y(_17503_));
 INVx1_ASAP7_75t_R _33764_ (.A(_18216_),
    .Y(_17500_));
 INVx1_ASAP7_75t_R _33765_ (.A(_18196_),
    .Y(_17501_));
 INVx1_ASAP7_75t_R _33766_ (.A(_18212_),
    .Y(_17495_));
 INVx1_ASAP7_75t_R _33767_ (.A(_18194_),
    .Y(_17496_));
 INVx1_ASAP7_75t_R _33768_ (.A(_02308_),
    .Y(_16802_));
 INVx1_ASAP7_75t_R _33769_ (.A(_01373_),
    .Y(_16779_));
 INVx1_ASAP7_75t_R _33770_ (.A(_02302_),
    .Y(_17851_));
 INVx1_ASAP7_75t_R _33771_ (.A(_18042_),
    .Y(_17138_));
 INVx1_ASAP7_75t_R _33772_ (.A(_18085_),
    .Y(_17235_));
 INVx1_ASAP7_75t_R _33773_ (.A(_01400_),
    .Y(_16827_));
 INVx1_ASAP7_75t_R _33774_ (.A(_17994_),
    .Y(_17028_));
 INVx1_ASAP7_75t_R _33775_ (.A(_17975_),
    .Y(_17029_));
 INVx1_ASAP7_75t_R _33776_ (.A(_02332_),
    .Y(_17014_));
 INVx1_ASAP7_75t_R _33777_ (.A(_01440_),
    .Y(_16973_));
 INVx1_ASAP7_75t_R _33778_ (.A(_02331_),
    .Y(_17000_));
 INVx1_ASAP7_75t_R _33779_ (.A(_18060_),
    .Y(_17236_));
 INVx1_ASAP7_75t_R _33780_ (.A(_18007_),
    .Y(_17059_));
 INVx1_ASAP7_75t_R _33781_ (.A(_02311_),
    .Y(_17870_));
 INVx1_ASAP7_75t_R _33782_ (.A(_01380_),
    .Y(_17871_));
 INVx1_ASAP7_75t_R _33783_ (.A(_02304_),
    .Y(_16792_));
 INVx1_ASAP7_75t_R _33784_ (.A(_18173_),
    .Y(_17410_));
 INVx1_ASAP7_75t_R _33785_ (.A(_18149_),
    .Y(_17411_));
 INVx1_ASAP7_75t_R _33786_ (.A(_18014_),
    .Y(_17118_));
 INVx1_ASAP7_75t_R _33787_ (.A(_18030_),
    .Y(_17117_));
 INVx1_ASAP7_75t_R _33788_ (.A(_18019_),
    .Y(_17145_));
 INVx1_ASAP7_75t_R _33789_ (.A(_18041_),
    .Y(_17144_));
 INVx1_ASAP7_75t_R _33790_ (.A(_16783_),
    .Y(_17855_));
 INVx1_ASAP7_75t_R _33791_ (.A(_01414_),
    .Y(_17893_));
 INVx1_ASAP7_75t_R _33792_ (.A(_02319_),
    .Y(_17884_));
 INVx1_ASAP7_75t_R _33793_ (.A(_01401_),
    .Y(_17885_));
 INVx1_ASAP7_75t_R _33794_ (.A(_18010_),
    .Y(_17064_));
 INVx1_ASAP7_75t_R _33795_ (.A(_02321_),
    .Y(_16868_));
 INVx1_ASAP7_75t_R _33796_ (.A(_01405_),
    .Y(_16836_));
 INVx1_ASAP7_75t_R _33797_ (.A(_02316_),
    .Y(_17879_));
 INVx1_ASAP7_75t_R _33798_ (.A(_01392_),
    .Y(_17880_));
 INVx1_ASAP7_75t_R _33799_ (.A(_02306_),
    .Y(_17862_));
 INVx1_ASAP7_75t_R _33800_ (.A(_01371_),
    .Y(_17863_));
 INVx1_ASAP7_75t_R _33801_ (.A(_00242_),
    .Y(_17753_));
 INVx1_ASAP7_75t_R _33802_ (.A(_17740_),
    .Y(_17739_));
 INVx1_ASAP7_75t_R _33803_ (.A(_18059_),
    .Y(_17179_));
 INVx1_ASAP7_75t_R _33804_ (.A(_02345_),
    .Y(_17316_));
 INVx1_ASAP7_75t_R _33805_ (.A(_00035_),
    .Y(_17269_));
 INVx1_ASAP7_75t_R _33806_ (.A(_18033_),
    .Y(_17180_));
 INVx1_ASAP7_75t_R _33807_ (.A(_18017_),
    .Y(_17136_));
 INVx1_ASAP7_75t_R _33808_ (.A(_18037_),
    .Y(_17135_));
 INVx1_ASAP7_75t_R _33809_ (.A(_02299_),
    .Y(_17841_));
 INVx1_ASAP7_75t_R _33810_ (.A(_18147_),
    .Y(_17353_));
 INVx1_ASAP7_75t_R _33811_ (.A(_01430_),
    .Y(_16907_));
 INVx1_ASAP7_75t_R _33812_ (.A(_18123_),
    .Y(_17354_));
 INVx1_ASAP7_75t_R _33813_ (.A(_01369_),
    .Y(_17858_));
 INVx1_ASAP7_75t_R _33814_ (.A(_18115_),
    .Y(_17296_));
 INVx1_ASAP7_75t_R _33815_ (.A(_18275_),
    .Y(_17647_));
 INVx1_ASAP7_75t_R _33816_ (.A(_18122_),
    .Y(_17352_));
 INVx1_ASAP7_75t_R _33817_ (.A(_17889_),
    .Y(_16812_));
 INVx1_ASAP7_75t_R _33818_ (.A(_17876_),
    .Y(_16813_));
 INVx1_ASAP7_75t_R _33819_ (.A(_17896_),
    .Y(_16831_));
 INVx1_ASAP7_75t_R _33820_ (.A(_17888_),
    .Y(_16832_));
 INVx1_ASAP7_75t_R _33821_ (.A(_18223_),
    .Y(_17560_));
 INVx1_ASAP7_75t_R _33822_ (.A(_18125_),
    .Y(_17306_));
 INVx1_ASAP7_75t_R _33823_ (.A(_18002_),
    .Y(_17095_));
 INVx1_ASAP7_75t_R _33824_ (.A(_02325_),
    .Y(_16919_));
 INVx1_ASAP7_75t_R _33825_ (.A(_01424_),
    .Y(_16891_));
 INVx1_ASAP7_75t_R _33826_ (.A(_17958_),
    .Y(_16955_));
 INVx1_ASAP7_75t_R _33827_ (.A(_17938_),
    .Y(_16956_));
 INVx1_ASAP7_75t_R _33828_ (.A(_01381_),
    .Y(_16799_));
 INVx1_ASAP7_75t_R _33829_ (.A(_02312_),
    .Y(_16820_));
 INVx1_ASAP7_75t_R _33830_ (.A(_18172_),
    .Y(_17451_));
 INVx1_ASAP7_75t_R _33831_ (.A(_18191_),
    .Y(_17450_));
 INVx1_ASAP7_75t_R _33832_ (.A(_18093_),
    .Y(_17307_));
 INVx1_ASAP7_75t_R _33833_ (.A(_17959_),
    .Y(_16951_));
 INVx1_ASAP7_75t_R _33834_ (.A(_17937_),
    .Y(_16952_));
 INVx1_ASAP7_75t_R _33835_ (.A(_17974_),
    .Y(_16989_));
 INVx1_ASAP7_75t_R _33836_ (.A(_17957_),
    .Y(_16990_));
 INVx1_ASAP7_75t_R _33837_ (.A(_18298_),
    .Y(_17666_));
 INVx1_ASAP7_75t_R _33838_ (.A(_17976_),
    .Y(_16985_));
 INVx1_ASAP7_75t_R _33839_ (.A(_17956_),
    .Y(_16986_));
 INVx1_ASAP7_75t_R _33840_ (.A(_17720_),
    .Y(_17717_));
 INVx1_ASAP7_75t_R _33841_ (.A(_17742_),
    .Y(_17716_));
 INVx1_ASAP7_75t_R _33842_ (.A(_18034_),
    .Y(_17124_));
 INVx1_ASAP7_75t_R _33843_ (.A(_18035_),
    .Y(_17186_));
 INVx1_ASAP7_75t_R _33844_ (.A(_18061_),
    .Y(_17185_));
 INVx1_ASAP7_75t_R _33845_ (.A(_18069_),
    .Y(_17256_));
 INVx1_ASAP7_75t_R _33846_ (.A(_18065_),
    .Y(_17246_));
 INVx1_ASAP7_75t_R _33847_ (.A(_18090_),
    .Y(_17245_));
 INVx1_ASAP7_75t_R _33848_ (.A(_17983_),
    .Y(_17005_));
 INVx1_ASAP7_75t_R _33849_ (.A(_18150_),
    .Y(_17359_));
 INVx1_ASAP7_75t_R _33850_ (.A(_18128_),
    .Y(_17360_));
 INVx1_ASAP7_75t_R _33851_ (.A(_17967_),
    .Y(_17006_));
 INVx1_ASAP7_75t_R _33852_ (.A(_18124_),
    .Y(_17311_));
 INVx1_ASAP7_75t_R _33853_ (.A(_18098_),
    .Y(_17312_));
 INVx1_ASAP7_75t_R _33854_ (.A(_18097_),
    .Y(_17310_));
 INVx1_ASAP7_75t_R _33855_ (.A(_18068_),
    .Y(_17201_));
 INVx1_ASAP7_75t_R _33856_ (.A(_18040_),
    .Y(_17202_));
 INVx1_ASAP7_75t_R _33857_ (.A(_18100_),
    .Y(_17255_));
 INVx1_ASAP7_75t_R _33858_ (.A(_18094_),
    .Y(_17243_));
 INVx1_ASAP7_75t_R _33859_ (.A(_18064_),
    .Y(_17244_));
 INVx1_ASAP7_75t_R _33860_ (.A(_18063_),
    .Y(_17190_));
 INVx2_ASAP7_75t_R _33861_ (.A(_18036_),
    .Y(_17191_));
 INVx1_ASAP7_75t_R _33862_ (.A(_17925_),
    .Y(_16890_));
 INVx1_ASAP7_75t_R _33863_ (.A(_18244_),
    .Y(_17561_));
 INVx1_ASAP7_75t_R _33864_ (.A(_18224_),
    .Y(_17562_));
 INVx1_ASAP7_75t_R _33865_ (.A(_00011_),
    .Y(_16998_));
 INVx1_ASAP7_75t_R _33866_ (.A(_02334_),
    .Y(_17041_));
 INVx1_ASAP7_75t_R _33867_ (.A(_18087_),
    .Y(_17240_));
 INVx1_ASAP7_75t_R _33868_ (.A(_18062_),
    .Y(_17241_));
 INVx1_ASAP7_75t_R _33869_ (.A(_17723_),
    .Y(_17690_));
 INVx1_ASAP7_75t_R _33870_ (.A(_00018_),
    .Y(_17068_));
 INVx1_ASAP7_75t_R _33871_ (.A(_02338_),
    .Y(_17114_));
 INVx1_ASAP7_75t_R _33872_ (.A(_02324_),
    .Y(_16906_));
 INVx1_ASAP7_75t_R _33873_ (.A(_01421_),
    .Y(_17901_));
 INVx1_ASAP7_75t_R _33874_ (.A(_02328_),
    .Y(_16940_));
 INVx1_ASAP7_75t_R _33875_ (.A(_01429_),
    .Y(_16905_));
 INVx1_ASAP7_75t_R _33876_ (.A(_02337_),
    .Y(_17089_));
 INVx1_ASAP7_75t_R _33877_ (.A(_18299_),
    .Y(_17698_));
 INVx1_ASAP7_75t_R _33878_ (.A(_18308_),
    .Y(_17697_));
 INVx1_ASAP7_75t_R _33879_ (.A(_18020_),
    .Y(_17094_));
 INVx1_ASAP7_75t_R _33880_ (.A(_17929_),
    .Y(_16933_));
 INVx1_ASAP7_75t_R _33881_ (.A(_17950_),
    .Y(_16971_));
 INVx1_ASAP7_75t_R _33882_ (.A(_17969_),
    .Y(_16970_));
 INVx1_ASAP7_75t_R _33883_ (.A(_01408_),
    .Y(_16841_));
 INVx2_ASAP7_75t_R _33884_ (.A(_01419_),
    .Y(_16840_));
 INVx1_ASAP7_75t_R _33885_ (.A(_18302_),
    .Y(_17699_));
 INVx1_ASAP7_75t_R _33886_ (.A(_01431_),
    .Y(_16908_));
 INVx1_ASAP7_75t_R _33887_ (.A(_17987_),
    .Y(_17056_));
 INVx1_ASAP7_75t_R _33888_ (.A(_00043_),
    .Y(_17407_));
 INVx1_ASAP7_75t_R _33889_ (.A(_02339_),
    .Y(_17130_));
 INVx1_ASAP7_75t_R _33890_ (.A(_17918_),
    .Y(_16875_));
 INVx1_ASAP7_75t_R _33891_ (.A(_17902_),
    .Y(_16876_));
 INVx1_ASAP7_75t_R _33892_ (.A(_18300_),
    .Y(_17670_));
 INVx1_ASAP7_75t_R _33893_ (.A(_02320_),
    .Y(_16865_));
 INVx1_ASAP7_75t_R _33894_ (.A(_18121_),
    .Y(_17308_));
 INVx1_ASAP7_75t_R _33895_ (.A(_18095_),
    .Y(_17309_));
 INVx1_ASAP7_75t_R _33896_ (.A(_01403_),
    .Y(_16834_));
 INVx1_ASAP7_75t_R _33897_ (.A(_18088_),
    .Y(_17295_));
 INVx1_ASAP7_75t_R _33898_ (.A(_18119_),
    .Y(_17294_));
 INVx1_ASAP7_75t_R _33899_ (.A(_18318_),
    .Y(_17747_));
 INVx1_ASAP7_75t_R _33900_ (.A(_18320_),
    .Y(_17749_));
 INVx1_ASAP7_75t_R _33901_ (.A(_17741_),
    .Y(_17715_));
 INVx1_ASAP7_75t_R _33902_ (.A(_18067_),
    .Y(_17251_));
 INVx1_ASAP7_75t_R _33903_ (.A(_18249_),
    .Y(_17609_));
 INVx1_ASAP7_75t_R _33904_ (.A(_18270_),
    .Y(_17608_));
 INVx1_ASAP7_75t_R _33905_ (.A(_18230_),
    .Y(_17572_));
 INVx1_ASAP7_75t_R _33906_ (.A(_18248_),
    .Y(_17571_));
 INVx1_ASAP7_75t_R _33907_ (.A(_18092_),
    .Y(_17250_));
 INVx1_ASAP7_75t_R _33908_ (.A(_01378_),
    .Y(_16797_));
 INVx1_ASAP7_75t_R _33909_ (.A(_02310_),
    .Y(_16816_));
 INVx1_ASAP7_75t_R _33910_ (.A(_01415_),
    .Y(_16864_));
 INVx1_ASAP7_75t_R _33911_ (.A(_02323_),
    .Y(_16892_));
 INVx1_ASAP7_75t_R _33912_ (.A(_02327_),
    .Y(_17914_));
 INVx1_ASAP7_75t_R _33913_ (.A(_01423_),
    .Y(_17905_));
 INVx1_ASAP7_75t_R _33914_ (.A(_00014_),
    .Y(_17022_));
 INVx1_ASAP7_75t_R _33915_ (.A(_00017_),
    .Y(_17043_));
 INVx1_ASAP7_75t_R _33916_ (.A(_02335_),
    .Y(_17069_));
 INVx1_ASAP7_75t_R _33917_ (.A(_18071_),
    .Y(_17258_));
 INVx1_ASAP7_75t_R _33918_ (.A(_18096_),
    .Y(_17257_));
 INVx1_ASAP7_75t_R _33919_ (.A(_18159_),
    .Y(_17429_));
 INVx1_ASAP7_75t_R _33920_ (.A(_18181_),
    .Y(_17428_));
 INVx1_ASAP7_75t_R _33921_ (.A(_18202_),
    .Y(_17510_));
 INVx1_ASAP7_75t_R _33922_ (.A(_18222_),
    .Y(_17509_));
 INVx1_ASAP7_75t_R _33923_ (.A(_18177_),
    .Y(_17467_));
 INVx1_ASAP7_75t_R _33924_ (.A(_18198_),
    .Y(_17466_));
 INVx1_ASAP7_75t_R _33925_ (.A(_17988_),
    .Y(_17060_));
 INVx1_ASAP7_75t_R _33926_ (.A(_18203_),
    .Y(_17512_));
 INVx1_ASAP7_75t_R _33927_ (.A(_18221_),
    .Y(_17511_));
 INVx1_ASAP7_75t_R _33928_ (.A(_18156_),
    .Y(_17424_));
 INVx1_ASAP7_75t_R _33929_ (.A(_18178_),
    .Y(_17423_));
 INVx1_ASAP7_75t_R _33930_ (.A(_17993_),
    .Y(_17073_));
 INVx1_ASAP7_75t_R _33931_ (.A(_18013_),
    .Y(_17072_));
 INVx1_ASAP7_75t_R _33932_ (.A(_18162_),
    .Y(_17433_));
 INVx1_ASAP7_75t_R _33933_ (.A(_18184_),
    .Y(_17432_));
 INVx1_ASAP7_75t_R _33934_ (.A(_18111_),
    .Y(_17336_));
 INVx1_ASAP7_75t_R _33935_ (.A(_18136_),
    .Y(_17335_));
 INVx1_ASAP7_75t_R _33936_ (.A(_18137_),
    .Y(_17384_));
 INVx1_ASAP7_75t_R _33937_ (.A(_18166_),
    .Y(_17383_));
 INVx1_ASAP7_75t_R _33938_ (.A(_18164_),
    .Y(_17437_));
 INVx1_ASAP7_75t_R _33939_ (.A(_17903_),
    .Y(_16845_));
 INVx1_ASAP7_75t_R _33940_ (.A(_18082_),
    .Y(_17281_));
 INVx1_ASAP7_75t_R _33941_ (.A(_18108_),
    .Y(_17280_));
 INVx1_ASAP7_75t_R _33942_ (.A(_18232_),
    .Y(_17577_));
 INVx1_ASAP7_75t_R _33943_ (.A(_18109_),
    .Y(_17331_));
 INVx1_ASAP7_75t_R _33944_ (.A(_18134_),
    .Y(_17330_));
 INVx1_ASAP7_75t_R _33945_ (.A(_18252_),
    .Y(_17576_));
 INVx1_ASAP7_75t_R _33946_ (.A(_18236_),
    .Y(_17583_));
 INVx1_ASAP7_75t_R _33947_ (.A(_18253_),
    .Y(_17582_));
 INVx1_ASAP7_75t_R _33948_ (.A(_18254_),
    .Y(_17619_));
 INVx1_ASAP7_75t_R _33949_ (.A(_18274_),
    .Y(_17618_));
 INVx1_ASAP7_75t_R _33950_ (.A(_17989_),
    .Y(_17065_));
 INVx1_ASAP7_75t_R _33951_ (.A(_01366_),
    .Y(_17850_));
 INVx1_ASAP7_75t_R _33952_ (.A(_02301_),
    .Y(_17849_));
 INVx1_ASAP7_75t_R _33953_ (.A(_01372_),
    .Y(_17865_));
 INVx1_ASAP7_75t_R _33954_ (.A(_02307_),
    .Y(_17864_));
 INVx1_ASAP7_75t_R _33955_ (.A(_01368_),
    .Y(_17854_));
 INVx1_ASAP7_75t_R _33956_ (.A(_02303_),
    .Y(_17853_));
 INVx1_ASAP7_75t_R _33957_ (.A(_16782_),
    .Y(_17867_));
 INVx1_ASAP7_75t_R _33958_ (.A(_02309_),
    .Y(_17866_));
 INVx1_ASAP7_75t_R _33959_ (.A(_01370_),
    .Y(_16777_));
 INVx1_ASAP7_75t_R _33960_ (.A(_02305_),
    .Y(_16798_));
 INVx2_ASAP7_75t_R _33961_ (.A(_01418_),
    .Y(_16870_));
 INVx1_ASAP7_75t_R _33962_ (.A(_01425_),
    .Y(_16869_));
 INVx1_ASAP7_75t_R _33963_ (.A(_18138_),
    .Y(_17386_));
 INVx1_ASAP7_75t_R _33964_ (.A(_18163_),
    .Y(_17385_));
 INVx1_ASAP7_75t_R _33965_ (.A(_18182_),
    .Y(_17474_));
 INVx1_ASAP7_75t_R _33966_ (.A(_18205_),
    .Y(_17473_));
 INVx1_ASAP7_75t_R _33967_ (.A(_01416_),
    .Y(_16867_));
 INVx1_ASAP7_75t_R _33968_ (.A(_17970_),
    .Y(_17020_));
 INVx1_ASAP7_75t_R _33969_ (.A(_17990_),
    .Y(_17019_));
 INVx1_ASAP7_75t_R _33970_ (.A(_00040_),
    .Y(_17356_));
 INVx1_ASAP7_75t_R _33971_ (.A(_02348_),
    .Y(_17408_));
 INVx1_ASAP7_75t_R _33972_ (.A(_18206_),
    .Y(_17522_));
 INVx1_ASAP7_75t_R _33973_ (.A(_17933_),
    .Y(_16946_));
 INVx1_ASAP7_75t_R _33974_ (.A(_17953_),
    .Y(_16945_));
 INVx1_ASAP7_75t_R _33975_ (.A(_18140_),
    .Y(_17391_));
 INVx1_ASAP7_75t_R _33976_ (.A(_18165_),
    .Y(_17390_));
 INVx1_ASAP7_75t_R _33977_ (.A(_18167_),
    .Y(_17439_));
 INVx1_ASAP7_75t_R _33978_ (.A(_18186_),
    .Y(_17438_));
 INVx1_ASAP7_75t_R _33979_ (.A(_18183_),
    .Y(_17476_));
 INVx1_ASAP7_75t_R _33980_ (.A(_18204_),
    .Y(_17475_));
 INVx1_ASAP7_75t_R _33981_ (.A(_00037_),
    .Y(_17315_));
 INVx1_ASAP7_75t_R _33982_ (.A(_02346_),
    .Y(_17357_));
 INVx1_ASAP7_75t_R _33983_ (.A(_18207_),
    .Y(_17524_));
 INVx1_ASAP7_75t_R _33984_ (.A(_18225_),
    .Y(_17523_));
 INVx1_ASAP7_75t_R _33985_ (.A(_02343_),
    .Y(_17270_));
 INVx1_ASAP7_75t_R _33986_ (.A(_17921_),
    .Y(_16913_));
 INVx1_ASAP7_75t_R _33987_ (.A(_17934_),
    .Y(_16912_));
 INVx1_ASAP7_75t_R _33988_ (.A(_18217_),
    .Y(_17550_));
 INVx1_ASAP7_75t_R _33989_ (.A(_18237_),
    .Y(_17549_));
 INVx1_ASAP7_75t_R _33990_ (.A(_17917_),
    .Y(_16900_));
 INVx1_ASAP7_75t_R _33991_ (.A(_17930_),
    .Y(_16899_));
 INVx1_ASAP7_75t_R _33992_ (.A(_18282_),
    .Y(_17665_));
 INVx1_ASAP7_75t_R _33993_ (.A(_18187_),
    .Y(_17482_));
 INVx1_ASAP7_75t_R _33994_ (.A(_17951_),
    .Y(_16938_));
 INVx1_ASAP7_75t_R _33995_ (.A(_18219_),
    .Y(_17552_));
 INVx1_ASAP7_75t_R _33996_ (.A(_01434_),
    .Y(_16939_));
 INVx1_ASAP7_75t_R _33997_ (.A(_02329_),
    .Y(_16974_));
 INVx1_ASAP7_75t_R _33998_ (.A(_18241_),
    .Y(_17551_));
 INVx1_ASAP7_75t_R _33999_ (.A(_18280_),
    .Y(_17662_));
 INVx1_ASAP7_75t_R _34000_ (.A(_17693_),
    .Y(_17661_));
 INVx1_ASAP7_75t_R _34001_ (.A(_18116_),
    .Y(_17346_));
 INVx1_ASAP7_75t_R _34002_ (.A(_18141_),
    .Y(_17345_));
 INVx1_ASAP7_75t_R _34003_ (.A(_18143_),
    .Y(_17399_));
 INVx1_ASAP7_75t_R _34004_ (.A(_18168_),
    .Y(_17398_));
 INVx1_ASAP7_75t_R _34005_ (.A(_18265_),
    .Y(_17634_));
 INVx1_ASAP7_75t_R _34006_ (.A(_18281_),
    .Y(_17633_));
 INVx1_ASAP7_75t_R _34007_ (.A(_01393_),
    .Y(_16817_));
 INVx1_ASAP7_75t_R _34008_ (.A(_02317_),
    .Y(_16839_));
 INVx1_ASAP7_75t_R _34009_ (.A(_18283_),
    .Y(_17667_));
 INVx1_ASAP7_75t_R _34010_ (.A(_17998_),
    .Y(_17086_));
 INVx1_ASAP7_75t_R _34011_ (.A(_18018_),
    .Y(_17085_));
 INVx1_ASAP7_75t_R _34012_ (.A(_18188_),
    .Y(_17484_));
 INVx1_ASAP7_75t_R _34013_ (.A(_18208_),
    .Y(_17483_));
 INVx1_ASAP7_75t_R _34014_ (.A(_18211_),
    .Y(_17538_));
 INVx1_ASAP7_75t_R _34015_ (.A(_18231_),
    .Y(_17537_));
 INVx1_ASAP7_75t_R _34016_ (.A(_18213_),
    .Y(_17543_));
 INVx1_ASAP7_75t_R _34017_ (.A(_18235_),
    .Y(_17542_));
 INVx1_ASAP7_75t_R _34018_ (.A(_18214_),
    .Y(_17545_));
 INVx1_ASAP7_75t_R _34019_ (.A(_18234_),
    .Y(_17544_));
 INVx1_ASAP7_75t_R _34020_ (.A(_18276_),
    .Y(_17649_));
 INVx1_ASAP7_75t_R _34021_ (.A(_18292_),
    .Y(_17648_));
 INVx1_ASAP7_75t_R _34022_ (.A(_18021_),
    .Y(_17087_));
 INVx1_ASAP7_75t_R _34023_ (.A(_18278_),
    .Y(_17653_));
 INVx1_ASAP7_75t_R _34024_ (.A(_18294_),
    .Y(_17652_));
 INVx1_ASAP7_75t_R _34025_ (.A(_18220_),
    .Y(_17554_));
 INVx1_ASAP7_75t_R _34026_ (.A(_18240_),
    .Y(_17553_));
 INVx1_ASAP7_75t_R _34027_ (.A(_17692_),
    .Y(_17683_));
 INVx1_ASAP7_75t_R _34028_ (.A(_18091_),
    .Y(_17302_));
 INVx1_ASAP7_75t_R _34029_ (.A(_18117_),
    .Y(_17301_));
 INVx1_ASAP7_75t_R _34030_ (.A(_18297_),
    .Y(_17691_));
 INVx1_ASAP7_75t_R _34031_ (.A(_18118_),
    .Y(_17349_));
 INVx1_ASAP7_75t_R _34032_ (.A(_18307_),
    .Y(_17722_));
 INVx1_ASAP7_75t_R _34033_ (.A(_18315_),
    .Y(_17721_));
 INVx1_ASAP7_75t_R _34034_ (.A(_01412_),
    .Y(_16849_));
 INVx1_ASAP7_75t_R _34035_ (.A(_17952_),
    .Y(_16980_));
 INVx1_ASAP7_75t_R _34036_ (.A(_17971_),
    .Y(_16979_));
 INVx1_ASAP7_75t_R _34037_ (.A(_02349_),
    .Y(_17448_));
 INVx1_ASAP7_75t_R _34038_ (.A(_18309_),
    .Y(_17728_));
 INVx1_ASAP7_75t_R _34039_ (.A(_18317_),
    .Y(_17727_));
 INVx1_ASAP7_75t_R _34040_ (.A(_18120_),
    .Y(_17351_));
 INVx1_ASAP7_75t_R _34041_ (.A(_18267_),
    .Y(_17639_));
 INVx1_ASAP7_75t_R _34042_ (.A(_18144_),
    .Y(_17350_));
 INVx1_ASAP7_75t_R _34043_ (.A(_01390_),
    .Y(_16815_));
 INVx1_ASAP7_75t_R _34044_ (.A(_02315_),
    .Y(_16835_));
 INVx1_ASAP7_75t_R _34045_ (.A(_01406_),
    .Y(_16838_));
 INVx1_ASAP7_75t_R _34046_ (.A(_01417_),
    .Y(_16837_));
 INVx1_ASAP7_75t_R _34047_ (.A(_18285_),
    .Y(_17638_));
 INVx1_ASAP7_75t_R _34048_ (.A(_18086_),
    .Y(_17292_));
 INVx1_ASAP7_75t_R _34049_ (.A(_18112_),
    .Y(_17291_));
 INVx1_ASAP7_75t_R _34050_ (.A(_18286_),
    .Y(_17669_));
 INVx1_ASAP7_75t_R _34051_ (.A(_18301_),
    .Y(_17668_));
 INVx1_ASAP7_75t_R _34052_ (.A(_18113_),
    .Y(_17339_));
 INVx1_ASAP7_75t_R _34053_ (.A(_17910_),
    .Y(_16863_));
 INVx1_ASAP7_75t_R _34054_ (.A(_18142_),
    .Y(_17338_));
 INVx1_ASAP7_75t_R _34055_ (.A(_00023_),
    .Y(_17115_));
 INVx1_ASAP7_75t_R _34056_ (.A(_02341_),
    .Y(_17169_));
 INVx1_ASAP7_75t_R _34057_ (.A(_18145_),
    .Y(_17400_));
 INVx1_ASAP7_75t_R _34058_ (.A(_18247_),
    .Y(_17604_));
 INVx1_ASAP7_75t_R _34059_ (.A(_18266_),
    .Y(_17603_));
 INVx1_ASAP7_75t_R _34060_ (.A(_18209_),
    .Y(_17529_));
 INVx1_ASAP7_75t_R _34061_ (.A(_18227_),
    .Y(_17528_));
 INVx1_ASAP7_75t_R _34062_ (.A(_18268_),
    .Y(_17641_));
 INVx1_ASAP7_75t_R _34063_ (.A(_18284_),
    .Y(_17640_));
 INVx1_ASAP7_75t_R _34064_ (.A(_18287_),
    .Y(_17671_));
 INVx1_ASAP7_75t_R _34065_ (.A(_01399_),
    .Y(_17883_));
 INVx1_ASAP7_75t_R _34066_ (.A(_02318_),
    .Y(_16851_));
 INVx1_ASAP7_75t_R _34067_ (.A(_18303_),
    .Y(_17701_));
 INVx1_ASAP7_75t_R _34068_ (.A(_18310_),
    .Y(_17700_));
 INVx1_ASAP7_75t_R _34069_ (.A(_18311_),
    .Y(_17732_));
 INVx1_ASAP7_75t_R _34070_ (.A(_18319_),
    .Y(_17731_));
 INVx1_ASAP7_75t_R _34071_ (.A(_01413_),
    .Y(_16853_));
 INVx1_ASAP7_75t_R _34072_ (.A(_01422_),
    .Y(_16852_));
 INVx1_ASAP7_75t_R _34073_ (.A(_18316_),
    .Y(_17745_));
 INVx2_ASAP7_75t_R _34074_ (.A(net295),
    .Y(_17556_));
 INVx2_ASAP7_75t_R _34075_ (.A(net2150),
    .Y(_17555_));
 INVx1_ASAP7_75t_R _34076_ (.A(_18058_),
    .Y(_17230_));
 INVx1_ASAP7_75t_R _34077_ (.A(_18083_),
    .Y(_17229_));
 INVx1_ASAP7_75t_R _34078_ (.A(_18084_),
    .Y(_17287_));
 INVx1_ASAP7_75t_R _34079_ (.A(_18110_),
    .Y(_17286_));
 INVx1_ASAP7_75t_R _34080_ (.A(_18233_),
    .Y(_17579_));
 INVx1_ASAP7_75t_R _34081_ (.A(_18251_),
    .Y(_17578_));
 INVx1_ASAP7_75t_R _34082_ (.A(_18255_),
    .Y(_17621_));
 INVx1_ASAP7_75t_R _34083_ (.A(_18273_),
    .Y(_17620_));
 INVx1_ASAP7_75t_R _34084_ (.A(_18238_),
    .Y(_17585_));
 INVx1_ASAP7_75t_R _34085_ (.A(_18257_),
    .Y(_17584_));
 INVx1_ASAP7_75t_R _34086_ (.A(_18258_),
    .Y(_17622_));
 INVx1_ASAP7_75t_R _34087_ (.A(_18239_),
    .Y(_17587_));
 INVx1_ASAP7_75t_R _34088_ (.A(_18256_),
    .Y(_17586_));
 INVx1_ASAP7_75t_R _34089_ (.A(_18259_),
    .Y(_17624_));
 INVx1_ASAP7_75t_R _34090_ (.A(_18277_),
    .Y(_17623_));
 INVx1_ASAP7_75t_R _34091_ (.A(_18242_),
    .Y(_17589_));
 INVx1_ASAP7_75t_R _34092_ (.A(_18243_),
    .Y(_17591_));
 INVx1_ASAP7_75t_R _34093_ (.A(_18260_),
    .Y(_17590_));
 INVx1_ASAP7_75t_R _34094_ (.A(_18261_),
    .Y(_17628_));
 INVx1_ASAP7_75t_R _34095_ (.A(_18279_),
    .Y(_17627_));
 INVx1_ASAP7_75t_R _34096_ (.A(_18245_),
    .Y(_17595_));
 INVx1_ASAP7_75t_R _34097_ (.A(_18262_),
    .Y(_17594_));
 INVx1_ASAP7_75t_R _34098_ (.A(_17906_),
    .Y(_16885_));
 INVx1_ASAP7_75t_R _34099_ (.A(_17922_),
    .Y(_16884_));
 INVx1_ASAP7_75t_R _34100_ (.A(_17895_),
    .Y(_16858_));
 INVx1_ASAP7_75t_R _34101_ (.A(_17907_),
    .Y(_16857_));
 INVx1_ASAP7_75t_R _34102_ (.A(_18226_),
    .Y(_17566_));
 INVx1_ASAP7_75t_R _34103_ (.A(_18246_),
    .Y(_17565_));
 INVx1_ASAP7_75t_R _34104_ (.A(_18073_),
    .Y(_17259_));
 INVx1_ASAP7_75t_R _34105_ (.A(_18074_),
    .Y(_17261_));
 INVx1_ASAP7_75t_R _34106_ (.A(_18099_),
    .Y(_17260_));
 INVx1_ASAP7_75t_R _34107_ (.A(_18103_),
    .Y(_17319_));
 INVx1_ASAP7_75t_R _34108_ (.A(_18129_),
    .Y(_17318_));
 INVx1_ASAP7_75t_R _34109_ (.A(_18079_),
    .Y(_17273_));
 INVx1_ASAP7_75t_R _34110_ (.A(_18104_),
    .Y(_17272_));
 INVx1_ASAP7_75t_R _34111_ (.A(_18114_),
    .Y(_17341_));
 INVx1_ASAP7_75t_R _34112_ (.A(_18139_),
    .Y(_17340_));
 INVx1_ASAP7_75t_R _34113_ (.A(_18271_),
    .Y(_17644_));
 INVx1_ASAP7_75t_R _34114_ (.A(_18289_),
    .Y(_17643_));
 INVx1_ASAP7_75t_R _34115_ (.A(_18146_),
    .Y(_17402_));
 INVx1_ASAP7_75t_R _34116_ (.A(_18171_),
    .Y(_17401_));
 INVx1_ASAP7_75t_R _34117_ (.A(_18250_),
    .Y(_17611_));
 INVx1_ASAP7_75t_R _34118_ (.A(_18269_),
    .Y(_17610_));
 INVx1_ASAP7_75t_R _34119_ (.A(_18169_),
    .Y(_17440_));
 INVx1_ASAP7_75t_R _34120_ (.A(_18170_),
    .Y(_17442_));
 INVx1_ASAP7_75t_R _34121_ (.A(_18189_),
    .Y(_17441_));
 INVx1_ASAP7_75t_R _34122_ (.A(_18272_),
    .Y(_17646_));
 INVx1_ASAP7_75t_R _34123_ (.A(_18288_),
    .Y(_17645_));
 INVx1_ASAP7_75t_R _34124_ (.A(_18190_),
    .Y(_17490_));
 INVx1_ASAP7_75t_R _34125_ (.A(_18210_),
    .Y(_17489_));
 INVx1_ASAP7_75t_R _34126_ (.A(_18290_),
    .Y(_17672_));
 INVx1_ASAP7_75t_R _34127_ (.A(_18305_),
    .Y(_17705_));
 INVx1_ASAP7_75t_R _34128_ (.A(_18321_),
    .Y(_17734_));
 INVx1_ASAP7_75t_R _34129_ (.A(_18304_),
    .Y(_17673_));
 INVx1_ASAP7_75t_R _34130_ (.A(_18291_),
    .Y(_17674_));
 INVx1_ASAP7_75t_R _34131_ (.A(_18312_),
    .Y(_17704_));
 INVx1_ASAP7_75t_R _34132_ (.A(_18032_),
    .Y(_17120_));
 INVx1_ASAP7_75t_R _34133_ (.A(_18008_),
    .Y(_17106_));
 INVx1_ASAP7_75t_R _34134_ (.A(_18026_),
    .Y(_17105_));
 INVx1_ASAP7_75t_R _34135_ (.A(_00013_),
    .Y(_17001_));
 INVx1_ASAP7_75t_R _34136_ (.A(_18009_),
    .Y(_17111_));
 INVx1_ASAP7_75t_R _34137_ (.A(_18028_),
    .Y(_17110_));
 INVx1_ASAP7_75t_R _34138_ (.A(_01389_),
    .Y(_17874_));
 INVx1_ASAP7_75t_R _34139_ (.A(_02314_),
    .Y(_17873_));
 INVx1_ASAP7_75t_R _34140_ (.A(_01402_),
    .Y(_17886_));
 INVx1_ASAP7_75t_R _34141_ (.A(_17877_),
    .Y(_16791_));
 INVx1_ASAP7_75t_R _34142_ (.A(_01394_),
    .Y(_16819_));
 INVx1_ASAP7_75t_R _34143_ (.A(_01407_),
    .Y(_16818_));
 INVx1_ASAP7_75t_R _34144_ (.A(_01391_),
    .Y(_16795_));
 INVx1_ASAP7_75t_R _34145_ (.A(_01384_),
    .Y(_16804_));
 INVx2_ASAP7_75t_R _34146_ (.A(_01397_),
    .Y(_16803_));
 INVx1_ASAP7_75t_R _34147_ (.A(_01388_),
    .Y(_16808_));
 INVx1_ASAP7_75t_R _34148_ (.A(_01396_),
    .Y(_16822_));
 INVx1_ASAP7_75t_R _34149_ (.A(_01409_),
    .Y(_16821_));
 INVx1_ASAP7_75t_R _34150_ (.A(_00027_),
    .Y(_17131_));
 INVx1_ASAP7_75t_R _34151_ (.A(_01404_),
    .Y(_17892_));
 INVx1_ASAP7_75t_R _34152_ (.A(_01374_),
    .Y(_16781_));
 INVx1_ASAP7_75t_R _34153_ (.A(_01383_),
    .Y(_16780_));
 INVx1_ASAP7_75t_R _34154_ (.A(_01377_),
    .Y(_16787_));
 INVx1_ASAP7_75t_R _34155_ (.A(_00012_),
    .Y(_16999_));
 INVx1_ASAP7_75t_R _34156_ (.A(_18293_),
    .Y(_17678_));
 INVx1_ASAP7_75t_R _34157_ (.A(_18306_),
    .Y(_17677_));
 FAx1_ASAP7_75t_R _34158_ (.SN(\ex_block_i.alu_adder_result_ex_o[1] ),
    .A(_16714_),
    .B(_16715_),
    .CI(_16716_),
    .CON(_02222_));
 FAx1_ASAP7_75t_R _34159_ (.SN(\ex_block_i.alu_adder_result_ex_o[0] ),
    .A(_16718_),
    .B(_16719_),
    .CI(_14002_),
    .CON(_17757_));
 FAx1_ASAP7_75t_R _34160_ (.SN(net174),
    .A(_16722_),
    .B(_16723_),
    .CI(_16724_),
    .CON(_02223_));
 FAx1_ASAP7_75t_R _34161_ (.SN(net176),
    .A(_16725_),
    .B(_16726_),
    .CI(_16727_),
    .CON(_02224_));
 FAx1_ASAP7_75t_R _34162_ (.SN(_00676_),
    .A(_16728_),
    .B(_16729_),
    .CI(_16730_),
    .CON(_00679_));
 FAx1_ASAP7_75t_R _34163_ (.SN(net180),
    .A(_16731_),
    .B(_16732_),
    .CI(_16733_),
    .CON(_02225_));
 FAx1_ASAP7_75t_R _34164_ (.SN(net152),
    .A(_16734_),
    .B(_16735_),
    .CI(_16736_),
    .CON(_02226_));
 FAx1_ASAP7_75t_R _34165_ (.SN(net154),
    .A(_16737_),
    .B(_16738_),
    .CI(_16739_),
    .CON(_02227_));
 FAx1_ASAP7_75t_R _34166_ (.SN(_00785_),
    .A(_16740_),
    .B(_16741_),
    .CI(_16742_),
    .CON(_00818_));
 FAx1_ASAP7_75t_R _34167_ (.SN(net158),
    .A(_16743_),
    .B(_16744_),
    .CI(_16745_),
    .CON(_02228_));
 FAx1_ASAP7_75t_R _34168_ (.SN(net160),
    .A(_16746_),
    .B(_16747_),
    .CI(_16748_),
    .CON(_02229_));
 FAx1_ASAP7_75t_R _34169_ (.SN(net162),
    .A(_16749_),
    .B(_16750_),
    .CI(_16751_),
    .CON(_01014_));
 FAx1_ASAP7_75t_R _34170_ (.SN(net164),
    .A(_16752_),
    .B(_16753_),
    .CI(_16754_),
    .CON(_02230_));
 FAx1_ASAP7_75t_R _34171_ (.SN(net166),
    .A(_16755_),
    .B(_16756_),
    .CI(_16757_),
    .CON(_01145_));
 FAx1_ASAP7_75t_R _34172_ (.SN(net168),
    .A(_16758_),
    .B(_16759_),
    .CI(_16760_),
    .CON(_01211_));
 FAx1_ASAP7_75t_R _34173_ (.SN(net170),
    .A(_16761_),
    .B(_16762_),
    .CI(_16763_),
    .CON(_01277_));
 FAx1_ASAP7_75t_R _34174_ (.SN(_17837_),
    .A(_16764_),
    .B(_16765_),
    .CI(_16766_),
    .CON(_17848_));
 FAx1_ASAP7_75t_R _34175_ (.SN(_17847_),
    .A(_16767_),
    .B(_16768_),
    .CI(_16769_),
    .CON(_17861_));
 FAx1_ASAP7_75t_R _34176_ (.SN(_02231_),
    .A(_16770_),
    .B(_16771_),
    .CI(_16772_),
    .CON(_17868_));
 FAx1_ASAP7_75t_R _34177_ (.SN(_17860_),
    .A(_16774_),
    .B(_16775_),
    .CI(_16776_),
    .CON(_16794_));
 FAx1_ASAP7_75t_R _34178_ (.SN(_01374_),
    .A(_16777_),
    .B(_16778_),
    .CI(_16779_),
    .CON(_01383_));
 FAx1_ASAP7_75t_R _34179_ (.SN(_01376_),
    .A(_16782_),
    .B(_16783_),
    .CI(_16773_),
    .CON(_01387_));
 FAx1_ASAP7_75t_R _34180_ (.SN(_01377_),
    .A(_16784_),
    .B(_16785_),
    .CI(_16786_),
    .CON(_16814_));
 FAx1_ASAP7_75t_R _34181_ (.SN(_16793_),
    .A(_16788_),
    .B(_16789_),
    .CI(_16790_),
    .CON(_17877_));
 FAx1_ASAP7_75t_R _34182_ (.SN(_01379_),
    .A(_16792_),
    .B(_16793_),
    .CI(_16794_),
    .CON(_01391_));
 FAx1_ASAP7_75t_R _34183_ (.SN(_01382_),
    .A(_16797_),
    .B(_16798_),
    .CI(_16799_),
    .CON(_01395_));
 FAx1_ASAP7_75t_R _34184_ (.SN(_01384_),
    .A(_16801_),
    .B(_16780_),
    .CI(_16802_),
    .CON(_01397_));
 FAx1_ASAP7_75t_R _34185_ (.SN(_01388_),
    .A(_16805_),
    .B(_16806_),
    .CI(_16807_),
    .CON(_16833_));
 FAx1_ASAP7_75t_R _34186_ (.SN(_17876_),
    .A(_16809_),
    .B(_16810_),
    .CI(_16811_),
    .CON(_17889_));
 FAx1_ASAP7_75t_R _34187_ (.SN(_17878_),
    .A(_16814_),
    .B(_16813_),
    .CI(_16791_),
    .CON(_17891_));
 FAx1_ASAP7_75t_R _34188_ (.SN(_01394_),
    .A(_16815_),
    .B(_16816_),
    .CI(_16817_),
    .CON(_01407_));
 FAx1_ASAP7_75t_R _34189_ (.SN(_01396_),
    .A(_16819_),
    .B(_16800_),
    .CI(_16820_),
    .CON(_01409_));
 FAx1_ASAP7_75t_R _34190_ (.SN(_02233_),
    .A(_16822_),
    .B(_16803_),
    .CI(_16823_),
    .CON(_02232_));
 FAx1_ASAP7_75t_R _34191_ (.SN(_01400_),
    .A(_16824_),
    .B(_16825_),
    .CI(_16826_),
    .CON(_16859_));
 FAx1_ASAP7_75t_R _34192_ (.SN(_17888_),
    .A(_16828_),
    .B(_16829_),
    .CI(_16830_),
    .CON(_17896_));
 FAx1_ASAP7_75t_R _34193_ (.SN(_17890_),
    .A(_16833_),
    .B(_16832_),
    .CI(_16812_),
    .CON(_17898_));
 FAx1_ASAP7_75t_R _34194_ (.SN(_01406_),
    .A(_16834_),
    .B(_16835_),
    .CI(_16836_),
    .CON(_01417_));
 FAx1_ASAP7_75t_R _34195_ (.SN(_01408_),
    .A(_16838_),
    .B(_16818_),
    .CI(_16839_),
    .CON(_01419_));
 FAx1_ASAP7_75t_R _34196_ (.SN(_16850_),
    .A(_16842_),
    .B(_16843_),
    .CI(_16844_),
    .CON(_17903_));
 FAx1_ASAP7_75t_R _34197_ (.SN(_01412_),
    .A(_16846_),
    .B(_16847_),
    .CI(_16848_),
    .CON(_16886_));
 FAx1_ASAP7_75t_R _34198_ (.SN(_01413_),
    .A(_16850_),
    .B(_16851_),
    .CI(_16849_),
    .CON(_01422_));
 FAx1_ASAP7_75t_R _34199_ (.SN(_17895_),
    .A(_16854_),
    .B(_16855_),
    .CI(_16856_),
    .CON(_17907_));
 FAx1_ASAP7_75t_R _34200_ (.SN(_17897_),
    .A(_16859_),
    .B(_16858_),
    .CI(_16831_),
    .CON(_17909_));
 FAx1_ASAP7_75t_R _34201_ (.SN(_16866_),
    .A(_16860_),
    .B(_16861_),
    .CI(_16862_),
    .CON(_17910_));
 FAx1_ASAP7_75t_R _34202_ (.SN(_01416_),
    .A(_16864_),
    .B(_16865_),
    .CI(_16866_),
    .CON(_16895_));
 FAx1_ASAP7_75t_R _34203_ (.SN(_01418_),
    .A(_16867_),
    .B(_16837_),
    .CI(_16868_),
    .CON(_01425_));
 FAx1_ASAP7_75t_R _34204_ (.SN(_02235_),
    .A(_16870_),
    .B(_16840_),
    .CI(_16871_),
    .CON(_02234_));
 FAx1_ASAP7_75t_R _34205_ (.SN(_17902_),
    .A(_16872_),
    .B(_16873_),
    .CI(_16874_),
    .CON(_17918_));
 FAx1_ASAP7_75t_R _34206_ (.SN(_16880_),
    .A(_16877_),
    .B(_16878_),
    .CI(_16879_),
    .CON(_16914_));
 FAx1_ASAP7_75t_R _34207_ (.SN(_17904_),
    .A(_16876_),
    .B(_16845_),
    .CI(_16880_),
    .CON(_17920_));
 FAx1_ASAP7_75t_R _34208_ (.SN(_17906_),
    .A(_16881_),
    .B(_16882_),
    .CI(_16883_),
    .CON(_17922_));
 FAx1_ASAP7_75t_R _34209_ (.SN(_17908_),
    .A(_16886_),
    .B(_16885_),
    .CI(_16857_),
    .CON(_17924_));
 FAx1_ASAP7_75t_R _34210_ (.SN(_16893_),
    .A(_16887_),
    .B(_16888_),
    .CI(_16889_),
    .CON(_17925_));
 FAx1_ASAP7_75t_R _34211_ (.SN(_16894_),
    .A(_16891_),
    .B(_16892_),
    .CI(_16893_),
    .CON(_16922_));
 FAx1_ASAP7_75t_R _34212_ (.SN(net2251),
    .A(_16894_),
    .B(_16895_),
    .CI(_16863_),
    .CON(_16924_));
 FAx1_ASAP7_75t_R _34213_ (.SN(_17917_),
    .A(_16896_),
    .B(_16897_),
    .CI(_16898_),
    .CON(_17930_));
 FAx1_ASAP7_75t_R _34214_ (.SN(_16904_),
    .A(_16901_),
    .B(_16902_),
    .CI(_16903_),
    .CON(_16947_));
 FAx1_ASAP7_75t_R _34215_ (.SN(_17919_),
    .A(_16900_),
    .B(_16875_),
    .CI(_16904_),
    .CON(_17932_));
 FAx1_ASAP7_75t_R _34216_ (.SN(_01431_),
    .A(_16905_),
    .B(_16906_),
    .CI(_16907_),
    .CON(_16954_));
 FAx1_ASAP7_75t_R _34217_ (.SN(_17921_),
    .A(_16909_),
    .B(_16910_),
    .CI(_16911_),
    .CON(_17934_));
 FAx1_ASAP7_75t_R _34218_ (.SN(_17923_),
    .A(_16914_),
    .B(_16913_),
    .CI(_16884_),
    .CON(_17936_));
 FAx1_ASAP7_75t_R _34219_ (.SN(_16920_),
    .A(_16915_),
    .B(_16916_),
    .CI(_16917_),
    .CON(_17939_));
 FAx1_ASAP7_75t_R _34220_ (.SN(_16921_),
    .A(_16908_),
    .B(_16919_),
    .CI(_16920_),
    .CON(_16957_));
 FAx1_ASAP7_75t_R _34221_ (.SN(_16923_),
    .A(_16921_),
    .B(_16922_),
    .CI(_16890_),
    .CON(_17941_));
 FAx1_ASAP7_75t_R _34222_ (.SN(_02237_),
    .A(net2169),
    .B(net2170),
    .CI(_16925_),
    .CON(_02236_));
 FAx1_ASAP7_75t_R _34223_ (.SN(_17926_),
    .A(_16926_),
    .B(_16927_),
    .CI(_16928_),
    .CON(_17946_));
 FAx1_ASAP7_75t_R _34224_ (.SN(_17929_),
    .A(_16929_),
    .B(_16930_),
    .CI(_16931_),
    .CON(_17949_));
 FAx1_ASAP7_75t_R _34225_ (.SN(_16937_),
    .A(_16934_),
    .B(_16935_),
    .CI(_16936_),
    .CON(_16981_));
 FAx1_ASAP7_75t_R _34226_ (.SN(_17931_),
    .A(_16933_),
    .B(_16899_),
    .CI(_16937_),
    .CON(_17951_));
 FAx1_ASAP7_75t_R _34227_ (.SN(_16953_),
    .A(_16939_),
    .B(_16940_),
    .CI(_16941_),
    .CON(_16988_));
 FAx1_ASAP7_75t_R _34228_ (.SN(_17933_),
    .A(_16942_),
    .B(_16943_),
    .CI(_16944_),
    .CON(_17953_));
 FAx1_ASAP7_75t_R _34229_ (.SN(_17935_),
    .A(_16947_),
    .B(_16946_),
    .CI(_16912_),
    .CON(_17955_));
 FAx1_ASAP7_75t_R _34230_ (.SN(_17937_),
    .A(_16948_),
    .B(_16949_),
    .CI(_16950_),
    .CON(_17959_));
 FAx1_ASAP7_75t_R _34231_ (.SN(_17938_),
    .A(_16953_),
    .B(_16954_),
    .CI(_16952_),
    .CON(_17958_));
 FAx1_ASAP7_75t_R _34232_ (.SN(_17940_),
    .A(_16956_),
    .B(_16957_),
    .CI(_16918_),
    .CON(_16993_));
 FAx1_ASAP7_75t_R _34233_ (.SN(_17945_),
    .A(_16958_),
    .B(_16959_),
    .CI(_16960_),
    .CON(_17965_));
 FAx1_ASAP7_75t_R _34234_ (.SN(_17948_),
    .A(_16961_),
    .B(_16962_),
    .CI(_16963_),
    .CON(_17966_));
 FAx1_ASAP7_75t_R _34235_ (.SN(_16969_),
    .A(_16966_),
    .B(_16967_),
    .CI(_16968_),
    .CON(_17021_));
 FAx1_ASAP7_75t_R _34236_ (.SN(_17950_),
    .A(_16965_),
    .B(_16932_),
    .CI(_16969_),
    .CON(_17969_));
 FAx1_ASAP7_75t_R _34237_ (.SN(_16975_),
    .A(_16972_),
    .B(_16971_),
    .CI(_16938_),
    .CON(_17023_));
 FAx1_ASAP7_75t_R _34238_ (.SN(_16987_),
    .A(_16973_),
    .B(_16974_),
    .CI(_16975_),
    .CON(_17027_));
 FAx1_ASAP7_75t_R _34239_ (.SN(_17952_),
    .A(_16976_),
    .B(_16977_),
    .CI(_16978_),
    .CON(_17971_));
 FAx1_ASAP7_75t_R _34240_ (.SN(_17954_),
    .A(_16981_),
    .B(_16980_),
    .CI(_16945_),
    .CON(_17973_));
 FAx1_ASAP7_75t_R _34241_ (.SN(_17956_),
    .A(_16982_),
    .B(_16983_),
    .CI(_16984_),
    .CON(_17976_));
 FAx1_ASAP7_75t_R _34242_ (.SN(_17957_),
    .A(_16987_),
    .B(_16988_),
    .CI(_16986_),
    .CON(_17974_));
 FAx1_ASAP7_75t_R _34243_ (.SN(_16991_),
    .A(_16990_),
    .B(_16955_),
    .CI(_16951_),
    .CON(_17977_));
 FAx1_ASAP7_75t_R _34244_ (.SN(_02239_),
    .A(net2168),
    .B(_16992_),
    .CI(_16993_),
    .CON(_02238_));
 FAx1_ASAP7_75t_R _34245_ (.SN(_17964_),
    .A(_16994_),
    .B(_16995_),
    .CI(_16996_),
    .CON(_17982_));
 FAx1_ASAP7_75t_R _34246_ (.SN(_00013_),
    .A(_16998_),
    .B(_16999_),
    .CI(_17000_),
    .CON(_17057_));
 FAx1_ASAP7_75t_R _34247_ (.SN(_17967_),
    .A(_17002_),
    .B(_17003_),
    .CI(_17004_),
    .CON(_17983_));
 FAx1_ASAP7_75t_R _34248_ (.SN(_17010_),
    .A(_17007_),
    .B(_17008_),
    .CI(_17009_),
    .CON(_17066_));
 FAx1_ASAP7_75t_R _34249_ (.SN(_17968_),
    .A(_16964_),
    .B(_17010_),
    .CI(_17006_),
    .CON(_17986_));
 FAx1_ASAP7_75t_R _34250_ (.SN(_17015_),
    .A(_16970_),
    .B(_17013_),
    .CI(_17012_),
    .CON(_17067_));
 FAx1_ASAP7_75t_R _34251_ (.SN(_17026_),
    .A(_17014_),
    .B(_17015_),
    .CI(_17001_),
    .CON(_17070_));
 FAx1_ASAP7_75t_R _34252_ (.SN(_17970_),
    .A(_17016_),
    .B(_17017_),
    .CI(_17018_),
    .CON(_17990_));
 FAx1_ASAP7_75t_R _34253_ (.SN(_17972_),
    .A(_17020_),
    .B(_17021_),
    .CI(_16979_),
    .CON(_17991_));
 FAx1_ASAP7_75t_R _34254_ (.SN(_17025_),
    .A(_17022_),
    .B(_17023_),
    .CI(_17024_),
    .CON(_17074_));
 FAx1_ASAP7_75t_R _34255_ (.SN(_17975_),
    .A(_17025_),
    .B(_17026_),
    .CI(_17027_),
    .CON(_17994_));
 FAx1_ASAP7_75t_R _34256_ (.SN(_17978_),
    .A(_16989_),
    .B(_16985_),
    .CI(_17029_),
    .CON(_17076_));
 FAx1_ASAP7_75t_R _34257_ (.SN(_17980_),
    .A(_17030_),
    .B(_17031_),
    .CI(_17032_),
    .CON(_17999_));
 FAx1_ASAP7_75t_R _34258_ (.SN(_17981_),
    .A(_17034_),
    .B(_17035_),
    .CI(_17036_),
    .CON(_18000_));
 FAx1_ASAP7_75t_R _34259_ (.SN(_17042_),
    .A(_17039_),
    .B(_16997_),
    .CI(_17038_),
    .CON(_18004_));
 FAx1_ASAP7_75t_R _34260_ (.SN(_17058_),
    .A(_17041_),
    .B(_17042_),
    .CI(_17043_),
    .CON(_17103_));
 FAx1_ASAP7_75t_R _34261_ (.SN(_17984_),
    .A(_17044_),
    .B(_17045_),
    .CI(_17046_),
    .CON(_18001_));
 FAx1_ASAP7_75t_R _34262_ (.SN(_17052_),
    .A(_17049_),
    .B(_17050_),
    .CI(_17051_),
    .CON(_17112_));
 FAx1_ASAP7_75t_R _34263_ (.SN(_17985_),
    .A(_17052_),
    .B(_17005_),
    .CI(_17048_),
    .CON(_18005_));
 FAx1_ASAP7_75t_R _34264_ (.SN(_17987_),
    .A(_17054_),
    .B(_17011_),
    .CI(_17055_),
    .CON(_17113_));
 FAx1_ASAP7_75t_R _34265_ (.SN(_17988_),
    .A(_17057_),
    .B(_17056_),
    .CI(_17058_),
    .CON(_18007_));
 FAx1_ASAP7_75t_R _34266_ (.SN(_17989_),
    .A(_17061_),
    .B(_17062_),
    .CI(_17063_),
    .CON(_18010_));
 FAx1_ASAP7_75t_R _34267_ (.SN(_17992_),
    .A(_17066_),
    .B(_17065_),
    .CI(_17019_),
    .CON(_18011_));
 FAx1_ASAP7_75t_R _34268_ (.SN(_17071_),
    .A(_17067_),
    .B(_17068_),
    .CI(_17069_),
    .CON(_17119_));
 FAx1_ASAP7_75t_R _34269_ (.SN(_17993_),
    .A(_17060_),
    .B(_17070_),
    .CI(_17071_),
    .CON(_18013_));
 FAx1_ASAP7_75t_R _34270_ (.SN(_17077_),
    .A(_17073_),
    .B(_17028_),
    .CI(_17074_),
    .CON(_18015_));
 FAx1_ASAP7_75t_R _34271_ (.SN(_02241_),
    .A(_17075_),
    .B(net2166),
    .CI(net2167),
    .CON(_02240_));
 FAx1_ASAP7_75t_R _34272_ (.SN(_00021_),
    .A(_17078_),
    .B(_17079_),
    .CI(_17080_),
    .CON(_17137_));
 FAx1_ASAP7_75t_R _34273_ (.SN(_17998_),
    .A(_17082_),
    .B(_17083_),
    .CI(_17084_),
    .CON(_18018_));
 FAx1_ASAP7_75t_R _34274_ (.SN(_17090_),
    .A(_17086_),
    .B(_17037_),
    .CI(_17033_),
    .CON(_18021_));
 FAx1_ASAP7_75t_R _34275_ (.SN(_17104_),
    .A(_17088_),
    .B(_17089_),
    .CI(_17090_),
    .CON(_17154_));
 FAx1_ASAP7_75t_R _34276_ (.SN(_18002_),
    .A(_17091_),
    .B(_17092_),
    .CI(_17093_),
    .CON(_18020_));
 FAx1_ASAP7_75t_R _34277_ (.SN(_17099_),
    .A(_17096_),
    .B(_17097_),
    .CI(_17098_),
    .CON(_17163_));
 FAx1_ASAP7_75t_R _34278_ (.SN(_18003_),
    .A(_17099_),
    .B(_17047_),
    .CI(_17095_),
    .CON(_18023_));
 FAx1_ASAP7_75t_R _34279_ (.SN(_18006_),
    .A(_17053_),
    .B(_17101_),
    .CI(_17040_),
    .CON(_17168_));
 FAx1_ASAP7_75t_R _34280_ (.SN(_18008_),
    .A(_17102_),
    .B(_17103_),
    .CI(_17104_),
    .CON(_18026_));
 FAx1_ASAP7_75t_R _34281_ (.SN(_18009_),
    .A(_17107_),
    .B(_17108_),
    .CI(_17109_),
    .CON(_18028_));
 FAx1_ASAP7_75t_R _34282_ (.SN(_18012_),
    .A(_17111_),
    .B(_17064_),
    .CI(_17112_),
    .CON(_17165_));
 FAx1_ASAP7_75t_R _34283_ (.SN(_17116_),
    .A(_17113_),
    .B(_17114_),
    .CI(_17115_),
    .CON(_17173_));
 FAx1_ASAP7_75t_R _34284_ (.SN(_18014_),
    .A(_17116_),
    .B(_17059_),
    .CI(_17106_),
    .CON(_18030_));
 FAx1_ASAP7_75t_R _34285_ (.SN(_18016_),
    .A(_17119_),
    .B(_17072_),
    .CI(_17118_),
    .CON(_18032_));
 FAx1_ASAP7_75t_R _34286_ (.SN(_17129_),
    .A(_05946_),
    .B(_17122_),
    .CI(_17123_),
    .CON(_18034_));
 FAx1_ASAP7_75t_R _34287_ (.SN(_00026_),
    .A(_17125_),
    .B(_17126_),
    .CI(_17127_),
    .CON(_17192_));
 FAx1_ASAP7_75t_R _34288_ (.SN(_00027_),
    .A(_17129_),
    .B(_17130_),
    .CI(_17128_),
    .CON(_17195_));
 FAx1_ASAP7_75t_R _34289_ (.SN(_18017_),
    .A(_17132_),
    .B(_17133_),
    .CI(_17134_),
    .CON(_18037_));
 FAx1_ASAP7_75t_R _34290_ (.SN(_17140_),
    .A(_17137_),
    .B(_17136_),
    .CI(_17085_),
    .CON(_18042_));
 FAx1_ASAP7_75t_R _34291_ (.SN(_17155_),
    .A(_17131_),
    .B(_17139_),
    .CI(_17140_),
    .CON(_17210_));
 FAx1_ASAP7_75t_R _34292_ (.SN(_18019_),
    .A(_17141_),
    .B(_17142_),
    .CI(_17143_),
    .CON(_18041_));
 FAx1_ASAP7_75t_R _34293_ (.SN(_17149_),
    .A(_17146_),
    .B(_17147_),
    .CI(_17148_),
    .CON(_17218_));
 FAx1_ASAP7_75t_R _34294_ (.SN(_18022_),
    .A(_17145_),
    .B(_17094_),
    .CI(_17149_),
    .CON(_18044_));
 FAx1_ASAP7_75t_R _34295_ (.SN(_18024_),
    .A(_17087_),
    .B(_17151_),
    .CI(_17100_),
    .CON(_18052_));
 FAx1_ASAP7_75t_R _34296_ (.SN(_18025_),
    .A(_17154_),
    .B(_17153_),
    .CI(_17155_),
    .CON(_18047_));
 FAx1_ASAP7_75t_R _34297_ (.SN(_18027_),
    .A(_17158_),
    .B(_17159_),
    .CI(_17160_),
    .CON(_18049_));
 FAx1_ASAP7_75t_R _34298_ (.SN(_17164_),
    .A(_17163_),
    .B(_17162_),
    .CI(_17110_),
    .CON(_18051_));
 FAx1_ASAP7_75t_R _34299_ (.SN(_00028_),
    .A(_17164_),
    .B(_17165_),
    .CI(_17166_),
    .CON(_17220_));
 FAx1_ASAP7_75t_R _34300_ (.SN(_17170_),
    .A(_17168_),
    .B(_17167_),
    .CI(_17169_),
    .CON(_17225_));
 FAx1_ASAP7_75t_R _34301_ (.SN(_18029_),
    .A(_17157_),
    .B(_17105_),
    .CI(_17170_),
    .CON(_18055_));
 FAx1_ASAP7_75t_R _34302_ (.SN(_18031_),
    .A(_17172_),
    .B(_17117_),
    .CI(_17173_),
    .CON(_18057_));
 FAx1_ASAP7_75t_R _34303_ (.SN(_00030_),
    .A(_17174_),
    .B(_17120_),
    .CI(_17175_),
    .CON(_00033_));
 FAx1_ASAP7_75t_R _34304_ (.SN(_18033_),
    .A(_17176_),
    .B(_17177_),
    .CI(_17178_),
    .CON(_18059_));
 FAx1_ASAP7_75t_R _34305_ (.SN(_17184_),
    .A(_17181_),
    .B(_17182_),
    .CI(_17183_),
    .CON(_17242_));
 FAx1_ASAP7_75t_R _34306_ (.SN(_18035_),
    .A(_17180_),
    .B(_17124_),
    .CI(_17184_),
    .CON(_18061_));
 FAx1_ASAP7_75t_R _34307_ (.SN(_18036_),
    .A(_17187_),
    .B(_17188_),
    .CI(_17189_),
    .CON(_18063_));
 FAx1_ASAP7_75t_R _34308_ (.SN(_18038_),
    .A(_17192_),
    .B(_17191_),
    .CI(_17135_),
    .CON(_18070_));
 FAx1_ASAP7_75t_R _34309_ (.SN(_18039_),
    .A(_17186_),
    .B(_17195_),
    .CI(_17194_),
    .CON(_18066_));
 FAx1_ASAP7_75t_R _34310_ (.SN(_18040_),
    .A(_17198_),
    .B(_17199_),
    .CI(_17200_),
    .CON(_18068_));
 FAx1_ASAP7_75t_R _34311_ (.SN(_17206_),
    .A(_17203_),
    .B(_17204_),
    .CI(_17205_),
    .CON(_17266_));
 FAx1_ASAP7_75t_R _34312_ (.SN(_18043_),
    .A(_17202_),
    .B(_17144_),
    .CI(_17206_),
    .CON(_18072_));
 FAx1_ASAP7_75t_R _34313_ (.SN(_18045_),
    .A(_17138_),
    .B(_17208_),
    .CI(_17150_),
    .CON(_17268_));
 FAx1_ASAP7_75t_R _34314_ (.SN(_18046_),
    .A(_17197_),
    .B(_17210_),
    .CI(_17209_),
    .CON(_18075_));
 FAx1_ASAP7_75t_R _34315_ (.SN(_18048_),
    .A(_17213_),
    .B(_17214_),
    .CI(_17215_),
    .CON(_18076_));
 FAx1_ASAP7_75t_R _34316_ (.SN(_18050_),
    .A(_17218_),
    .B(_17217_),
    .CI(_17161_),
    .CON(_18078_));
 FAx1_ASAP7_75t_R _34317_ (.SN(_18053_),
    .A(_17152_),
    .B(_17219_),
    .CI(_17220_),
    .CON(_18081_));
 FAx1_ASAP7_75t_R _34318_ (.SN(_18054_),
    .A(_17212_),
    .B(_17156_),
    .CI(_17222_),
    .CON(_18080_));
 FAx1_ASAP7_75t_R _34319_ (.SN(_18056_),
    .A(_17224_),
    .B(_17171_),
    .CI(_17225_),
    .CON(_17275_));
 FAx1_ASAP7_75t_R _34320_ (.SN(_18058_),
    .A(_17226_),
    .B(_17227_),
    .CI(_17228_),
    .CON(_18083_));
 FAx1_ASAP7_75t_R _34321_ (.SN(_17234_),
    .A(_17231_),
    .B(_17232_),
    .CI(_17233_),
    .CON(_17293_));
 FAx1_ASAP7_75t_R _34322_ (.SN(_18060_),
    .A(_17230_),
    .B(_17179_),
    .CI(_17234_),
    .CON(_18085_));
 FAx1_ASAP7_75t_R _34323_ (.SN(_18062_),
    .A(_17237_),
    .B(_17238_),
    .CI(_17239_),
    .CON(_18087_));
 FAx1_ASAP7_75t_R _34324_ (.SN(_18064_),
    .A(_17242_),
    .B(_17241_),
    .CI(_17190_),
    .CON(_18094_));
 FAx1_ASAP7_75t_R _34325_ (.SN(_18065_),
    .A(_17236_),
    .B(_17185_),
    .CI(_17244_),
    .CON(_18090_));
 FAx1_ASAP7_75t_R _34326_ (.SN(_18067_),
    .A(_17247_),
    .B(_17248_),
    .CI(_17249_),
    .CON(_18092_));
 FAx1_ASAP7_75t_R _34327_ (.SN(_18069_),
    .A(_17252_),
    .B(_17253_),
    .CI(_17254_),
    .CON(_18100_));
 FAx1_ASAP7_75t_R _34328_ (.SN(_18071_),
    .A(_17251_),
    .B(_17201_),
    .CI(_17256_),
    .CON(_18096_));
 FAx1_ASAP7_75t_R _34329_ (.SN(_18073_),
    .A(_17193_),
    .B(_17258_),
    .CI(_17207_),
    .CON(_17314_));
 FAx1_ASAP7_75t_R _34330_ (.SN(_18074_),
    .A(_17246_),
    .B(_17196_),
    .CI(_17259_),
    .CON(_18099_));
 FAx1_ASAP7_75t_R _34331_ (.SN(_17267_),
    .A(_17166_),
    .B(_17262_),
    .CI(_17263_),
    .CON(_17313_));
 FAx1_ASAP7_75t_R _34332_ (.SN(_18077_),
    .A(_17266_),
    .B(net2128),
    .CI(_17216_),
    .CON(_18102_));
 FAx1_ASAP7_75t_R _34333_ (.SN(_17271_),
    .A(_17268_),
    .B(_17269_),
    .CI(_17270_),
    .CON(_17320_));
 FAx1_ASAP7_75t_R _34334_ (.SN(_18079_),
    .A(_17261_),
    .B(_17211_),
    .CI(_17271_),
    .CON(_18104_));
 FAx1_ASAP7_75t_R _34335_ (.SN(_17274_),
    .A(_17273_),
    .B(_17223_),
    .CI(_17221_),
    .CON(_18106_));
 FAx1_ASAP7_75t_R _34336_ (.SN(_02243_),
    .A(net2162),
    .B(_17275_),
    .CI(_17276_),
    .CON(_02242_));
 FAx1_ASAP7_75t_R _34337_ (.SN(_18082_),
    .A(_17277_),
    .B(_17278_),
    .CI(_17279_),
    .CON(_18108_));
 FAx1_ASAP7_75t_R _34338_ (.SN(_17285_),
    .A(_17282_),
    .B(_17283_),
    .CI(_17284_),
    .CON(_17337_));
 FAx1_ASAP7_75t_R _34339_ (.SN(_18084_),
    .A(_17281_),
    .B(_17229_),
    .CI(_17285_),
    .CON(_18110_));
 FAx1_ASAP7_75t_R _34340_ (.SN(_18086_),
    .A(_17288_),
    .B(_17289_),
    .CI(_17290_),
    .CON(_18112_));
 FAx1_ASAP7_75t_R _34341_ (.SN(_18088_),
    .A(_17293_),
    .B(_17292_),
    .CI(_17240_),
    .CON(_18119_));
 FAx1_ASAP7_75t_R _34342_ (.SN(_18089_),
    .A(_17287_),
    .B(_17235_),
    .CI(_17295_),
    .CON(_18115_));
 FAx1_ASAP7_75t_R _34343_ (.SN(_18091_),
    .A(_17298_),
    .B(_17299_),
    .CI(_17300_),
    .CON(_18117_));
 FAx1_ASAP7_75t_R _34344_ (.SN(_18093_),
    .A(_17303_),
    .B(_17304_),
    .CI(_17305_),
    .CON(_18125_));
 FAx1_ASAP7_75t_R _34345_ (.SN(_18095_),
    .A(_17302_),
    .B(_17250_),
    .CI(_17307_),
    .CON(_18121_));
 FAx1_ASAP7_75t_R _34346_ (.SN(_18097_),
    .A(_17243_),
    .B(_17309_),
    .CI(_17257_),
    .CON(_17355_));
 FAx1_ASAP7_75t_R _34347_ (.SN(_18098_),
    .A(_17297_),
    .B(_17245_),
    .CI(_17310_),
    .CON(_18124_));
 FAx1_ASAP7_75t_R _34348_ (.SN(_18101_),
    .A(net2127),
    .B(_17255_),
    .CI(_17313_),
    .CON(_18127_));
 FAx1_ASAP7_75t_R _34349_ (.SN(_17317_),
    .A(_17314_),
    .B(_17315_),
    .CI(_17316_),
    .CON(_17361_));
 FAx1_ASAP7_75t_R _34350_ (.SN(_18103_),
    .A(_17312_),
    .B(_17260_),
    .CI(_17317_),
    .CON(_18129_));
 FAx1_ASAP7_75t_R _34351_ (.SN(_18105_),
    .A(_17319_),
    .B(_17272_),
    .CI(_17320_),
    .CON(_17363_));
 FAx1_ASAP7_75t_R _34352_ (.SN(_18107_),
    .A(_17321_),
    .B(_17322_),
    .CI(_17323_),
    .CON(_18131_));
 FAx1_ASAP7_75t_R _34353_ (.SN(_17329_),
    .A(_17326_),
    .B(_17327_),
    .CI(_17328_),
    .CON(_17382_));
 FAx1_ASAP7_75t_R _34354_ (.SN(_18109_),
    .A(_17325_),
    .B(_17280_),
    .CI(_17329_),
    .CON(_18134_));
 FAx1_ASAP7_75t_R _34355_ (.SN(_18111_),
    .A(_17332_),
    .B(_17333_),
    .CI(_17334_),
    .CON(_18136_));
 FAx1_ASAP7_75t_R _34356_ (.SN(_18113_),
    .A(_17337_),
    .B(_17336_),
    .CI(_17291_),
    .CON(_18142_));
 FAx1_ASAP7_75t_R _34357_ (.SN(_18114_),
    .A(_17331_),
    .B(_17286_),
    .CI(_17339_),
    .CON(_18139_));
 FAx1_ASAP7_75t_R _34358_ (.SN(_18116_),
    .A(_17342_),
    .B(_17343_),
    .CI(_17344_),
    .CON(_18141_));
 FAx1_ASAP7_75t_R _34359_ (.SN(_18118_),
    .A(_17305_),
    .B(_17347_),
    .CI(_17348_),
    .CON(_17403_));
 FAx1_ASAP7_75t_R _34360_ (.SN(_18120_),
    .A(_17346_),
    .B(_17301_),
    .CI(_17349_),
    .CON(_18144_));
 FAx1_ASAP7_75t_R _34361_ (.SN(_18122_),
    .A(_17294_),
    .B(_17351_),
    .CI(_17308_),
    .CON(_17406_));
 FAx1_ASAP7_75t_R _34362_ (.SN(_18123_),
    .A(_17341_),
    .B(_17296_),
    .CI(_17352_),
    .CON(_18147_));
 FAx1_ASAP7_75t_R _34363_ (.SN(_18126_),
    .A(net2130),
    .B(net2250),
    .CI(_17306_),
    .CON(_18148_));
 FAx1_ASAP7_75t_R _34364_ (.SN(_17358_),
    .A(_17355_),
    .B(_17356_),
    .CI(_17357_),
    .CON(_17412_));
 FAx1_ASAP7_75t_R _34365_ (.SN(_18128_),
    .A(_17354_),
    .B(_17311_),
    .CI(_17358_),
    .CON(_18150_));
 FAx1_ASAP7_75t_R _34366_ (.SN(_17362_),
    .A(_17360_),
    .B(_17318_),
    .CI(_17361_),
    .CON(_18152_));
 FAx1_ASAP7_75t_R _34367_ (.SN(_02245_),
    .A(_17362_),
    .B(_17363_),
    .CI(_17364_),
    .CON(_02244_));
 FAx1_ASAP7_75t_R _34368_ (.SN(_18130_),
    .A(_17365_),
    .B(_17366_),
    .CI(_17367_),
    .CON(_18154_));
 FAx1_ASAP7_75t_R _34369_ (.SN(_18132_),
    .A(_17370_),
    .B(_17371_),
    .CI(_17372_),
    .CON(_18158_));
 FAx1_ASAP7_75t_R _34370_ (.SN(_18133_),
    .A(_17369_),
    .B(_17324_),
    .CI(_17374_),
    .CON(_18157_));
 FAx1_ASAP7_75t_R _34371_ (.SN(_18135_),
    .A(_17377_),
    .B(_17378_),
    .CI(_17379_),
    .CON(_18160_));
 FAx1_ASAP7_75t_R _34372_ (.SN(_18137_),
    .A(_17382_),
    .B(_17381_),
    .CI(_17335_),
    .CON(_18166_));
 FAx1_ASAP7_75t_R _34373_ (.SN(_18138_),
    .A(_17376_),
    .B(_17330_),
    .CI(_17384_),
    .CON(_18163_));
 FAx1_ASAP7_75t_R _34374_ (.SN(_18140_),
    .A(_17387_),
    .B(_17388_),
    .CI(_17389_),
    .CON(_18165_));
 FAx1_ASAP7_75t_R _34375_ (.SN(_17397_),
    .A(_17392_),
    .B(_17393_),
    .CI(_17394_),
    .CON(_17445_));
 FAx1_ASAP7_75t_R _34376_ (.SN(_18143_),
    .A(_17391_),
    .B(_17345_),
    .CI(net2131),
    .CON(_18168_));
 FAx1_ASAP7_75t_R _34377_ (.SN(_18145_),
    .A(_17338_),
    .B(_17399_),
    .CI(_17350_),
    .CON(_17446_));
 FAx1_ASAP7_75t_R _34378_ (.SN(_18146_),
    .A(_17386_),
    .B(_17340_),
    .CI(_17400_),
    .CON(_18171_));
 FAx1_ASAP7_75t_R _34379_ (.SN(_00042_),
    .A(_17265_),
    .B(_17264_),
    .CI(_17403_),
    .CON(_00047_));
 FAx1_ASAP7_75t_R _34380_ (.SN(_17409_),
    .A(_17406_),
    .B(_17407_),
    .CI(_17408_),
    .CON(_17452_));
 FAx1_ASAP7_75t_R _34381_ (.SN(_18149_),
    .A(_17402_),
    .B(_17353_),
    .CI(_17409_),
    .CON(_18173_));
 FAx1_ASAP7_75t_R _34382_ (.SN(_18151_),
    .A(_17411_),
    .B(_17359_),
    .CI(_17412_),
    .CON(_17454_));
 FAx1_ASAP7_75t_R _34383_ (.SN(_18153_),
    .A(_17413_),
    .B(_17414_),
    .CI(_17415_),
    .CON(_18175_));
 FAx1_ASAP7_75t_R _34384_ (.SN(_18155_),
    .A(_17418_),
    .B(_17419_),
    .CI(_17420_),
    .CON(_18179_));
 FAx1_ASAP7_75t_R _34385_ (.SN(_18156_),
    .A(_17417_),
    .B(_17368_),
    .CI(_17422_),
    .CON(_18178_));
 FAx1_ASAP7_75t_R _34386_ (.SN(_18159_),
    .A(_17425_),
    .B(_17426_),
    .CI(_17427_),
    .CON(_18181_));
 FAx1_ASAP7_75t_R _34387_ (.SN(_18161_),
    .A(_17373_),
    .B(_17429_),
    .CI(_17380_),
    .CON(_18185_));
 FAx1_ASAP7_75t_R _34388_ (.SN(_18162_),
    .A(_17424_),
    .B(_17375_),
    .CI(_17431_),
    .CON(_18184_));
 FAx1_ASAP7_75t_R _34389_ (.SN(_18164_),
    .A(_17434_),
    .B(_17435_),
    .CI(_17436_),
    .CON(_17480_));
 FAx1_ASAP7_75t_R _34390_ (.SN(_18167_),
    .A(net2132),
    .B(_17437_),
    .CI(_17390_),
    .CON(_18186_));
 FAx1_ASAP7_75t_R _34391_ (.SN(_18169_),
    .A(_17383_),
    .B(_17439_),
    .CI(_17398_),
    .CON(_17485_));
 FAx1_ASAP7_75t_R _34392_ (.SN(_18170_),
    .A(_17433_),
    .B(_17385_),
    .CI(_17440_),
    .CON(_18189_));
 FAx1_ASAP7_75t_R _34393_ (.SN(_00046_),
    .A(_17265_),
    .B(_17264_),
    .CI(_17395_),
    .CON(_00050_));
 FAx1_ASAP7_75t_R _34394_ (.SN(_17449_),
    .A(_17446_),
    .B(_17447_),
    .CI(_17448_),
    .CON(_17491_));
 FAx1_ASAP7_75t_R _34395_ (.SN(_18172_),
    .A(_17442_),
    .B(_17401_),
    .CI(_17449_),
    .CON(_18191_));
 FAx1_ASAP7_75t_R _34396_ (.SN(_17453_),
    .A(_17451_),
    .B(_17410_),
    .CI(_17452_),
    .CON(_18193_));
 FAx1_ASAP7_75t_R _34397_ (.SN(_02247_),
    .A(_17453_),
    .B(_17454_),
    .CI(_17455_),
    .CON(_02246_));
 FAx1_ASAP7_75t_R _34398_ (.SN(_18174_),
    .A(_17456_),
    .B(_17457_),
    .CI(_17458_),
    .CON(_18195_));
 FAx1_ASAP7_75t_R _34399_ (.SN(_18176_),
    .A(_17461_),
    .B(_17462_),
    .CI(_17463_),
    .CON(_18199_));
 FAx1_ASAP7_75t_R _34400_ (.SN(_18177_),
    .A(_17460_),
    .B(_17416_),
    .CI(_17465_),
    .CON(_18198_));
 FAx1_ASAP7_75t_R _34401_ (.SN(_18180_),
    .A(_17468_),
    .B(_17469_),
    .CI(_17470_),
    .CON(_18201_));
 FAx1_ASAP7_75t_R _34402_ (.SN(_18182_),
    .A(_17421_),
    .B(_17472_),
    .CI(_17428_),
    .CON(_18205_));
 FAx1_ASAP7_75t_R _34403_ (.SN(_18183_),
    .A(_17467_),
    .B(_17423_),
    .CI(_17474_),
    .CON(_18204_));
 FAx1_ASAP7_75t_R _34404_ (.SN(_17479_),
    .A(_17436_),
    .B(_17477_),
    .CI(_17478_),
    .CON(_17518_));
 FAx1_ASAP7_75t_R _34405_ (.SN(_17481_),
    .A(_17396_),
    .B(_17479_),
    .CI(_17480_),
    .CON(_17521_));
 FAx1_ASAP7_75t_R _34406_ (.SN(_18187_),
    .A(_17430_),
    .B(_17481_),
    .CI(_17438_),
    .CON(_17525_));
 FAx1_ASAP7_75t_R _34407_ (.SN(_18188_),
    .A(_17476_),
    .B(_17432_),
    .CI(_17482_),
    .CON(_18208_));
 FAx1_ASAP7_75t_R _34408_ (.SN(_17488_),
    .A(_17485_),
    .B(_17486_),
    .CI(_17487_),
    .CON(_17530_));
 FAx1_ASAP7_75t_R _34409_ (.SN(_18190_),
    .A(_17484_),
    .B(_17441_),
    .CI(_17488_),
    .CON(_18210_));
 FAx1_ASAP7_75t_R _34410_ (.SN(_18192_),
    .A(_17490_),
    .B(_17450_),
    .CI(_17491_),
    .CON(_17532_));
 FAx1_ASAP7_75t_R _34411_ (.SN(_18194_),
    .A(_17492_),
    .B(_17493_),
    .CI(_17494_),
    .CON(_18212_));
 FAx1_ASAP7_75t_R _34412_ (.SN(_18196_),
    .A(_17497_),
    .B(_17498_),
    .CI(_17499_),
    .CON(_18216_));
 FAx1_ASAP7_75t_R _34413_ (.SN(_18197_),
    .A(_17496_),
    .B(_17459_),
    .CI(_17501_),
    .CON(_18215_));
 FAx1_ASAP7_75t_R _34414_ (.SN(_18200_),
    .A(_17504_),
    .B(_17505_),
    .CI(_17506_),
    .CON(_18218_));
 FAx1_ASAP7_75t_R _34415_ (.SN(_18202_),
    .A(_17464_),
    .B(_17508_),
    .CI(_17471_),
    .CON(_18222_));
 FAx1_ASAP7_75t_R _34416_ (.SN(_18203_),
    .A(_17503_),
    .B(_17466_),
    .CI(_17510_),
    .CON(_18221_));
 FAx1_ASAP7_75t_R _34417_ (.SN(_17519_),
    .A(_17513_),
    .B(_17514_),
    .CI(_17515_),
    .CON(_17557_));
 FAx1_ASAP7_75t_R _34418_ (.SN(_17520_),
    .A(_17396_),
    .B(_17517_),
    .CI(_17518_),
    .CON(_17559_));
 FAx1_ASAP7_75t_R _34419_ (.SN(_18206_),
    .A(_17473_),
    .B(_17520_),
    .CI(_17521_),
    .CON(_17563_));
 FAx1_ASAP7_75t_R _34420_ (.SN(_18207_),
    .A(_17512_),
    .B(_17475_),
    .CI(_17522_),
    .CON(_18225_));
 FAx1_ASAP7_75t_R _34421_ (.SN(_17527_),
    .A(_17486_),
    .B(_17525_),
    .CI(_17526_),
    .CON(_17567_));
 FAx1_ASAP7_75t_R _34422_ (.SN(_18209_),
    .A(_17524_),
    .B(_17483_),
    .CI(_17527_),
    .CON(_18227_));
 FAx1_ASAP7_75t_R _34423_ (.SN(_17531_),
    .A(_17529_),
    .B(_17489_),
    .CI(_17530_),
    .CON(_18229_));
 FAx1_ASAP7_75t_R _34424_ (.SN(_02249_),
    .A(net2151),
    .B(_17532_),
    .CI(_17533_),
    .CON(_02248_));
 FAx1_ASAP7_75t_R _34425_ (.SN(_18211_),
    .A(_17534_),
    .B(_17535_),
    .CI(_17536_),
    .CON(_18231_));
 FAx1_ASAP7_75t_R _34426_ (.SN(_18213_),
    .A(_17539_),
    .B(_17540_),
    .CI(_17541_),
    .CON(_18235_));
 FAx1_ASAP7_75t_R _34427_ (.SN(_18214_),
    .A(_17538_),
    .B(_17495_),
    .CI(_17543_),
    .CON(_18234_));
 FAx1_ASAP7_75t_R _34428_ (.SN(_18217_),
    .A(_17546_),
    .B(_17547_),
    .CI(_17548_),
    .CON(_18237_));
 FAx1_ASAP7_75t_R _34429_ (.SN(_18219_),
    .A(_17500_),
    .B(_17550_),
    .CI(_17507_),
    .CON(_18241_));
 FAx1_ASAP7_75t_R _34430_ (.SN(_18220_),
    .A(_17545_),
    .B(_17502_),
    .CI(_17552_),
    .CON(_18240_));
 FAx1_ASAP7_75t_R _34431_ (.SN(_17558_),
    .A(_17396_),
    .B(_17517_),
    .CI(_17516_),
    .CON(_17588_));
 FAx1_ASAP7_75t_R _34432_ (.SN(_18223_),
    .A(_17509_),
    .B(net2193),
    .CI(_17559_),
    .CON(_17592_));
 FAx1_ASAP7_75t_R _34433_ (.SN(_18224_),
    .A(_17554_),
    .B(_17511_),
    .CI(_17560_),
    .CON(_18244_));
 FAx1_ASAP7_75t_R _34434_ (.SN(_17564_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17563_),
    .CON(_17596_));
 FAx1_ASAP7_75t_R _34435_ (.SN(_18226_),
    .A(_17562_),
    .B(_17523_),
    .CI(_17564_),
    .CON(_18246_));
 FAx1_ASAP7_75t_R _34436_ (.SN(_18228_),
    .A(_17566_),
    .B(_17528_),
    .CI(_17567_),
    .CON(_17598_));
 FAx1_ASAP7_75t_R _34437_ (.SN(_18230_),
    .A(_17568_),
    .B(_17569_),
    .CI(_17570_),
    .CON(_18248_));
 FAx1_ASAP7_75t_R _34438_ (.SN(_18232_),
    .A(_17573_),
    .B(_17574_),
    .CI(_17575_),
    .CON(_18252_));
 FAx1_ASAP7_75t_R _34439_ (.SN(_18233_),
    .A(_17572_),
    .B(_17537_),
    .CI(_17577_),
    .CON(_18251_));
 FAx1_ASAP7_75t_R _34440_ (.SN(_18236_),
    .A(_17548_),
    .B(_17580_),
    .CI(_17581_),
    .CON(_18253_));
 FAx1_ASAP7_75t_R _34441_ (.SN(_18238_),
    .A(_17542_),
    .B(_17583_),
    .CI(_17549_),
    .CON(_18257_));
 FAx1_ASAP7_75t_R _34442_ (.SN(_18239_),
    .A(_17579_),
    .B(_17544_),
    .CI(_17585_),
    .CON(_18256_));
 FAx1_ASAP7_75t_R _34443_ (.SN(_18242_),
    .A(net2195),
    .B(_17551_),
    .CI(_17588_),
    .CON(_17625_));
 FAx1_ASAP7_75t_R _34444_ (.SN(_18243_),
    .A(_17587_),
    .B(_17553_),
    .CI(_17589_),
    .CON(_18260_));
 FAx1_ASAP7_75t_R _34445_ (.SN(_17593_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17592_),
    .CON(_17629_));
 FAx1_ASAP7_75t_R _34446_ (.SN(_18245_),
    .A(_17591_),
    .B(_17561_),
    .CI(_17593_),
    .CON(_18262_));
 FAx1_ASAP7_75t_R _34447_ (.SN(_17597_),
    .A(_17595_),
    .B(_17565_),
    .CI(_17596_),
    .CON(_18264_));
 FAx1_ASAP7_75t_R _34448_ (.SN(_02251_),
    .A(_17597_),
    .B(_17598_),
    .CI(_17599_),
    .CON(_02250_));
 FAx1_ASAP7_75t_R _34449_ (.SN(_18247_),
    .A(_17600_),
    .B(_17601_),
    .CI(_17602_),
    .CON(_18266_));
 FAx1_ASAP7_75t_R _34450_ (.SN(_18249_),
    .A(_17605_),
    .B(_17606_),
    .CI(_17607_),
    .CON(_18270_));
 FAx1_ASAP7_75t_R _34451_ (.SN(_18250_),
    .A(_17604_),
    .B(_17571_),
    .CI(_17609_),
    .CON(_18269_));
 FAx1_ASAP7_75t_R _34452_ (.SN(_17617_),
    .A(_17612_),
    .B(_17613_),
    .CI(_17614_),
    .CON(_17642_));
 FAx1_ASAP7_75t_R _34453_ (.SN(_18254_),
    .A(_17576_),
    .B(net2241),
    .CI(_17582_),
    .CON(_18274_));
 FAx1_ASAP7_75t_R _34454_ (.SN(_18255_),
    .A(_17611_),
    .B(_17578_),
    .CI(_17619_),
    .CON(_18273_));
 FAx1_ASAP7_75t_R _34455_ (.SN(_18258_),
    .A(net295),
    .B(net2147),
    .CI(_17584_),
    .CON(_17650_));
 FAx1_ASAP7_75t_R _34456_ (.SN(_18259_),
    .A(_17621_),
    .B(_17586_),
    .CI(_17622_),
    .CON(_18277_));
 FAx1_ASAP7_75t_R _34457_ (.SN(_17626_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17625_),
    .CON(_17654_));
 FAx1_ASAP7_75t_R _34458_ (.SN(_18261_),
    .A(_17624_),
    .B(_17590_),
    .CI(_17626_),
    .CON(_18279_));
 FAx1_ASAP7_75t_R _34459_ (.SN(_18263_),
    .A(_17628_),
    .B(_17594_),
    .CI(_17629_),
    .CON(_17656_));
 FAx1_ASAP7_75t_R _34460_ (.SN(_18265_),
    .A(_17630_),
    .B(_17631_),
    .CI(_17632_),
    .CON(_18281_));
 FAx1_ASAP7_75t_R _34461_ (.SN(_18267_),
    .A(_17635_),
    .B(_17636_),
    .CI(_17637_),
    .CON(_18285_));
 FAx1_ASAP7_75t_R _34462_ (.SN(_18268_),
    .A(_17634_),
    .B(_17603_),
    .CI(_17639_),
    .CON(_18284_));
 FAx1_ASAP7_75t_R _34463_ (.SN(_18271_),
    .A(net2238),
    .B(_17608_),
    .CI(_17642_),
    .CON(_18289_));
 FAx1_ASAP7_75t_R _34464_ (.SN(_18272_),
    .A(_17641_),
    .B(_17610_),
    .CI(_17644_),
    .CON(_18288_));
 FAx1_ASAP7_75t_R _34465_ (.SN(_18275_),
    .A(net295),
    .B(net2147),
    .CI(_17618_),
    .CON(_17675_));
 FAx1_ASAP7_75t_R _34466_ (.SN(_18276_),
    .A(_17646_),
    .B(_17620_),
    .CI(_17647_),
    .CON(_18292_));
 FAx1_ASAP7_75t_R _34467_ (.SN(_17651_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17650_),
    .CON(_17679_));
 FAx1_ASAP7_75t_R _34468_ (.SN(_18278_),
    .A(_17649_),
    .B(_17623_),
    .CI(_17651_),
    .CON(_18294_));
 FAx1_ASAP7_75t_R _34469_ (.SN(_17655_),
    .A(_17653_),
    .B(_17627_),
    .CI(_17654_),
    .CON(_18296_));
 FAx1_ASAP7_75t_R _34470_ (.SN(_02253_),
    .A(_17655_),
    .B(_17656_),
    .CI(_17657_),
    .CON(_02252_));
 FAx1_ASAP7_75t_R _34471_ (.SN(_18280_),
    .A(_17658_),
    .B(_17659_),
    .CI(_17660_),
    .CON(_17693_));
 FAx1_ASAP7_75t_R _34472_ (.SN(_18282_),
    .A(_17637_),
    .B(_17663_),
    .CI(_17664_),
    .CON(_17694_));
 FAx1_ASAP7_75t_R _34473_ (.SN(_18283_),
    .A(_17662_),
    .B(_17633_),
    .CI(_17665_),
    .CON(_18298_));
 FAx1_ASAP7_75t_R _34474_ (.SN(_18286_),
    .A(net2240),
    .B(_17642_),
    .CI(_17638_),
    .CON(_18301_));
 FAx1_ASAP7_75t_R _34475_ (.SN(_18287_),
    .A(_17667_),
    .B(_17640_),
    .CI(_17669_),
    .CON(_18300_));
 FAx1_ASAP7_75t_R _34476_ (.SN(_18290_),
    .A(net295),
    .B(net2148),
    .CI(_17643_),
    .CON(_17702_));
 FAx1_ASAP7_75t_R _34477_ (.SN(_18291_),
    .A(_17671_),
    .B(_17645_),
    .CI(_17672_),
    .CON(_18304_));
 FAx1_ASAP7_75t_R _34478_ (.SN(_17676_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17675_),
    .CON(_17706_));
 FAx1_ASAP7_75t_R _34479_ (.SN(_18293_),
    .A(_17674_),
    .B(_17648_),
    .CI(_17676_),
    .CON(_18306_));
 FAx1_ASAP7_75t_R _34480_ (.SN(_18295_),
    .A(_17678_),
    .B(_17652_),
    .CI(_17679_),
    .CON(_17708_));
 FAx1_ASAP7_75t_R _34481_ (.SN(_17692_),
    .A(_17680_),
    .B(_17681_),
    .CI(_17682_),
    .CON(_17714_));
 FAx1_ASAP7_75t_R _34482_ (.SN(_17689_),
    .A(_17684_),
    .B(_17685_),
    .CI(_17686_),
    .CON(_17718_));
 FAx1_ASAP7_75t_R _34483_ (.SN(_18297_),
    .A(_17683_),
    .B(_17661_),
    .CI(_17689_),
    .CON(_17723_));
 FAx1_ASAP7_75t_R _34484_ (.SN(_17696_),
    .A(_17616_),
    .B(_17615_),
    .CI(_17694_),
    .CON(_17725_));
 FAx1_ASAP7_75t_R _34485_ (.SN(_18299_),
    .A(_17691_),
    .B(_17666_),
    .CI(_17696_),
    .CON(_18308_));
 FAx1_ASAP7_75t_R _34486_ (.SN(_18302_),
    .A(net295),
    .B(net2149),
    .CI(_17668_),
    .CON(_17729_));
 FAx1_ASAP7_75t_R _34487_ (.SN(_18303_),
    .A(_17698_),
    .B(_17670_),
    .CI(_17699_),
    .CON(_18310_));
 FAx1_ASAP7_75t_R _34488_ (.SN(_17703_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17702_),
    .CON(_17733_));
 FAx1_ASAP7_75t_R _34489_ (.SN(_18305_),
    .A(_17701_),
    .B(_17673_),
    .CI(_17703_),
    .CON(_18312_));
 FAx1_ASAP7_75t_R _34490_ (.SN(_17707_),
    .A(_17705_),
    .B(_17677_),
    .CI(_17706_),
    .CON(_18314_));
 FAx1_ASAP7_75t_R _34491_ (.SN(_02255_),
    .A(_17707_),
    .B(_17708_),
    .CI(_17709_),
    .CON(_02254_));
 FAx1_ASAP7_75t_R _34492_ (.SN(_17713_),
    .A(_17710_),
    .B(_17711_),
    .CI(_17712_),
    .CON(_17738_));
 FAx1_ASAP7_75t_R _34493_ (.SN(_17719_),
    .A(_17688_),
    .B(_17713_),
    .CI(_17714_),
    .CON(_17741_));
 FAx1_ASAP7_75t_R _34494_ (.SN(_17720_),
    .A(_17616_),
    .B(_17615_),
    .CI(_17687_),
    .CON(_17742_));
 FAx1_ASAP7_75t_R _34495_ (.SN(_18307_),
    .A(_17719_),
    .B(_17690_),
    .CI(_17720_),
    .CON(_18315_));
 FAx1_ASAP7_75t_R _34496_ (.SN(_17726_),
    .A(_17556_),
    .B(_17555_),
    .CI(_17695_),
    .CON(_00066_));
 FAx1_ASAP7_75t_R _34497_ (.SN(_18309_),
    .A(_17722_),
    .B(_17697_),
    .CI(_17726_),
    .CON(_18317_));
 FAx1_ASAP7_75t_R _34498_ (.SN(_17730_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17729_),
    .CON(_17748_));
 FAx1_ASAP7_75t_R _34499_ (.SN(_18311_),
    .A(_17728_),
    .B(_17700_),
    .CI(_17730_),
    .CON(_18319_));
 FAx1_ASAP7_75t_R _34500_ (.SN(_18313_),
    .A(_17732_),
    .B(_17704_),
    .CI(_17733_),
    .CON(_18321_));
 FAx1_ASAP7_75t_R _34501_ (.SN(_17737_),
    .A(_17712_),
    .B(_17735_),
    .CI(_17736_),
    .CON(_02256_));
 FAx1_ASAP7_75t_R _34502_ (.SN(_17740_),
    .A(_17688_),
    .B(_17737_),
    .CI(_17738_),
    .CON(_00068_));
 FAx1_ASAP7_75t_R _34503_ (.SN(_17743_),
    .A(_17717_),
    .B(_17739_),
    .CI(_17715_),
    .CON(_00069_));
 FAx1_ASAP7_75t_R _34504_ (.SN(_17744_),
    .A(_17556_),
    .B(_17555_),
    .CI(_17716_),
    .CON(_00070_));
 FAx1_ASAP7_75t_R _34505_ (.SN(_18316_),
    .A(_17743_),
    .B(_17721_),
    .CI(_17744_),
    .CON(_02257_));
 FAx1_ASAP7_75t_R _34506_ (.SN(_17746_),
    .A(_17486_),
    .B(_17526_),
    .CI(_17724_),
    .CON(_00071_));
 FAx1_ASAP7_75t_R _34507_ (.SN(_18318_),
    .A(_17745_),
    .B(_17727_),
    .CI(_17746_),
    .CON(_02258_));
 FAx1_ASAP7_75t_R _34508_ (.SN(_18320_),
    .A(_17747_),
    .B(_17731_),
    .CI(_17748_),
    .CON(_02259_));
 FAx1_ASAP7_75t_R _34509_ (.SN(_02261_),
    .A(_17749_),
    .B(_17734_),
    .CI(_17750_),
    .CON(_02260_));
 FAx1_ASAP7_75t_R _34510_ (.SN(_00241_),
    .A(_17751_),
    .B(_17752_),
    .CI(\cs_registers_i.pc_if_i[2] ),
    .CON(_00242_));
 HAxp5_ASAP7_75t_R _34511_ (.A(_17755_),
    .B(_17756_),
    .CON(_00664_),
    .SN(_00292_));
 HAxp5_ASAP7_75t_R _34512_ (.A(_17758_),
    .B(_17759_),
    .CON(_00667_),
    .SN(_02262_));
 HAxp5_ASAP7_75t_R _34513_ (.A(_17760_),
    .B(_17761_),
    .CON(_00669_),
    .SN(_00666_));
 HAxp5_ASAP7_75t_R _34514_ (.A(_17762_),
    .B(_17763_),
    .CON(_02263_),
    .SN(_02264_));
 HAxp5_ASAP7_75t_R _34515_ (.A(_17764_),
    .B(_17765_),
    .CON(_00673_),
    .SN(_00671_));
 HAxp5_ASAP7_75t_R _34516_ (.A(_17766_),
    .B(_17767_),
    .CON(_02265_),
    .SN(_02266_));
 HAxp5_ASAP7_75t_R _34517_ (.A(_16728_),
    .B(_16729_),
    .CON(_00678_),
    .SN(_00675_));
 HAxp5_ASAP7_75t_R _34518_ (.A(_17768_),
    .B(_17769_),
    .CON(_02267_),
    .SN(_02268_));
 HAxp5_ASAP7_75t_R _34519_ (.A(_17770_),
    .B(_17771_),
    .CON(_00683_),
    .SN(_00681_));
 HAxp5_ASAP7_75t_R _34520_ (.A(_17772_),
    .B(_17773_),
    .CON(_02269_),
    .SN(_02270_));
 HAxp5_ASAP7_75t_R _34521_ (.A(_17774_),
    .B(_17775_),
    .CON(_00687_),
    .SN(_00685_));
 HAxp5_ASAP7_75t_R _34522_ (.A(_17776_),
    .B(_17777_),
    .CON(_02271_),
    .SN(_02272_));
 HAxp5_ASAP7_75t_R _34523_ (.A(_17778_),
    .B(_17779_),
    .CON(_00752_),
    .SN(_00719_));
 HAxp5_ASAP7_75t_R _34524_ (.A(_17780_),
    .B(_17781_),
    .CON(_02273_),
    .SN(_00751_));
 HAxp5_ASAP7_75t_R _34525_ (.A(_16740_),
    .B(_16742_),
    .CON(_00817_),
    .SN(_00784_));
 HAxp5_ASAP7_75t_R _34526_ (.A(_17782_),
    .B(_17783_),
    .CON(_02274_),
    .SN(_02275_));
 HAxp5_ASAP7_75t_R _34527_ (.A(_17784_),
    .B(_17785_),
    .CON(_00883_),
    .SN(_00850_));
 HAxp5_ASAP7_75t_R _34528_ (.A(_17786_),
    .B(_17787_),
    .CON(_02276_),
    .SN(_00882_));
 HAxp5_ASAP7_75t_R _34529_ (.A(_17788_),
    .B(_17789_),
    .CON(_00948_),
    .SN(_00915_));
 HAxp5_ASAP7_75t_R _34530_ (.A(_17790_),
    .B(_17791_),
    .CON(_02277_),
    .SN(_00947_));
 HAxp5_ASAP7_75t_R _34531_ (.A(_16750_),
    .B(_16751_),
    .CON(_01013_),
    .SN(_00980_));
 HAxp5_ASAP7_75t_R _34532_ (.A(_17792_),
    .B(_17793_),
    .CON(_02278_),
    .SN(_01012_));
 HAxp5_ASAP7_75t_R _34533_ (.A(_17794_),
    .B(_17795_),
    .CON(_01079_),
    .SN(_01046_));
 HAxp5_ASAP7_75t_R _34534_ (.A(_17796_),
    .B(_17797_),
    .CON(_02279_),
    .SN(_01078_));
 HAxp5_ASAP7_75t_R _34535_ (.A(_16756_),
    .B(_16757_),
    .CON(_01144_),
    .SN(_01111_));
 HAxp5_ASAP7_75t_R _34536_ (.A(_17798_),
    .B(_17799_),
    .CON(_02280_),
    .SN(_01143_));
 HAxp5_ASAP7_75t_R _34537_ (.A(_16758_),
    .B(_16760_),
    .CON(_01210_),
    .SN(_01177_));
 HAxp5_ASAP7_75t_R _34538_ (.A(_17800_),
    .B(_17801_),
    .CON(_02281_),
    .SN(_01209_));
 HAxp5_ASAP7_75t_R _34539_ (.A(_16761_),
    .B(_16762_),
    .CON(_01276_),
    .SN(_01243_));
 HAxp5_ASAP7_75t_R _34540_ (.A(_17802_),
    .B(_17803_),
    .CON(_01309_),
    .SN(_01275_));
 HAxp5_ASAP7_75t_R _34541_ (.A(_17804_),
    .B(_17805_),
    .CON(_02282_),
    .SN(_01310_));
 HAxp5_ASAP7_75t_R _34542_ (.A(_17806_),
    .B(_17807_),
    .CON(_00160_),
    .SN(_17808_));
 HAxp5_ASAP7_75t_R _34543_ (.A(_17809_),
    .B(_17810_),
    .CON(_02283_),
    .SN(_02284_));
 HAxp5_ASAP7_75t_R _34544_ (.A(_17811_),
    .B(\cs_registers_i.priv_lvl_q[0] ),
    .CON(_02285_),
    .SN(_01313_));
 HAxp5_ASAP7_75t_R _34545_ (.A(_17812_),
    .B(_14713_),
    .CON(_02286_),
    .SN(_02287_));
 HAxp5_ASAP7_75t_R _34546_ (.A(_17812_),
    .B(_14714_),
    .CON(_02288_),
    .SN(_17815_));
 HAxp5_ASAP7_75t_R _34547_ (.A(_17816_),
    .B(_14713_),
    .CON(_02289_),
    .SN(_17817_));
 HAxp5_ASAP7_75t_R _34548_ (.A(_17818_),
    .B(_17819_),
    .CON(_01321_),
    .SN(_02290_));
 HAxp5_ASAP7_75t_R _34549_ (.A(_17818_),
    .B(_17819_),
    .CON(_02291_),
    .SN(_17820_));
 HAxp5_ASAP7_75t_R _34550_ (.A(_17818_),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_01326_),
    .SN(_17822_));
 HAxp5_ASAP7_75t_R _34551_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_17819_),
    .CON(_01319_),
    .SN(_17823_));
 HAxp5_ASAP7_75t_R _34552_ (.A(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\ex_block_i.genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .CON(_01320_),
    .SN(_17824_));
 HAxp5_ASAP7_75t_R _34553_ (.A(_17825_),
    .B(_17821_),
    .CON(_02292_),
    .SN(_02293_));
 HAxp5_ASAP7_75t_R _34554_ (.A(_17826_),
    .B(_17827_),
    .CON(_02294_),
    .SN(_01356_));
 HAxp5_ASAP7_75t_R _34555_ (.A(_17829_),
    .B(_17830_),
    .CON(_02295_),
    .SN(_01358_));
 HAxp5_ASAP7_75t_R _34556_ (.A(_17833_),
    .B(_17832_),
    .CON(_02296_),
    .SN(_01359_));
 HAxp5_ASAP7_75t_R _34557_ (.A(_17835_),
    .B(_17828_),
    .CON(_02297_),
    .SN(_01360_));
 HAxp5_ASAP7_75t_R _34558_ (.A(_17837_),
    .B(_17831_),
    .CON(_02298_),
    .SN(_01361_));
 HAxp5_ASAP7_75t_R _34559_ (.A(_17840_),
    .B(_17839_),
    .CON(_02299_),
    .SN(_01362_));
 HAxp5_ASAP7_75t_R _34560_ (.A(_17842_),
    .B(_17834_),
    .CON(_16771_),
    .SN(_01363_));
 HAxp5_ASAP7_75t_R _34561_ (.A(_17843_),
    .B(_17836_),
    .CON(_16772_),
    .SN(_01364_));
 HAxp5_ASAP7_75t_R _34562_ (.A(_17844_),
    .B(_17845_),
    .CON(_02300_),
    .SN(_01365_));
 HAxp5_ASAP7_75t_R _34563_ (.A(_17847_),
    .B(_17848_),
    .CON(_02301_),
    .SN(_01366_));
 HAxp5_ASAP7_75t_R _34564_ (.A(_17850_),
    .B(_17838_),
    .CON(_02302_),
    .SN(_01367_));
 HAxp5_ASAP7_75t_R _34565_ (.A(_17846_),
    .B(_17852_),
    .CON(_02303_),
    .SN(_01368_));
 HAxp5_ASAP7_75t_R _34566_ (.A(_17854_),
    .B(_17841_),
    .CON(_16783_),
    .SN(_16770_));
 HAxp5_ASAP7_75t_R _34567_ (.A(_17856_),
    .B(_17857_),
    .CON(_02304_),
    .SN(_01369_));
 HAxp5_ASAP7_75t_R _34568_ (.A(_17859_),
    .B(_17858_),
    .CON(_02305_),
    .SN(_01370_));
 HAxp5_ASAP7_75t_R _34569_ (.A(_17860_),
    .B(_17861_),
    .CON(_02306_),
    .SN(_01371_));
 HAxp5_ASAP7_75t_R _34570_ (.A(_17863_),
    .B(_17849_),
    .CON(_02307_),
    .SN(_01372_));
 HAxp5_ASAP7_75t_R _34571_ (.A(_17865_),
    .B(_17851_),
    .CON(_02308_),
    .SN(_01373_));
 HAxp5_ASAP7_75t_R _34572_ (.A(_16781_),
    .B(_17853_),
    .CON(_02309_),
    .SN(_16782_));
 HAxp5_ASAP7_75t_R _34573_ (.A(_17867_),
    .B(_17855_),
    .CON(_01386_),
    .SN(_01375_));
 HAxp5_ASAP7_75t_R _34574_ (.A(_17869_),
    .B(_16787_),
    .CON(_02310_),
    .SN(_01378_));
 HAxp5_ASAP7_75t_R _34575_ (.A(_16796_),
    .B(_17862_),
    .CON(_02311_),
    .SN(_01380_));
 HAxp5_ASAP7_75t_R _34576_ (.A(_17871_),
    .B(_17864_),
    .CON(_02312_),
    .SN(_01381_));
 HAxp5_ASAP7_75t_R _34577_ (.A(_16804_),
    .B(_17866_),
    .CON(_02313_),
    .SN(_01385_));
 HAxp5_ASAP7_75t_R _34578_ (.A(_17872_),
    .B(_16808_),
    .CON(_02314_),
    .SN(_01389_));
 HAxp5_ASAP7_75t_R _34579_ (.A(_17875_),
    .B(_17874_),
    .CON(_02315_),
    .SN(_01390_));
 HAxp5_ASAP7_75t_R _34580_ (.A(_17878_),
    .B(_16795_),
    .CON(_02316_),
    .SN(_01392_));
 HAxp5_ASAP7_75t_R _34581_ (.A(_17880_),
    .B(_17870_),
    .CON(_02317_),
    .SN(_01393_));
 HAxp5_ASAP7_75t_R _34582_ (.A(_16822_),
    .B(_16803_),
    .CON(_01411_),
    .SN(_01398_));
 HAxp5_ASAP7_75t_R _34583_ (.A(_17881_),
    .B(_17882_),
    .CON(_02318_),
    .SN(_01399_));
 HAxp5_ASAP7_75t_R _34584_ (.A(_17883_),
    .B(_16827_),
    .CON(_02319_),
    .SN(_01401_));
 HAxp5_ASAP7_75t_R _34585_ (.A(_17885_),
    .B(_17873_),
    .CON(_16860_),
    .SN(_01402_));
 HAxp5_ASAP7_75t_R _34586_ (.A(_17887_),
    .B(_17886_),
    .CON(_02320_),
    .SN(_01403_));
 HAxp5_ASAP7_75t_R _34587_ (.A(_17890_),
    .B(_17891_),
    .CON(_16862_),
    .SN(_01404_));
 HAxp5_ASAP7_75t_R _34588_ (.A(_17892_),
    .B(_17879_),
    .CON(_02321_),
    .SN(_01405_));
 HAxp5_ASAP7_75t_R _34589_ (.A(_16841_),
    .B(_16821_),
    .CON(_02322_),
    .SN(_01410_));
 HAxp5_ASAP7_75t_R _34590_ (.A(_16853_),
    .B(_17884_),
    .CON(_16887_),
    .SN(_01414_));
 HAxp5_ASAP7_75t_R _34591_ (.A(_17894_),
    .B(_17893_),
    .CON(_02323_),
    .SN(_01415_));
 HAxp5_ASAP7_75t_R _34592_ (.A(_17897_),
    .B(_17898_),
    .CON(_16889_),
    .SN(_16861_));
 HAxp5_ASAP7_75t_R _34593_ (.A(_16870_),
    .B(_16840_),
    .CON(_01427_),
    .SN(_01420_));
 HAxp5_ASAP7_75t_R _34594_ (.A(_17899_),
    .B(_17900_),
    .CON(_02324_),
    .SN(_01421_));
 HAxp5_ASAP7_75t_R _34595_ (.A(_17904_),
    .B(_16852_),
    .CON(_16915_),
    .SN(_01423_));
 HAxp5_ASAP7_75t_R _34596_ (.A(_17901_),
    .B(_17905_),
    .CON(_02325_),
    .SN(_01424_));
 HAxp5_ASAP7_75t_R _34597_ (.A(_17908_),
    .B(_17909_),
    .CON(_16917_),
    .SN(_16888_));
 HAxp5_ASAP7_75t_R _34598_ (.A(_17911_),
    .B(_16869_),
    .CON(_02326_),
    .SN(_01426_));
 HAxp5_ASAP7_75t_R _34599_ (.A(_17912_),
    .B(_17913_),
    .CON(_02327_),
    .SN(_01428_));
 HAxp5_ASAP7_75t_R _34600_ (.A(_17916_),
    .B(_17915_),
    .CON(_02328_),
    .SN(_01429_));
 HAxp5_ASAP7_75t_R _34601_ (.A(_17919_),
    .B(_17920_),
    .CON(_16948_),
    .SN(_01430_));
 HAxp5_ASAP7_75t_R _34602_ (.A(_17923_),
    .B(_17924_),
    .CON(_16950_),
    .SN(_16916_));
 HAxp5_ASAP7_75t_R _34603_ (.A(_16923_),
    .B(net2251),
    .CON(_01437_),
    .SN(_01432_));
 HAxp5_ASAP7_75t_R _34604_ (.A(_17926_),
    .B(_17914_),
    .CON(_16972_),
    .SN(_01433_));
 HAxp5_ASAP7_75t_R _34605_ (.A(_17928_),
    .B(_17927_),
    .CON(_02329_),
    .SN(_01434_));
 HAxp5_ASAP7_75t_R _34606_ (.A(_17931_),
    .B(_17932_),
    .CON(_16982_),
    .SN(_01435_));
 HAxp5_ASAP7_75t_R _34607_ (.A(_17935_),
    .B(_17936_),
    .CON(_16984_),
    .SN(_16949_));
 HAxp5_ASAP7_75t_R _34608_ (.A(_17940_),
    .B(_17941_),
    .CON(_02330_),
    .SN(_01436_));
 HAxp5_ASAP7_75t_R _34609_ (.A(_17942_),
    .B(_17943_),
    .CON(_02331_),
    .SN(_01438_));
 HAxp5_ASAP7_75t_R _34610_ (.A(_17945_),
    .B(_17946_),
    .CON(_17013_),
    .SN(_01439_));
 HAxp5_ASAP7_75t_R _34611_ (.A(_17944_),
    .B(_17947_),
    .CON(_02332_),
    .SN(_01440_));
 HAxp5_ASAP7_75t_R _34612_ (.A(_17954_),
    .B(_17955_),
    .CON(_02333_),
    .SN(_16983_));
 HAxp5_ASAP7_75t_R _34613_ (.A(_16991_),
    .B(_16993_),
    .CON(_00016_),
    .SN(_00009_));
 HAxp5_ASAP7_75t_R _34614_ (.A(_17960_),
    .B(_17961_),
    .CON(_17039_),
    .SN(_00010_));
 HAxp5_ASAP7_75t_R _34615_ (.A(_17962_),
    .B(_17963_),
    .CON(_02334_),
    .SN(_00011_));
 HAxp5_ASAP7_75t_R _34616_ (.A(_17964_),
    .B(_17965_),
    .CON(_17055_),
    .SN(_00012_));
 HAxp5_ASAP7_75t_R _34617_ (.A(_17972_),
    .B(_17973_),
    .CON(_02335_),
    .SN(_00014_));
 HAxp5_ASAP7_75t_R _34618_ (.A(_17977_),
    .B(_17978_),
    .CON(_02336_),
    .SN(_00015_));
 HAxp5_ASAP7_75t_R _34619_ (.A(_17979_),
    .B(_17980_),
    .CON(_02337_),
    .SN(_00017_));
 HAxp5_ASAP7_75t_R _34620_ (.A(_17991_),
    .B(_17992_),
    .CON(_02338_),
    .SN(_00018_));
 HAxp5_ASAP7_75t_R _34621_ (.A(_17076_),
    .B(_17077_),
    .CON(_00025_),
    .SN(_00019_));
 HAxp5_ASAP7_75t_R _34622_ (.A(_17995_),
    .B(_17996_),
    .CON(_02339_),
    .SN(_00020_));
 HAxp5_ASAP7_75t_R _34623_ (.A(_17997_),
    .B(_17081_),
    .CON(_02340_),
    .SN(_00022_));
 HAxp5_ASAP7_75t_R _34624_ (.A(_18011_),
    .B(_18012_),
    .CON(_02341_),
    .SN(_00023_));
 HAxp5_ASAP7_75t_R _34625_ (.A(_18015_),
    .B(_18016_),
    .CON(_02342_),
    .SN(_00024_));
 HAxp5_ASAP7_75t_R _34626_ (.A(net2232),
    .B(_18032_),
    .CON(_00032_),
    .SN(_00029_));
 HAxp5_ASAP7_75t_R _34627_ (.A(_18050_),
    .B(_18051_),
    .CON(_02343_),
    .SN(_17219_));
 HAxp5_ASAP7_75t_R _34628_ (.A(_18056_),
    .B(_18057_),
    .CON(_02344_),
    .SN(_00031_));
 HAxp5_ASAP7_75t_R _34629_ (.A(_18077_),
    .B(_18078_),
    .CON(_02345_),
    .SN(_00035_));
 HAxp5_ASAP7_75t_R _34630_ (.A(net2161),
    .B(_17275_),
    .CON(_00039_),
    .SN(_00036_));
 HAxp5_ASAP7_75t_R _34631_ (.A(_18101_),
    .B(_18102_),
    .CON(_02346_),
    .SN(_00037_));
 HAxp5_ASAP7_75t_R _34632_ (.A(_18105_),
    .B(_18106_),
    .CON(_02347_),
    .SN(_00038_));
 HAxp5_ASAP7_75t_R _34633_ (.A(_18126_),
    .B(_18127_),
    .CON(_02348_),
    .SN(_00040_));
 HAxp5_ASAP7_75t_R _34634_ (.A(_17362_),
    .B(_17363_),
    .CON(_00045_),
    .SN(_00041_));
 HAxp5_ASAP7_75t_R _34635_ (.A(_17405_),
    .B(_18148_),
    .CON(_02349_),
    .SN(_00043_));
 HAxp5_ASAP7_75t_R _34636_ (.A(_18151_),
    .B(_18152_),
    .CON(_02350_),
    .SN(_00044_));
 HAxp5_ASAP7_75t_R _34637_ (.A(_17444_),
    .B(_17404_),
    .CON(_02351_),
    .SN(_00048_));
 HAxp5_ASAP7_75t_R _34638_ (.A(_17453_),
    .B(_17454_),
    .CON(_00053_),
    .SN(_00049_));
 HAxp5_ASAP7_75t_R _34639_ (.A(_17444_),
    .B(_17443_),
    .CON(_02352_),
    .SN(_00051_));
 HAxp5_ASAP7_75t_R _34640_ (.A(_18192_),
    .B(_18193_),
    .CON(_02353_),
    .SN(_00052_));
 HAxp5_ASAP7_75t_R _34641_ (.A(_17531_),
    .B(_17532_),
    .CON(_00056_),
    .SN(_00054_));
 HAxp5_ASAP7_75t_R _34642_ (.A(_18228_),
    .B(_18229_),
    .CON(_02354_),
    .SN(_00055_));
 HAxp5_ASAP7_75t_R _34643_ (.A(_17597_),
    .B(_17598_),
    .CON(_00059_),
    .SN(_00057_));
 HAxp5_ASAP7_75t_R _34644_ (.A(_18263_),
    .B(_18264_),
    .CON(_02355_),
    .SN(_00058_));
 HAxp5_ASAP7_75t_R _34645_ (.A(_17655_),
    .B(_17656_),
    .CON(_00062_),
    .SN(_00060_));
 HAxp5_ASAP7_75t_R _34646_ (.A(_18295_),
    .B(_18296_),
    .CON(_02356_),
    .SN(_00061_));
 HAxp5_ASAP7_75t_R _34647_ (.A(_17707_),
    .B(_17708_),
    .CON(_00065_),
    .SN(_00063_));
 HAxp5_ASAP7_75t_R _34648_ (.A(_18313_),
    .B(_18314_),
    .CON(_00067_),
    .SN(_00064_));
 HAxp5_ASAP7_75t_R _34649_ (.A(net304),
    .B(_13523_),
    .CON(_02357_),
    .SN(_00072_));
 HAxp5_ASAP7_75t_R _34650_ (.A(_14180_),
    .B(_18324_),
    .CON(_02358_),
    .SN(_00073_));
 HAxp5_ASAP7_75t_R _34651_ (.A(_13893_),
    .B(_18326_),
    .CON(_00074_),
    .SN(_02359_));
 HAxp5_ASAP7_75t_R _34652_ (.A(_13894_),
    .B(_13999_),
    .CON(_02360_),
    .SN(_18329_));
 HAxp5_ASAP7_75t_R _34653_ (.A(_18330_),
    .B(_13525_),
    .CON(_00076_),
    .SN(_00075_));
 HAxp5_ASAP7_75t_R _34654_ (.A(_18332_),
    .B(_13523_),
    .CON(_02361_),
    .SN(_18333_));
 HAxp5_ASAP7_75t_R _34655_ (.A(_14179_),
    .B(_18335_),
    .CON(_00078_),
    .SN(_00077_));
 HAxp5_ASAP7_75t_R _34656_ (.A(_14180_),
    .B(_18336_),
    .CON(_02362_),
    .SN(_18337_));
 HAxp5_ASAP7_75t_R _34657_ (.A(_14238_),
    .B(_18339_),
    .CON(_02363_),
    .SN(_00079_));
 HAxp5_ASAP7_75t_R _34658_ (.A(_14239_),
    .B(_18341_),
    .CON(_00080_),
    .SN(_18342_));
 HAxp5_ASAP7_75t_R _34659_ (.A(_14296_),
    .B(_18344_),
    .CON(_02364_),
    .SN(_00082_));
 HAxp5_ASAP7_75t_R _34660_ (.A(_14297_),
    .B(_18346_),
    .CON(_00083_),
    .SN(_18347_));
 HAxp5_ASAP7_75t_R _34661_ (.A(_14358_),
    .B(_15115_),
    .CON(_00086_),
    .SN(_00085_));
 HAxp5_ASAP7_75t_R _34662_ (.A(_14359_),
    .B(_18351_),
    .CON(_02365_),
    .SN(_18352_));
 HAxp5_ASAP7_75t_R _34663_ (.A(_18353_),
    .B(_15172_),
    .CON(_00089_),
    .SN(_00088_));
 HAxp5_ASAP7_75t_R _34664_ (.A(_18355_),
    .B(_18356_),
    .CON(_02366_),
    .SN(_18357_));
 HAxp5_ASAP7_75t_R _34665_ (.A(_14481_),
    .B(_15226_),
    .CON(_00092_),
    .SN(_00091_));
 HAxp5_ASAP7_75t_R _34666_ (.A(_18360_),
    .B(_18361_),
    .CON(_02367_),
    .SN(_18362_));
 HAxp5_ASAP7_75t_R _34667_ (.A(_18363_),
    .B(_15280_),
    .CON(_00094_),
    .SN(_00093_));
 HAxp5_ASAP7_75t_R _34668_ (.A(_18365_),
    .B(_18366_),
    .CON(_02368_),
    .SN(_18367_));
 HAxp5_ASAP7_75t_R _34669_ (.A(_14599_),
    .B(_15337_),
    .CON(_00097_),
    .SN(_00096_));
 HAxp5_ASAP7_75t_R _34670_ (.A(_18370_),
    .B(_18371_),
    .CON(_02369_),
    .SN(_18372_));
 HAxp5_ASAP7_75t_R _34671_ (.A(_14653_),
    .B(_15401_),
    .CON(_00100_),
    .SN(_00099_));
 HAxp5_ASAP7_75t_R _34672_ (.A(_18375_),
    .B(_18376_),
    .CON(_02370_),
    .SN(_18377_));
 HAxp5_ASAP7_75t_R _34673_ (.A(_14710_),
    .B(_18379_),
    .CON(_02371_),
    .SN(_00102_));
 HAxp5_ASAP7_75t_R _34674_ (.A(_18380_),
    .B(_18381_),
    .CON(_00103_),
    .SN(_18382_));
 HAxp5_ASAP7_75t_R _34675_ (.A(_18383_),
    .B(_18384_),
    .CON(_00105_),
    .SN(_00104_));
 HAxp5_ASAP7_75t_R _34676_ (.A(_18385_),
    .B(_18386_),
    .CON(_02372_),
    .SN(_18387_));
 HAxp5_ASAP7_75t_R _34677_ (.A(_18388_),
    .B(_18389_),
    .CON(_00107_),
    .SN(_00106_));
 HAxp5_ASAP7_75t_R _34678_ (.A(_18390_),
    .B(_18391_),
    .CON(_02373_),
    .SN(_18392_));
 HAxp5_ASAP7_75t_R _34679_ (.A(_18393_),
    .B(_18394_),
    .CON(_02374_),
    .SN(_00109_));
 HAxp5_ASAP7_75t_R _34680_ (.A(_18395_),
    .B(_18396_),
    .CON(_00110_),
    .SN(_18397_));
 HAxp5_ASAP7_75t_R _34681_ (.A(_15887_),
    .B(_18399_),
    .CON(_00113_),
    .SN(_00112_));
 HAxp5_ASAP7_75t_R _34682_ (.A(_18400_),
    .B(_15841_),
    .CON(_02375_),
    .SN(_18402_));
 HAxp5_ASAP7_75t_R _34683_ (.A(_18403_),
    .B(_18404_),
    .CON(_02376_),
    .SN(_00115_));
 HAxp5_ASAP7_75t_R _34684_ (.A(_18405_),
    .B(_16020_),
    .CON(_00116_),
    .SN(_18407_));
 HAxp5_ASAP7_75t_R _34685_ (.A(_18408_),
    .B(_18409_),
    .CON(_02377_),
    .SN(_00118_));
 HAxp5_ASAP7_75t_R _34686_ (.A(_18410_),
    .B(_16145_),
    .CON(_00119_),
    .SN(_18412_));
 HAxp5_ASAP7_75t_R _34687_ (.A(_18413_),
    .B(_16262_),
    .CON(_02378_),
    .SN(_00121_));
 HAxp5_ASAP7_75t_R _34688_ (.A(_18415_),
    .B(_18416_),
    .CON(_00122_),
    .SN(_18417_));
 HAxp5_ASAP7_75t_R _34689_ (.A(_18418_),
    .B(_18419_),
    .CON(_00125_),
    .SN(_00124_));
 HAxp5_ASAP7_75t_R _34690_ (.A(_16386_),
    .B(_18421_),
    .CON(_02379_),
    .SN(_18422_));
 HAxp5_ASAP7_75t_R _34691_ (.A(_18423_),
    .B(_18424_),
    .CON(_02380_),
    .SN(_00127_));
 HAxp5_ASAP7_75t_R _34692_ (.A(_18425_),
    .B(_18426_),
    .CON(_00128_),
    .SN(_18427_));
 HAxp5_ASAP7_75t_R _34693_ (.A(_16571_),
    .B(_18429_),
    .CON(_02381_),
    .SN(_00130_));
 HAxp5_ASAP7_75t_R _34694_ (.A(_18430_),
    .B(_16620_),
    .CON(_00131_),
    .SN(_18432_));
 HAxp5_ASAP7_75t_R _34695_ (.A(_04516_),
    .B(_18434_),
    .CON(_00134_),
    .SN(_00133_));
 HAxp5_ASAP7_75t_R _34696_ (.A(_18435_),
    .B(_18436_),
    .CON(_02382_),
    .SN(_18437_));
 HAxp5_ASAP7_75t_R _34697_ (.A(_04632_),
    .B(_18439_),
    .CON(_00137_),
    .SN(_00136_));
 HAxp5_ASAP7_75t_R _34698_ (.A(_18440_),
    .B(_18441_),
    .CON(_02383_),
    .SN(_18442_));
 HAxp5_ASAP7_75t_R _34699_ (.A(_04700_),
    .B(_18444_),
    .CON(_02384_),
    .SN(_00139_));
 HAxp5_ASAP7_75t_R _34700_ (.A(_18445_),
    .B(_18446_),
    .CON(_00140_),
    .SN(_18447_));
 HAxp5_ASAP7_75t_R _34701_ (.A(_04810_),
    .B(_18449_),
    .CON(_02385_),
    .SN(_00142_));
 HAxp5_ASAP7_75t_R _34702_ (.A(_18450_),
    .B(_04857_),
    .CON(_00143_),
    .SN(_18452_));
 HAxp5_ASAP7_75t_R _34703_ (.A(_04967_),
    .B(_04919_),
    .CON(_00146_),
    .SN(_00145_));
 HAxp5_ASAP7_75t_R _34704_ (.A(_18455_),
    .B(_18456_),
    .CON(_02386_),
    .SN(_18457_));
 HAxp5_ASAP7_75t_R _34705_ (.A(_05077_),
    .B(_18459_),
    .CON(_00149_),
    .SN(_00148_));
 HAxp5_ASAP7_75t_R _34706_ (.A(_18460_),
    .B(_05030_),
    .CON(_02387_),
    .SN(_18462_));
 HAxp5_ASAP7_75t_R _34707_ (.A(_05138_),
    .B(_05184_),
    .CON(_02388_),
    .SN(_00151_));
 HAxp5_ASAP7_75t_R _34708_ (.A(_18465_),
    .B(_18466_),
    .CON(_00152_),
    .SN(_18467_));
 HAxp5_ASAP7_75t_R _34709_ (.A(_05247_),
    .B(_18469_),
    .CON(_02389_),
    .SN(_00154_));
 HAxp5_ASAP7_75t_R _34710_ (.A(_18470_),
    .B(_18471_),
    .CON(_00155_),
    .SN(_18472_));
 HAxp5_ASAP7_75t_R _34711_ (.A(_05357_),
    .B(_18474_),
    .CON(_02390_),
    .SN(_00157_));
 HAxp5_ASAP7_75t_R _34712_ (.A(_18475_),
    .B(_18476_),
    .CON(_00158_),
    .SN(_18477_));
 HAxp5_ASAP7_75t_R _34713_ (.A(\cs_registers_i.mhpmcounter[2][0] ),
    .B(\cs_registers_i.mhpmcounter[2][1] ),
    .CON(_02391_),
    .SN(_02392_));
 HAxp5_ASAP7_75t_R _34714_ (.A(\cs_registers_i.mhpmcounter[2][2] ),
    .B(_18478_),
    .CON(_02393_),
    .SN(_02394_));
 HAxp5_ASAP7_75t_R _34715_ (.A(\cs_registers_i.mhpmcounter[2][4] ),
    .B(_18479_),
    .CON(_02395_),
    .SN(_02396_));
 HAxp5_ASAP7_75t_R _34716_ (.A(\cs_registers_i.mhpmcounter[2][6] ),
    .B(_18480_),
    .CON(_02397_),
    .SN(_02398_));
 HAxp5_ASAP7_75t_R _34717_ (.A(\cs_registers_i.mhpmcounter[2][8] ),
    .B(_18481_),
    .CON(_02399_),
    .SN(_02400_));
 HAxp5_ASAP7_75t_R _34718_ (.A(\cs_registers_i.mhpmcounter[2][10] ),
    .B(_18482_),
    .CON(_02401_),
    .SN(_02402_));
 HAxp5_ASAP7_75t_R _34719_ (.A(\cs_registers_i.mhpmcounter[2][12] ),
    .B(_18483_),
    .CON(_02403_),
    .SN(_02404_));
 HAxp5_ASAP7_75t_R _34720_ (.A(\cs_registers_i.mhpmcounter[2][14] ),
    .B(_18484_),
    .CON(_02405_),
    .SN(_02406_));
 HAxp5_ASAP7_75t_R _34721_ (.A(\cs_registers_i.mhpmcounter[2][16] ),
    .B(_18485_),
    .CON(_02407_),
    .SN(_02408_));
 HAxp5_ASAP7_75t_R _34722_ (.A(\cs_registers_i.mhpmcounter[2][18] ),
    .B(_18486_),
    .CON(_02409_),
    .SN(_02410_));
 HAxp5_ASAP7_75t_R _34723_ (.A(\cs_registers_i.mhpmcounter[2][20] ),
    .B(_18487_),
    .CON(_02411_),
    .SN(_02412_));
 HAxp5_ASAP7_75t_R _34724_ (.A(\cs_registers_i.mhpmcounter[2][22] ),
    .B(_18488_),
    .CON(_02413_),
    .SN(_02414_));
 HAxp5_ASAP7_75t_R _34725_ (.A(\cs_registers_i.mhpmcounter[2][24] ),
    .B(_18489_),
    .CON(_02415_),
    .SN(_02416_));
 HAxp5_ASAP7_75t_R _34726_ (.A(\cs_registers_i.mhpmcounter[2][26] ),
    .B(_18490_),
    .CON(_02417_),
    .SN(_02418_));
 HAxp5_ASAP7_75t_R _34727_ (.A(\cs_registers_i.mhpmcounter[2][28] ),
    .B(_18491_),
    .CON(_02419_),
    .SN(_02420_));
 HAxp5_ASAP7_75t_R _34728_ (.A(\cs_registers_i.mhpmcounter[2][30] ),
    .B(_18492_),
    .CON(_02421_),
    .SN(_02422_));
 HAxp5_ASAP7_75t_R _34729_ (.A(\cs_registers_i.mhpmcounter[2][32] ),
    .B(_18493_),
    .CON(_02423_),
    .SN(_02424_));
 HAxp5_ASAP7_75t_R _34730_ (.A(\cs_registers_i.mhpmcounter[2][34] ),
    .B(_18494_),
    .CON(_02425_),
    .SN(_02426_));
 HAxp5_ASAP7_75t_R _34731_ (.A(\cs_registers_i.mhpmcounter[2][36] ),
    .B(_18495_),
    .CON(_02427_),
    .SN(_02428_));
 HAxp5_ASAP7_75t_R _34732_ (.A(\cs_registers_i.mhpmcounter[2][38] ),
    .B(_18496_),
    .CON(_02429_),
    .SN(_02430_));
 HAxp5_ASAP7_75t_R _34733_ (.A(\cs_registers_i.mhpmcounter[2][40] ),
    .B(_18497_),
    .CON(_02431_),
    .SN(_02432_));
 HAxp5_ASAP7_75t_R _34734_ (.A(\cs_registers_i.mhpmcounter[2][42] ),
    .B(_18498_),
    .CON(_02433_),
    .SN(_02434_));
 HAxp5_ASAP7_75t_R _34735_ (.A(\cs_registers_i.mhpmcounter[2][44] ),
    .B(_18499_),
    .CON(_02435_),
    .SN(_02436_));
 HAxp5_ASAP7_75t_R _34736_ (.A(\cs_registers_i.mhpmcounter[2][46] ),
    .B(_18500_),
    .CON(_02437_),
    .SN(_02438_));
 HAxp5_ASAP7_75t_R _34737_ (.A(\cs_registers_i.mhpmcounter[2][48] ),
    .B(_18501_),
    .CON(_02439_),
    .SN(_02440_));
 HAxp5_ASAP7_75t_R _34738_ (.A(\cs_registers_i.mhpmcounter[2][50] ),
    .B(_18502_),
    .CON(_02441_),
    .SN(_02442_));
 HAxp5_ASAP7_75t_R _34739_ (.A(\cs_registers_i.mhpmcounter[2][52] ),
    .B(_18503_),
    .CON(_02443_),
    .SN(_02444_));
 HAxp5_ASAP7_75t_R _34740_ (.A(\cs_registers_i.mhpmcounter[2][54] ),
    .B(_18504_),
    .CON(_02445_),
    .SN(_02446_));
 HAxp5_ASAP7_75t_R _34741_ (.A(\cs_registers_i.mhpmcounter[2][56] ),
    .B(_18505_),
    .CON(_02447_),
    .SN(_02448_));
 HAxp5_ASAP7_75t_R _34742_ (.A(\cs_registers_i.mhpmcounter[2][58] ),
    .B(_18506_),
    .CON(_02449_),
    .SN(_02450_));
 HAxp5_ASAP7_75t_R _34743_ (.A(\cs_registers_i.mhpmcounter[2][60] ),
    .B(_18507_),
    .CON(_02451_),
    .SN(_02452_));
 HAxp5_ASAP7_75t_R _34744_ (.A(\cs_registers_i.mhpmcounter[2][62] ),
    .B(_18508_),
    .CON(_02453_),
    .SN(_02454_));
 HAxp5_ASAP7_75t_R _34745_ (.A(\cs_registers_i.mcycle_counter_i.counter[0] ),
    .B(\cs_registers_i.mcycle_counter_i.counter[1] ),
    .CON(_02455_),
    .SN(_02456_));
 HAxp5_ASAP7_75t_R _34746_ (.A(\cs_registers_i.mcycle_counter_i.counter[2] ),
    .B(_18509_),
    .CON(_02457_),
    .SN(_02458_));
 HAxp5_ASAP7_75t_R _34747_ (.A(\cs_registers_i.mcycle_counter_i.counter[4] ),
    .B(_18510_),
    .CON(_02459_),
    .SN(_02460_));
 HAxp5_ASAP7_75t_R _34748_ (.A(\cs_registers_i.mcycle_counter_i.counter[6] ),
    .B(_18511_),
    .CON(_02461_),
    .SN(_02462_));
 HAxp5_ASAP7_75t_R _34749_ (.A(\cs_registers_i.mcycle_counter_i.counter[8] ),
    .B(_18512_),
    .CON(_02463_),
    .SN(_02464_));
 HAxp5_ASAP7_75t_R _34750_ (.A(\cs_registers_i.mcycle_counter_i.counter[10] ),
    .B(_18513_),
    .CON(_02465_),
    .SN(_02466_));
 HAxp5_ASAP7_75t_R _34751_ (.A(\cs_registers_i.mcycle_counter_i.counter[12] ),
    .B(_18514_),
    .CON(_02467_),
    .SN(_02468_));
 HAxp5_ASAP7_75t_R _34752_ (.A(\cs_registers_i.mcycle_counter_i.counter[14] ),
    .B(_18515_),
    .CON(_02469_),
    .SN(_02470_));
 HAxp5_ASAP7_75t_R _34753_ (.A(\cs_registers_i.mcycle_counter_i.counter[16] ),
    .B(_18516_),
    .CON(_02471_),
    .SN(_02472_));
 HAxp5_ASAP7_75t_R _34754_ (.A(\cs_registers_i.mcycle_counter_i.counter[18] ),
    .B(_18517_),
    .CON(_02473_),
    .SN(_02474_));
 HAxp5_ASAP7_75t_R _34755_ (.A(\cs_registers_i.mcycle_counter_i.counter[20] ),
    .B(_18518_),
    .CON(_02475_),
    .SN(_02476_));
 HAxp5_ASAP7_75t_R _34756_ (.A(\cs_registers_i.mcycle_counter_i.counter[22] ),
    .B(_18519_),
    .CON(_02477_),
    .SN(_02478_));
 HAxp5_ASAP7_75t_R _34757_ (.A(\cs_registers_i.mcycle_counter_i.counter[24] ),
    .B(_18520_),
    .CON(_02479_),
    .SN(_02480_));
 HAxp5_ASAP7_75t_R _34758_ (.A(\cs_registers_i.mcycle_counter_i.counter[26] ),
    .B(_18521_),
    .CON(_02481_),
    .SN(_02482_));
 HAxp5_ASAP7_75t_R _34759_ (.A(\cs_registers_i.mcycle_counter_i.counter[28] ),
    .B(_18522_),
    .CON(_02483_),
    .SN(_02484_));
 HAxp5_ASAP7_75t_R _34760_ (.A(\cs_registers_i.mcycle_counter_i.counter[30] ),
    .B(_18523_),
    .CON(_02485_),
    .SN(_02486_));
 HAxp5_ASAP7_75t_R _34761_ (.A(\cs_registers_i.mcycle_counter_i.counter[32] ),
    .B(_18524_),
    .CON(_02487_),
    .SN(_02488_));
 HAxp5_ASAP7_75t_R _34762_ (.A(\cs_registers_i.mcycle_counter_i.counter[34] ),
    .B(_18525_),
    .CON(_02489_),
    .SN(_02490_));
 HAxp5_ASAP7_75t_R _34763_ (.A(\cs_registers_i.mcycle_counter_i.counter[36] ),
    .B(_18526_),
    .CON(_02491_),
    .SN(_02492_));
 HAxp5_ASAP7_75t_R _34764_ (.A(\cs_registers_i.mcycle_counter_i.counter[38] ),
    .B(_18527_),
    .CON(_02493_),
    .SN(_02494_));
 HAxp5_ASAP7_75t_R _34765_ (.A(\cs_registers_i.mcycle_counter_i.counter[40] ),
    .B(_18528_),
    .CON(_02495_),
    .SN(_02496_));
 HAxp5_ASAP7_75t_R _34766_ (.A(\cs_registers_i.mcycle_counter_i.counter[42] ),
    .B(_18529_),
    .CON(_02497_),
    .SN(_02498_));
 HAxp5_ASAP7_75t_R _34767_ (.A(\cs_registers_i.mcycle_counter_i.counter[44] ),
    .B(_18530_),
    .CON(_02499_),
    .SN(_02500_));
 HAxp5_ASAP7_75t_R _34768_ (.A(\cs_registers_i.mcycle_counter_i.counter[46] ),
    .B(_18531_),
    .CON(_02501_),
    .SN(_02502_));
 HAxp5_ASAP7_75t_R _34769_ (.A(\cs_registers_i.mcycle_counter_i.counter[48] ),
    .B(_18532_),
    .CON(_02503_),
    .SN(_02504_));
 HAxp5_ASAP7_75t_R _34770_ (.A(\cs_registers_i.mcycle_counter_i.counter[50] ),
    .B(_18533_),
    .CON(_02505_),
    .SN(_02506_));
 HAxp5_ASAP7_75t_R _34771_ (.A(\cs_registers_i.mcycle_counter_i.counter[52] ),
    .B(_18534_),
    .CON(_02507_),
    .SN(_02508_));
 HAxp5_ASAP7_75t_R _34772_ (.A(\cs_registers_i.mcycle_counter_i.counter[54] ),
    .B(_18535_),
    .CON(_02509_),
    .SN(_02510_));
 HAxp5_ASAP7_75t_R _34773_ (.A(\cs_registers_i.mcycle_counter_i.counter[56] ),
    .B(_18536_),
    .CON(_02511_),
    .SN(_02512_));
 HAxp5_ASAP7_75t_R _34774_ (.A(\cs_registers_i.mcycle_counter_i.counter[58] ),
    .B(_18537_),
    .CON(_02513_),
    .SN(_02514_));
 HAxp5_ASAP7_75t_R _34775_ (.A(\cs_registers_i.mcycle_counter_i.counter[60] ),
    .B(_18538_),
    .CON(_02515_),
    .SN(_02516_));
 HAxp5_ASAP7_75t_R _34776_ (.A(\cs_registers_i.mcycle_counter_i.counter[62] ),
    .B(_18539_),
    .CON(_02517_),
    .SN(_02518_));
 HAxp5_ASAP7_75t_R _34777_ (.A(\cs_registers_i.pc_id_i[1] ),
    .B(\cs_registers_i.pc_id_i[2] ),
    .CON(_02519_),
    .SN(_00167_));
 HAxp5_ASAP7_75t_R _34778_ (.A(\cs_registers_i.pc_id_i[3] ),
    .B(_18540_),
    .CON(_02520_),
    .SN(_00171_));
 HAxp5_ASAP7_75t_R _34779_ (.A(\cs_registers_i.pc_id_i[5] ),
    .B(_18541_),
    .CON(_02521_),
    .SN(_00178_));
 HAxp5_ASAP7_75t_R _34780_ (.A(\cs_registers_i.pc_id_i[7] ),
    .B(_18542_),
    .CON(_02522_),
    .SN(_00183_));
 HAxp5_ASAP7_75t_R _34781_ (.A(\cs_registers_i.pc_id_i[9] ),
    .B(_18543_),
    .CON(_02523_),
    .SN(_00190_));
 HAxp5_ASAP7_75t_R _34782_ (.A(\cs_registers_i.pc_id_i[11] ),
    .B(_18544_),
    .CON(_02524_),
    .SN(_00197_));
 HAxp5_ASAP7_75t_R _34783_ (.A(\cs_registers_i.pc_id_i[13] ),
    .B(_18545_),
    .CON(_02525_),
    .SN(_00202_));
 HAxp5_ASAP7_75t_R _34784_ (.A(\cs_registers_i.pc_id_i[15] ),
    .B(_18546_),
    .CON(_02526_),
    .SN(_00207_));
 HAxp5_ASAP7_75t_R _34785_ (.A(\cs_registers_i.pc_id_i[17] ),
    .B(_18547_),
    .CON(_02527_),
    .SN(_00210_));
 HAxp5_ASAP7_75t_R _34786_ (.A(\cs_registers_i.pc_id_i[19] ),
    .B(_18548_),
    .CON(_02528_),
    .SN(_00213_));
 HAxp5_ASAP7_75t_R _34787_ (.A(\cs_registers_i.pc_id_i[21] ),
    .B(_18549_),
    .CON(_02529_),
    .SN(_00216_));
 HAxp5_ASAP7_75t_R _34788_ (.A(\cs_registers_i.pc_id_i[23] ),
    .B(_18550_),
    .CON(_02530_),
    .SN(_00219_));
 HAxp5_ASAP7_75t_R _34789_ (.A(\cs_registers_i.pc_id_i[25] ),
    .B(_18551_),
    .CON(_02531_),
    .SN(_00222_));
 HAxp5_ASAP7_75t_R _34790_ (.A(\cs_registers_i.pc_id_i[27] ),
    .B(_18552_),
    .CON(_02532_),
    .SN(_00225_));
 HAxp5_ASAP7_75t_R _34791_ (.A(\cs_registers_i.pc_id_i[29] ),
    .B(_18553_),
    .CON(_02533_),
    .SN(_00228_));
 HAxp5_ASAP7_75t_R _34792_ (.A(_18554_),
    .B(net292),
    .CON(_02534_),
    .SN(_02535_));
 HAxp5_ASAP7_75t_R _34793_ (.A(net296),
    .B(_18554_),
    .CON(_00236_),
    .SN(_02536_));
 HAxp5_ASAP7_75t_R _34794_ (.A(_16717_),
    .B(_18554_),
    .CON(_00233_),
    .SN(_18556_));
 HAxp5_ASAP7_75t_R _34795_ (.A(net296),
    .B(net298),
    .CON(_00234_),
    .SN(_00235_));
 HAxp5_ASAP7_75t_R _34796_ (.A(net296),
    .B(net298),
    .CON(_02537_),
    .SN(_18557_));
 HAxp5_ASAP7_75t_R _34797_ (.A(net296),
    .B(_16721_),
    .CON(_00231_),
    .SN(_18558_));
 HAxp5_ASAP7_75t_R _34798_ (.A(_16717_),
    .B(net298),
    .CON(_00232_),
    .SN(_18559_));
 HAxp5_ASAP7_75t_R _34799_ (.A(_16717_),
    .B(_16721_),
    .CON(_18555_),
    .SN(_18560_));
 HAxp5_ASAP7_75t_R _34800_ (.A(_17753_),
    .B(\cs_registers_i.pc_if_i[3] ),
    .CON(_02538_),
    .SN(_02539_));
 HAxp5_ASAP7_75t_R _34801_ (.A(_18561_),
    .B(\cs_registers_i.pc_if_i[5] ),
    .CON(_02540_),
    .SN(_02541_));
 HAxp5_ASAP7_75t_R _34802_ (.A(_18562_),
    .B(\cs_registers_i.pc_if_i[7] ),
    .CON(_02542_),
    .SN(_02543_));
 HAxp5_ASAP7_75t_R _34803_ (.A(_18563_),
    .B(\cs_registers_i.pc_if_i[9] ),
    .CON(_02544_),
    .SN(_02545_));
 HAxp5_ASAP7_75t_R _34804_ (.A(_18564_),
    .B(\cs_registers_i.pc_if_i[11] ),
    .CON(_02546_),
    .SN(_02547_));
 HAxp5_ASAP7_75t_R _34805_ (.A(_18565_),
    .B(\cs_registers_i.pc_if_i[13] ),
    .CON(_02548_),
    .SN(_02549_));
 HAxp5_ASAP7_75t_R _34806_ (.A(_18566_),
    .B(\cs_registers_i.pc_if_i[15] ),
    .CON(_02550_),
    .SN(_02551_));
 HAxp5_ASAP7_75t_R _34807_ (.A(_18567_),
    .B(\cs_registers_i.pc_if_i[17] ),
    .CON(_02552_),
    .SN(_02553_));
 HAxp5_ASAP7_75t_R _34808_ (.A(_18568_),
    .B(\cs_registers_i.pc_if_i[19] ),
    .CON(_02554_),
    .SN(_02555_));
 HAxp5_ASAP7_75t_R _34809_ (.A(_18569_),
    .B(\cs_registers_i.pc_if_i[21] ),
    .CON(_02556_),
    .SN(_02557_));
 HAxp5_ASAP7_75t_R _34810_ (.A(_18570_),
    .B(\cs_registers_i.pc_if_i[23] ),
    .CON(_02558_),
    .SN(_02559_));
 HAxp5_ASAP7_75t_R _34811_ (.A(_18571_),
    .B(\cs_registers_i.pc_if_i[25] ),
    .CON(_02560_),
    .SN(_02561_));
 HAxp5_ASAP7_75t_R _34812_ (.A(_18572_),
    .B(\cs_registers_i.pc_if_i[27] ),
    .CON(_02562_),
    .SN(_02563_));
 HAxp5_ASAP7_75t_R _34813_ (.A(_18573_),
    .B(\cs_registers_i.pc_if_i[29] ),
    .CON(_02564_),
    .SN(_02565_));
 HAxp5_ASAP7_75t_R _34814_ (.A(_18574_),
    .B(_18575_),
    .CON(_02566_),
    .SN(_02567_));
 HAxp5_ASAP7_75t_R _34815_ (.A(_18576_),
    .B(_18577_),
    .CON(_02568_),
    .SN(_02569_));
 HAxp5_ASAP7_75t_R _34816_ (.A(_18578_),
    .B(_18579_),
    .CON(_02570_),
    .SN(_02571_));
 HAxp5_ASAP7_75t_R _34817_ (.A(_18580_),
    .B(_18581_),
    .CON(_02572_),
    .SN(_02573_));
 HAxp5_ASAP7_75t_R _34818_ (.A(_18582_),
    .B(_18583_),
    .CON(_02574_),
    .SN(_02575_));
 HAxp5_ASAP7_75t_R _34819_ (.A(_18584_),
    .B(_18585_),
    .CON(_02576_),
    .SN(_02577_));
 HAxp5_ASAP7_75t_R _34820_ (.A(_18586_),
    .B(_18587_),
    .CON(_02578_),
    .SN(_02579_));
 HAxp5_ASAP7_75t_R _34821_ (.A(_18588_),
    .B(_18589_),
    .CON(_02580_),
    .SN(_02581_));
 HAxp5_ASAP7_75t_R _34822_ (.A(_18590_),
    .B(_18591_),
    .CON(_02582_),
    .SN(_02583_));
 HAxp5_ASAP7_75t_R _34823_ (.A(_18592_),
    .B(_18593_),
    .CON(_02584_),
    .SN(_02585_));
 HAxp5_ASAP7_75t_R _34824_ (.A(_18594_),
    .B(_18595_),
    .CON(_02586_),
    .SN(_02587_));
 HAxp5_ASAP7_75t_R _34825_ (.A(_18596_),
    .B(_18597_),
    .CON(_02588_),
    .SN(_02589_));
 HAxp5_ASAP7_75t_R _34826_ (.A(_18598_),
    .B(_18599_),
    .CON(_02590_),
    .SN(_02591_));
 HAxp5_ASAP7_75t_R _34827_ (.A(_18600_),
    .B(_18601_),
    .CON(_02592_),
    .SN(_02593_));
 HAxp5_ASAP7_75t_R _34828_ (.A(_18602_),
    .B(_18603_),
    .CON(_02594_),
    .SN(_02595_));
 HAxp5_ASAP7_75t_R _34829_ (.A(_18604_),
    .B(_18605_),
    .CON(_00243_),
    .SN(_02596_));
 DFFHQNx1_ASAP7_75t_R _34830_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02597_),
    .QN(_01723_));
 DFFHQNx1_ASAP7_75t_R _34831_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02598_),
    .QN(_00164_));
 DFFHQNx1_ASAP7_75t_R _34832_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02599_),
    .QN(_00166_));
 DFFHQNx1_ASAP7_75t_R _34833_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02600_),
    .QN(_00169_));
 DFFHQNx1_ASAP7_75t_R _34834_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02601_),
    .QN(_00173_));
 DFFHQNx1_ASAP7_75t_R _34835_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02602_),
    .QN(_00176_));
 DFFHQNx1_ASAP7_75t_R _34836_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02603_),
    .QN(_00179_));
 DFFHQNx1_ASAP7_75t_R _34837_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02604_),
    .QN(_00181_));
 DFFHQNx1_ASAP7_75t_R _34838_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02605_),
    .QN(_00185_));
 DFFHQNx1_ASAP7_75t_R _34839_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02606_),
    .QN(_00188_));
 DFFHQNx1_ASAP7_75t_R _34840_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02607_),
    .QN(_00192_));
 DFFHQNx1_ASAP7_75t_R _34841_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02608_),
    .QN(_00195_));
 DFFHQNx1_ASAP7_75t_R _34842_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02609_),
    .QN(_00198_));
 DFFHQNx1_ASAP7_75t_R _34843_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02610_),
    .QN(_00200_));
 DFFHQNx1_ASAP7_75t_R _34844_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02611_),
    .QN(_00203_));
 DFFHQNx1_ASAP7_75t_R _34845_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_02612_),
    .QN(_00205_));
 DFFHQNx1_ASAP7_75t_R _34846_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02613_),
    .QN(_00385_));
 DFFHQNx1_ASAP7_75t_R _34847_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02614_),
    .QN(_01722_));
 DFFHQNx1_ASAP7_75t_R _34848_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02615_),
    .QN(_01721_));
 DFFHQNx1_ASAP7_75t_R _34849_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02616_),
    .QN(_01720_));
 DFFHQNx1_ASAP7_75t_R _34850_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02617_),
    .QN(_00162_));
 DFFHQNx1_ASAP7_75t_R _34851_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02618_),
    .QN(_00170_));
 DFFHQNx1_ASAP7_75t_R _34852_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02619_),
    .QN(_00174_));
 DFFHQNx1_ASAP7_75t_R _34853_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02620_),
    .QN(_00177_));
 DFFHQNx1_ASAP7_75t_R _34854_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02621_),
    .QN(_00180_));
 DFFHQNx1_ASAP7_75t_R _34855_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02622_),
    .QN(_00182_));
 DFFHQNx1_ASAP7_75t_R _34856_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02623_),
    .QN(_00186_));
 DFFHQNx1_ASAP7_75t_R _34857_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02624_),
    .QN(_00189_));
 DFFHQNx1_ASAP7_75t_R _34858_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02625_),
    .QN(_00193_));
 DFFHQNx1_ASAP7_75t_R _34859_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02626_),
    .QN(_00196_));
 DFFHQNx1_ASAP7_75t_R _34860_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02627_),
    .QN(_00199_));
 DFFHQNx1_ASAP7_75t_R _34861_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02628_),
    .QN(_00201_));
 DFFHQNx1_ASAP7_75t_R _34862_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02629_),
    .QN(_00204_));
 DFFHQNx1_ASAP7_75t_R _34863_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02630_),
    .QN(_00206_));
 DFFHQNx1_ASAP7_75t_R _34864_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02631_),
    .QN(_00208_));
 DFFHQNx1_ASAP7_75t_R _34865_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02632_),
    .QN(_00209_));
 DFFHQNx1_ASAP7_75t_R _34866_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02633_),
    .QN(_00211_));
 DFFHQNx1_ASAP7_75t_R _34867_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02634_),
    .QN(_00212_));
 DFFHQNx1_ASAP7_75t_R _34868_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02635_),
    .QN(_00214_));
 DFFHQNx1_ASAP7_75t_R _34869_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02636_),
    .QN(_00215_));
 DFFHQNx1_ASAP7_75t_R _34870_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02637_),
    .QN(_00217_));
 DFFHQNx1_ASAP7_75t_R _34871_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02638_),
    .QN(_00218_));
 DFFHQNx1_ASAP7_75t_R _34872_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02639_),
    .QN(_00220_));
 DFFHQNx1_ASAP7_75t_R _34873_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02640_),
    .QN(_00221_));
 DFFHQNx1_ASAP7_75t_R _34874_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02641_),
    .QN(_00223_));
 DFFHQNx1_ASAP7_75t_R _34875_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02642_),
    .QN(_00224_));
 DFFHQNx1_ASAP7_75t_R _34876_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02643_),
    .QN(_00226_));
 DFFHQNx1_ASAP7_75t_R _34877_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02644_),
    .QN(_00227_));
 DFFHQNx1_ASAP7_75t_R _34878_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02645_),
    .QN(_00229_));
 DFFHQNx1_ASAP7_75t_R _34879_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02646_),
    .QN(_00230_));
 DFFASRHQNx1_ASAP7_75t_R _34880_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.instr_valid_id_d ),
    .QN(_01317_),
    .RESETN(net467),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _34881_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.illegal_insn_d ),
    .QN(_01312_),
    .RESETN(net468),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34882_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.controller_i.exc_req_d ),
    .QN(_01724_),
    .RESETN(net469),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34883_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(net3059),
    .QN(_01725_),
    .RESETN(net470),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34884_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(net3039),
    .QN(_01719_),
    .RESETN(net471),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34885_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(net2644),
    .QN(_01718_),
    .RESETN(net472),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _34886_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02648_),
    .QN(_01717_),
    .RESETN(net473),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _34887_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02649_),
    .QN(_01716_),
    .RESETN(net474),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34888_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02650_),
    .QN(_01715_),
    .RESETN(net475),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _34889_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02651_),
    .QN(_01714_),
    .RESETN(net476),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _34890_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02652_),
    .QN(_01713_),
    .RESETN(net477),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34891_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02653_),
    .QN(_01712_),
    .RESETN(net478),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34892_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(net2533),
    .QN(_01711_),
    .RESETN(net479),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34893_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02655_),
    .QN(_01726_),
    .RESETN(net480),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34894_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(\id_stage_i.branch_set_d ),
    .QN(_01710_),
    .RESETN(net481),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _34895_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_02656_),
    .QN(_01709_),
    .RESETN(net482),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34896_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02657_),
    .QN(_01708_),
    .RESETN(net483),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34897_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_02658_),
    .QN(_01707_),
    .RESETN(net484),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _34898_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02659_),
    .QN(_01706_),
    .RESETN(net485),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34899_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02660_),
    .QN(_01705_),
    .RESETN(net486),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _34900_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02661_),
    .QN(_01704_),
    .RESETN(net487),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34901_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02662_),
    .QN(_01703_),
    .RESETN(net488),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34902_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02663_),
    .QN(_01702_),
    .RESETN(net489),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _34903_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_02664_),
    .QN(_01701_),
    .RESETN(net490),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34904_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02665_),
    .QN(_01700_),
    .RESETN(net491),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34905_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02666_),
    .QN(_01699_),
    .RESETN(net492),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _34906_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_02667_),
    .QN(_01698_),
    .RESETN(net493),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34907_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02668_),
    .QN(_01697_),
    .RESETN(net494),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34908_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02669_),
    .QN(_01696_),
    .RESETN(net495),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34909_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_02670_),
    .QN(_01695_),
    .RESETN(net496),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34910_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02671_),
    .QN(_01694_),
    .RESETN(net497),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34911_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_02672_),
    .QN(_01693_),
    .RESETN(net498),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _34912_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02673_),
    .QN(_01692_),
    .RESETN(net499),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34913_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02674_),
    .QN(_01691_),
    .RESETN(net500),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34914_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02675_),
    .QN(_01690_),
    .RESETN(net501),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34915_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02676_),
    .QN(_01689_),
    .RESETN(net502),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _34916_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02677_),
    .QN(_01688_),
    .RESETN(net503),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _34917_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02678_),
    .QN(_01687_),
    .RESETN(net504),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34918_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_02679_),
    .QN(_01686_),
    .RESETN(net505),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _34919_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02680_),
    .QN(_01685_),
    .RESETN(net506),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _34920_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02681_),
    .QN(_01684_),
    .RESETN(net507),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34921_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_02682_),
    .QN(_01683_),
    .RESETN(net508),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _34922_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02683_),
    .QN(_01682_),
    .RESETN(net509),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _34923_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02684_),
    .QN(_01681_),
    .RESETN(net510),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _34924_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_02685_),
    .QN(_01680_),
    .RESETN(net511),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _34925_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02686_),
    .QN(_01679_),
    .RESETN(net512),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _34926_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_02687_),
    .QN(_01678_),
    .RESETN(net513),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _34927_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02688_),
    .QN(_00324_),
    .RESETN(net514),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34928_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02689_),
    .QN(_00291_),
    .RESETN(net515),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34929_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02690_),
    .QN(_00663_),
    .RESETN(net516),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34930_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02691_),
    .QN(_00665_),
    .RESETN(net517),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34931_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02692_),
    .QN(_00668_),
    .RESETN(net518),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34932_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02693_),
    .QN(_00670_),
    .RESETN(net519),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34933_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02694_),
    .QN(_00672_),
    .RESETN(net520),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34934_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02695_),
    .QN(_00674_),
    .RESETN(net521),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34935_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02696_),
    .QN(_00677_),
    .RESETN(net522),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34936_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02697_),
    .QN(_00680_),
    .RESETN(net523),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34937_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02698_),
    .QN(_00682_),
    .RESETN(net524),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34938_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02699_),
    .QN(_00684_),
    .RESETN(net525),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34939_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02700_),
    .QN(_00686_),
    .RESETN(net526),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34940_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02701_),
    .QN(_00718_),
    .RESETN(net527),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34941_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02702_),
    .QN(_00750_),
    .RESETN(net528),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34942_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02703_),
    .QN(_00783_),
    .RESETN(net529),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34943_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02704_),
    .QN(_00816_),
    .RESETN(net530),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34944_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02705_),
    .QN(_00849_),
    .RESETN(net531),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34945_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02706_),
    .QN(_00881_),
    .RESETN(net532),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34946_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02707_),
    .QN(_00914_),
    .RESETN(net533),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34947_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02708_),
    .QN(_00946_),
    .RESETN(net534),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34948_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02709_),
    .QN(_00979_),
    .RESETN(net535),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34949_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02710_),
    .QN(_01011_),
    .RESETN(net536),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34950_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02711_),
    .QN(_01045_),
    .RESETN(net537),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34951_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02712_),
    .QN(_01077_),
    .RESETN(net538),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34952_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02713_),
    .QN(_01110_),
    .RESETN(net539),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34953_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02714_),
    .QN(_01142_),
    .RESETN(net540),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34954_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02715_),
    .QN(_01176_),
    .RESETN(net541),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34955_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02716_),
    .QN(_01208_),
    .RESETN(net542),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34956_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02717_),
    .QN(_01242_),
    .RESETN(net543),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34957_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02718_),
    .QN(_01274_),
    .RESETN(net544),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34958_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_02719_),
    .QN(_01308_),
    .RESETN(net545),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _34959_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02720_),
    .QN(_01677_),
    .RESETN(net546),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34960_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_02721_),
    .QN(_00034_),
    .RESETN(net547),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _34961_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_00002_),
    .QN(_01727_),
    .RESETN(net548),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _34962_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_00003_),
    .QN(_01728_),
    .RESETN(net549),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34963_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_00004_),
    .QN(_00284_),
    .RESETN(net550),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34964_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_00005_),
    .QN(_01357_),
    .RESETN(net551),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _34965_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02722_),
    .QN(_01676_),
    .RESETN(net552),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34966_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02723_),
    .QN(_01675_),
    .RESETN(net553),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34967_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02724_),
    .QN(_01674_),
    .RESETN(net554),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34968_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02725_),
    .QN(_01673_),
    .RESETN(net555),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34969_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02726_),
    .QN(_01672_),
    .RESETN(net556),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34970_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02727_),
    .QN(_01671_),
    .RESETN(net557),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34971_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02728_),
    .QN(_01670_),
    .RESETN(net558),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34972_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02729_),
    .QN(_01669_),
    .RESETN(net559),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34973_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02730_),
    .QN(_01668_),
    .RESETN(net560),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34974_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02731_),
    .QN(_01667_),
    .RESETN(net561),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34975_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02732_),
    .QN(_01666_),
    .RESETN(net562),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34976_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02733_),
    .QN(_01665_),
    .RESETN(net563),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34977_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02734_),
    .QN(_01664_),
    .RESETN(net564),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34978_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02735_),
    .QN(_01663_),
    .RESETN(net565),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34979_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02736_),
    .QN(_01662_),
    .RESETN(net566),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34980_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02737_),
    .QN(_01661_),
    .RESETN(net567),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34981_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02738_),
    .QN(_01660_),
    .RESETN(net568),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34982_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02739_),
    .QN(_01659_),
    .RESETN(net569),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34983_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02740_),
    .QN(_01658_),
    .RESETN(net570),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34984_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02741_),
    .QN(_01657_),
    .RESETN(net571),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34985_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02742_),
    .QN(_01656_),
    .RESETN(net572),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34986_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02743_),
    .QN(_01655_),
    .RESETN(net573),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34987_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02744_),
    .QN(_01654_),
    .RESETN(net574),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34988_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02745_),
    .QN(_01653_),
    .RESETN(net575),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34989_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02746_),
    .QN(_01652_),
    .RESETN(net576),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34990_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02747_),
    .QN(_01651_),
    .RESETN(net577),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34991_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02748_),
    .QN(_01650_),
    .RESETN(net578),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34992_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02749_),
    .QN(_01649_),
    .RESETN(net579),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34993_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02750_),
    .QN(_01648_),
    .RESETN(net580),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34994_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02751_),
    .QN(_01647_),
    .RESETN(net581),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34995_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02752_),
    .QN(_01646_),
    .RESETN(net582),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _34996_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02753_),
    .QN(_01645_),
    .RESETN(net583),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _34997_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02754_),
    .QN(_01323_),
    .RESETN(net584),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _34998_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02755_),
    .QN(_01324_),
    .RESETN(net585),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _34999_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02756_),
    .QN(_01325_),
    .RESETN(net586),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35000_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02757_),
    .QN(_01327_),
    .RESETN(net587),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35001_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02758_),
    .QN(_01328_),
    .RESETN(net588),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35002_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02759_),
    .QN(_01329_),
    .RESETN(net589),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35003_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02760_),
    .QN(_01330_),
    .RESETN(net590),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35004_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02761_),
    .QN(_01331_),
    .RESETN(net591),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35005_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02762_),
    .QN(_01332_),
    .RESETN(net592),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35006_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02763_),
    .QN(_01333_),
    .RESETN(net593),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35007_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02764_),
    .QN(_01334_),
    .RESETN(net594),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35008_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02765_),
    .QN(_01335_),
    .RESETN(net595),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35009_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02766_),
    .QN(_01336_),
    .RESETN(net596),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35010_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02767_),
    .QN(_01337_),
    .RESETN(net597),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35011_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02768_),
    .QN(_01338_),
    .RESETN(net598),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35012_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02769_),
    .QN(_01339_),
    .RESETN(net599),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35013_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02770_),
    .QN(_01340_),
    .RESETN(net600),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35014_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02771_),
    .QN(_01341_),
    .RESETN(net601),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35015_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02772_),
    .QN(_01342_),
    .RESETN(net602),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35016_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02773_),
    .QN(_01343_),
    .RESETN(net603),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35017_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02774_),
    .QN(_01344_),
    .RESETN(net604),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35018_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02775_),
    .QN(_01345_),
    .RESETN(net605),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35019_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02776_),
    .QN(_01346_),
    .RESETN(net606),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35020_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02777_),
    .QN(_01347_),
    .RESETN(net607),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35021_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02778_),
    .QN(_01348_),
    .RESETN(net608),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35022_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02779_),
    .QN(_01349_),
    .RESETN(net609),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35023_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02780_),
    .QN(_01350_),
    .RESETN(net610),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35024_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_02781_),
    .QN(_01351_),
    .RESETN(net611),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35025_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02782_),
    .QN(_01352_),
    .RESETN(net612),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35026_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02783_),
    .QN(_01353_),
    .RESETN(net613),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35027_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02784_),
    .QN(_01354_),
    .RESETN(net614),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35028_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02785_),
    .QN(_01355_),
    .RESETN(net615),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35029_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02786_),
    .QN(_17818_),
    .RESETN(net616),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35030_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02787_),
    .QN(_17819_),
    .RESETN(net617),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35031_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_02788_),
    .QN(_17825_),
    .RESETN(net618),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35032_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02789_),
    .QN(_01322_),
    .RESETN(net619),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35033_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_02790_),
    .QN(_01318_),
    .RESETN(net620),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35034_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_02791_),
    .QN(_01316_),
    .RESETN(net621),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35035_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02792_),
    .QN(_01644_),
    .RESETN(net622),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35036_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02793_),
    .QN(_01643_),
    .RESETN(net623),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35037_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_02794_),
    .QN(_01642_),
    .RESETN(net624),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35038_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02795_),
    .QN(_01641_),
    .RESETN(net625),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35039_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02796_),
    .QN(_01640_),
    .RESETN(net626),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35040_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02797_),
    .QN(_01639_),
    .RESETN(net627),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35041_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02798_),
    .QN(_01638_),
    .RESETN(net628),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35042_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02799_),
    .QN(_01637_),
    .RESETN(net629),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35043_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02800_),
    .QN(_01636_),
    .RESETN(net630),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35044_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02801_),
    .QN(_01635_),
    .RESETN(net631),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35045_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02802_),
    .QN(_01634_),
    .RESETN(net632),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35046_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02803_),
    .QN(_01633_),
    .RESETN(net633),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35047_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02804_),
    .QN(_01632_),
    .RESETN(net634),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35048_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02805_),
    .QN(_01631_),
    .RESETN(net635),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35049_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02806_),
    .QN(_01630_),
    .RESETN(net636),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35050_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02807_),
    .QN(_01629_),
    .RESETN(net637),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35051_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02808_),
    .QN(_01628_),
    .RESETN(net638),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35052_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02809_),
    .QN(_01627_),
    .RESETN(net639),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35053_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02810_),
    .QN(_01626_),
    .RESETN(net640),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35054_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02811_),
    .QN(_01625_),
    .RESETN(net641),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35055_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02812_),
    .QN(_01624_),
    .RESETN(net642),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35056_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02813_),
    .QN(_01623_),
    .RESETN(net643),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35057_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02814_),
    .QN(_01622_),
    .RESETN(net644),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35058_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02815_),
    .QN(_01621_),
    .RESETN(net645),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35059_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02816_),
    .QN(_01620_),
    .RESETN(net646),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35060_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02817_),
    .QN(_01619_),
    .RESETN(net647),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35061_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02818_),
    .QN(_01618_),
    .RESETN(net648),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35062_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02819_),
    .QN(_01617_),
    .RESETN(net649),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35063_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02820_),
    .QN(_01616_),
    .RESETN(net650),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35064_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02821_),
    .QN(_01615_),
    .RESETN(net651),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35065_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02822_),
    .QN(_01614_),
    .RESETN(net652),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35066_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02823_),
    .QN(_01613_),
    .RESETN(net653),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35067_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02824_),
    .QN(_01612_),
    .RESETN(net654),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35068_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_02825_),
    .QN(_01611_),
    .RESETN(net655),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35069_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_02826_),
    .QN(_01610_),
    .RESETN(net656),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35070_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(net3032),
    .QN(_01609_),
    .RESETN(net657),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35071_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02828_),
    .QN(_01608_),
    .RESETN(net658),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35072_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(net2806),
    .QN(_00277_),
    .RESETN(net659),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35073_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(net2735),
    .QN(_01607_),
    .RESETN(net660),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35074_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_02831_),
    .QN(_18554_),
    .RESETN(net661),
    .SETN(net449));
 DFFHQNx1_ASAP7_75t_R _35075_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02832_),
    .QN(_00662_));
 DFFHQNx1_ASAP7_75t_R _35076_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02833_),
    .QN(_17754_));
 DFFHQNx1_ASAP7_75t_R _35077_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02834_),
    .QN(_01606_));
 DFFHQNx1_ASAP7_75t_R _35078_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02835_),
    .QN(_01605_));
 DFFHQNx1_ASAP7_75t_R _35079_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02836_),
    .QN(_01604_));
 DFFHQNx1_ASAP7_75t_R _35080_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02837_),
    .QN(_01603_));
 DFFHQNx1_ASAP7_75t_R _35081_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02838_),
    .QN(_01602_));
 DFFHQNx1_ASAP7_75t_R _35082_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02839_),
    .QN(_01601_));
 DFFHQNx1_ASAP7_75t_R _35083_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02840_),
    .QN(_01600_));
 DFFHQNx1_ASAP7_75t_R _35084_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02841_),
    .QN(_01599_));
 DFFHQNx1_ASAP7_75t_R _35085_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02842_),
    .QN(_01598_));
 DFFHQNx1_ASAP7_75t_R _35086_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02843_),
    .QN(_01597_));
 DFFHQNx1_ASAP7_75t_R _35087_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02844_),
    .QN(_01596_));
 DFFHQNx1_ASAP7_75t_R _35088_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02845_),
    .QN(_01595_));
 DFFHQNx1_ASAP7_75t_R _35089_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02846_),
    .QN(_01594_));
 DFFHQNx1_ASAP7_75t_R _35090_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02847_),
    .QN(_01593_));
 DFFHQNx1_ASAP7_75t_R _35091_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02848_),
    .QN(_01592_));
 DFFHQNx1_ASAP7_75t_R _35092_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02849_),
    .QN(_01591_));
 DFFHQNx1_ASAP7_75t_R _35093_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02850_),
    .QN(_01590_));
 DFFHQNx1_ASAP7_75t_R _35094_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02851_),
    .QN(_01589_));
 DFFHQNx1_ASAP7_75t_R _35095_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02852_),
    .QN(_01588_));
 DFFHQNx1_ASAP7_75t_R _35096_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02853_),
    .QN(_01587_));
 DFFHQNx1_ASAP7_75t_R _35097_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02854_),
    .QN(_01586_));
 DFFHQNx1_ASAP7_75t_R _35098_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02855_),
    .QN(_01585_));
 DFFHQNx1_ASAP7_75t_R _35099_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02856_),
    .QN(_01584_));
 DFFHQNx1_ASAP7_75t_R _35100_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02857_),
    .QN(_01583_));
 DFFHQNx1_ASAP7_75t_R _35101_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02858_),
    .QN(_01582_));
 DFFHQNx1_ASAP7_75t_R _35102_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02859_),
    .QN(_01581_));
 DFFHQNx1_ASAP7_75t_R _35103_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02860_),
    .QN(_01580_));
 DFFHQNx1_ASAP7_75t_R _35104_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02861_),
    .QN(_01579_));
 DFFHQNx1_ASAP7_75t_R _35105_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02862_),
    .QN(_01578_));
 DFFASRHQNx1_ASAP7_75t_R _35106_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02863_),
    .QN(_01577_),
    .RESETN(net453),
    .SETN(net662));
 DFFASRHQNx1_ASAP7_75t_R _35107_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02864_),
    .QN(_01576_),
    .RESETN(net453),
    .SETN(net663));
 DFFASRHQNx1_ASAP7_75t_R _35108_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02865_),
    .QN(_00658_),
    .RESETN(net664),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35109_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(net3528),
    .QN(_01575_),
    .RESETN(net665),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35110_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02867_),
    .QN(_00081_),
    .RESETN(net666),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35111_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_02868_),
    .QN(_00084_),
    .RESETN(net667),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35112_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(net3633),
    .QN(_00087_),
    .RESETN(net668),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _35113_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02870_),
    .QN(_00090_),
    .RESETN(net669),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35114_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02871_),
    .QN(_01574_),
    .RESETN(net670),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35115_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02872_),
    .QN(_01573_),
    .RESETN(net671),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35116_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02873_),
    .QN(_01572_),
    .RESETN(net672),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35117_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02874_),
    .QN(_01571_),
    .RESETN(net673),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35118_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02875_),
    .QN(_01570_),
    .RESETN(net674),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35119_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02876_),
    .QN(_01569_),
    .RESETN(net675),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35120_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02877_),
    .QN(_01568_),
    .RESETN(net676),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35121_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02878_),
    .QN(_01567_),
    .RESETN(net677),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35122_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_02879_),
    .QN(_01566_),
    .RESETN(net678),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35123_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02880_),
    .QN(_01565_),
    .RESETN(net679),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35124_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02881_),
    .QN(_01564_),
    .RESETN(net680),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35125_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02882_),
    .QN(_01563_),
    .RESETN(net681),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35126_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02883_),
    .QN(_01562_),
    .RESETN(net682),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35127_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_02884_),
    .QN(_01561_),
    .RESETN(net683),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35128_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02885_),
    .QN(_01560_),
    .RESETN(net684),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _35129_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02886_),
    .QN(_01559_),
    .RESETN(net685),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35130_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02887_),
    .QN(_01558_),
    .RESETN(net686),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _35131_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_02888_),
    .QN(_01557_),
    .RESETN(net687),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _35132_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_02889_),
    .QN(_01556_),
    .RESETN(net688),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _35133_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02890_),
    .QN(_01555_),
    .RESETN(net689),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _35134_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_02891_),
    .QN(_01554_),
    .RESETN(net690),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35135_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_02892_),
    .QN(_01553_),
    .RESETN(net691),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _35136_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02893_),
    .QN(_01552_),
    .RESETN(net692),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _35137_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_02894_),
    .QN(_01551_),
    .RESETN(net693),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _35138_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_02895_),
    .QN(_01550_),
    .RESETN(net694),
    .SETN(net456));
 DFFHQNx1_ASAP7_75t_R _35139_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02896_),
    .QN(_01549_));
 DFFHQNx1_ASAP7_75t_R _35140_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_02897_),
    .QN(_01548_));
 DFFHQNx1_ASAP7_75t_R _35141_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02898_),
    .QN(_01547_));
 DFFHQNx1_ASAP7_75t_R _35142_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02899_),
    .QN(_01546_));
 DFFHQNx1_ASAP7_75t_R _35143_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02900_),
    .QN(_01545_));
 DFFHQNx1_ASAP7_75t_R _35144_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02901_),
    .QN(_01544_));
 DFFHQNx1_ASAP7_75t_R _35145_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02902_),
    .QN(_01543_));
 DFFHQNx1_ASAP7_75t_R _35146_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02903_),
    .QN(_01542_));
 DFFHQNx1_ASAP7_75t_R _35147_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02904_),
    .QN(_01541_));
 DFFHQNx1_ASAP7_75t_R _35148_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02905_),
    .QN(_01540_));
 DFFHQNx1_ASAP7_75t_R _35149_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02906_),
    .QN(_01539_));
 DFFHQNx1_ASAP7_75t_R _35150_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02907_),
    .QN(_01538_));
 DFFHQNx1_ASAP7_75t_R _35151_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02908_),
    .QN(_01537_));
 DFFHQNx1_ASAP7_75t_R _35152_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_02909_),
    .QN(_01536_));
 DFFHQNx1_ASAP7_75t_R _35153_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02910_),
    .QN(_01535_));
 DFFHQNx1_ASAP7_75t_R _35154_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02911_),
    .QN(_01534_));
 DFFHQNx1_ASAP7_75t_R _35155_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02912_),
    .QN(_01533_));
 DFFHQNx1_ASAP7_75t_R _35156_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02913_),
    .QN(_01532_));
 DFFHQNx1_ASAP7_75t_R _35157_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02914_),
    .QN(_01531_));
 DFFHQNx1_ASAP7_75t_R _35158_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02915_),
    .QN(_01530_));
 DFFHQNx1_ASAP7_75t_R _35159_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02916_),
    .QN(_01529_));
 DFFHQNx1_ASAP7_75t_R _35160_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02917_),
    .QN(_01528_));
 DFFHQNx1_ASAP7_75t_R _35161_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02918_),
    .QN(_01527_));
 DFFHQNx1_ASAP7_75t_R _35162_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_02919_),
    .QN(_01526_));
 DFFHQNx1_ASAP7_75t_R _35163_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02920_),
    .QN(_01525_));
 DFFHQNx1_ASAP7_75t_R _35164_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02921_),
    .QN(_01524_));
 DFFHQNx1_ASAP7_75t_R _35165_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02922_),
    .QN(_01523_));
 DFFHQNx1_ASAP7_75t_R _35166_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02923_),
    .QN(_01522_));
 DFFHQNx1_ASAP7_75t_R _35167_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02924_),
    .QN(_01521_));
 DFFHQNx1_ASAP7_75t_R _35168_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_02925_),
    .QN(_01520_));
 DFFASRHQNx1_ASAP7_75t_R _35169_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02926_),
    .QN(_00293_),
    .RESETN(net695),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35170_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02927_),
    .QN(_00247_),
    .RESETN(net696),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35171_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_02928_),
    .QN(_00355_),
    .RESETN(net697),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35172_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02929_),
    .QN(_00386_),
    .RESETN(net698),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35173_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02930_),
    .QN(_00416_),
    .RESETN(net699),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35174_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02931_),
    .QN(_00446_),
    .RESETN(net700),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35175_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02932_),
    .QN(_00476_),
    .RESETN(net701),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35176_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_02933_),
    .QN(_00506_),
    .RESETN(net702),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35177_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_02934_),
    .QN(_00536_),
    .RESETN(net703),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35178_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02935_),
    .QN(_00566_),
    .RESETN(net704),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35179_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02936_),
    .QN(_00596_),
    .RESETN(net705),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35180_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_02937_),
    .QN(_00626_),
    .RESETN(net706),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35181_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02938_),
    .QN(_00325_),
    .RESETN(net707),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35182_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02939_),
    .QN(_00688_),
    .RESETN(net708),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35183_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_02940_),
    .QN(_00720_),
    .RESETN(net709),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35184_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02941_),
    .QN(_00753_),
    .RESETN(net710),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35185_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_02942_),
    .QN(_00786_),
    .RESETN(net711),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35186_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02943_),
    .QN(_00819_),
    .RESETN(net712),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35187_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02944_),
    .QN(_00851_),
    .RESETN(net713),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35188_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02945_),
    .QN(_00884_),
    .RESETN(net714),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35189_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02946_),
    .QN(_00916_),
    .RESETN(net715),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35190_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02947_),
    .QN(_00949_),
    .RESETN(net716),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35191_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_02948_),
    .QN(_00981_),
    .RESETN(net717),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35192_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02949_),
    .QN(_01015_),
    .RESETN(net718),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35193_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02950_),
    .QN(_01047_),
    .RESETN(net719),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35194_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_02951_),
    .QN(_01080_),
    .RESETN(net720),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35195_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_02952_),
    .QN(_01112_),
    .RESETN(net721),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35196_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02953_),
    .QN(_01146_),
    .RESETN(net722),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35197_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02954_),
    .QN(_01178_),
    .RESETN(net723),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35198_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02955_),
    .QN(_01212_),
    .RESETN(net724),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35199_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02956_),
    .QN(_01244_),
    .RESETN(net725),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35200_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02957_),
    .QN(_01278_),
    .RESETN(net726),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35201_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_02958_),
    .QN(_00294_),
    .RESETN(net727),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35202_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02959_),
    .QN(_00248_),
    .RESETN(net728),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35203_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_02960_),
    .QN(_00356_),
    .RESETN(net729),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35204_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02961_),
    .QN(_00387_),
    .RESETN(net730),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35205_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02962_),
    .QN(_00417_),
    .RESETN(net731),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35206_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02963_),
    .QN(_00447_),
    .RESETN(net732),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35207_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02964_),
    .QN(_00477_),
    .RESETN(net733),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35208_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_02965_),
    .QN(_00507_),
    .RESETN(net734),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35209_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_02966_),
    .QN(_00537_),
    .RESETN(net735),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35210_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02967_),
    .QN(_00567_),
    .RESETN(net736),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35211_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_02968_),
    .QN(_00597_),
    .RESETN(net737),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35212_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_02969_),
    .QN(_00627_),
    .RESETN(net738),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35213_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02970_),
    .QN(_00326_),
    .RESETN(net739),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35214_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02971_),
    .QN(_00689_),
    .RESETN(net740),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35215_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_02972_),
    .QN(_00721_),
    .RESETN(net741),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35216_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02973_),
    .QN(_00754_),
    .RESETN(net742),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35217_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_02974_),
    .QN(_00787_),
    .RESETN(net743),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35218_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_02975_),
    .QN(_00820_),
    .RESETN(net744),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35219_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02976_),
    .QN(_00852_),
    .RESETN(net745),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35220_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02977_),
    .QN(_00885_),
    .RESETN(net746),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35221_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_02978_),
    .QN(_00917_),
    .RESETN(net747),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35222_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02979_),
    .QN(_00950_),
    .RESETN(net748),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35223_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_02980_),
    .QN(_00982_),
    .RESETN(net749),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35224_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_02981_),
    .QN(_01016_),
    .RESETN(net750),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35225_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_02982_),
    .QN(_01048_),
    .RESETN(net751),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35226_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_02983_),
    .QN(_01081_),
    .RESETN(net752),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35227_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_02984_),
    .QN(_01113_),
    .RESETN(net753),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35228_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_02985_),
    .QN(_01147_),
    .RESETN(net754),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35229_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02986_),
    .QN(_01179_),
    .RESETN(net755),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35230_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_02987_),
    .QN(_01213_),
    .RESETN(net756),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35231_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_02988_),
    .QN(_01245_),
    .RESETN(net757),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35232_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_02989_),
    .QN(_01279_),
    .RESETN(net758),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35233_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_02990_),
    .QN(_00295_),
    .RESETN(net759),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35234_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_02991_),
    .QN(_00249_),
    .RESETN(net760),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35235_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_02992_),
    .QN(_00357_),
    .RESETN(net761),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35236_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_02993_),
    .QN(_00388_),
    .RESETN(net762),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35237_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_02994_),
    .QN(_00418_),
    .RESETN(net763),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35238_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_02995_),
    .QN(_00448_),
    .RESETN(net764),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35239_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_02996_),
    .QN(_00478_),
    .RESETN(net765),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35240_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_02997_),
    .QN(_00508_),
    .RESETN(net766),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35241_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_02998_),
    .QN(_00538_),
    .RESETN(net767),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35242_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_02999_),
    .QN(_00568_),
    .RESETN(net768),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35243_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03000_),
    .QN(_00598_),
    .RESETN(net769),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35244_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03001_),
    .QN(_00628_),
    .RESETN(net770),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35245_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03002_),
    .QN(_00327_),
    .RESETN(net771),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35246_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03003_),
    .QN(_00690_),
    .RESETN(net772),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35247_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03004_),
    .QN(_00722_),
    .RESETN(net773),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35248_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03005_),
    .QN(_00755_),
    .RESETN(net774),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35249_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03006_),
    .QN(_00788_),
    .RESETN(net775),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35250_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03007_),
    .QN(_00821_),
    .RESETN(net776),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35251_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03008_),
    .QN(_00853_),
    .RESETN(net777),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35252_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03009_),
    .QN(_00886_),
    .RESETN(net778),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35253_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03010_),
    .QN(_00918_),
    .RESETN(net779),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35254_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03011_),
    .QN(_00951_),
    .RESETN(net780),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35255_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03012_),
    .QN(_00983_),
    .RESETN(net781),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35256_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03013_),
    .QN(_01017_),
    .RESETN(net782),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35257_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03014_),
    .QN(_01049_),
    .RESETN(net783),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35258_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03015_),
    .QN(_01082_),
    .RESETN(net784),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35259_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03016_),
    .QN(_01114_),
    .RESETN(net785),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35260_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03017_),
    .QN(_01148_),
    .RESETN(net786),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35261_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03018_),
    .QN(_01180_),
    .RESETN(net787),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35262_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03019_),
    .QN(_01214_),
    .RESETN(net788),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35263_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03020_),
    .QN(_01246_),
    .RESETN(net789),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35264_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03021_),
    .QN(_01280_),
    .RESETN(net790),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35265_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03022_),
    .QN(_00296_),
    .RESETN(net791),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35266_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03023_),
    .QN(_00250_),
    .RESETN(net792),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35267_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03024_),
    .QN(_00358_),
    .RESETN(net793),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35268_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03025_),
    .QN(_00389_),
    .RESETN(net794),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35269_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03026_),
    .QN(_00419_),
    .RESETN(net795),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35270_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03027_),
    .QN(_00449_),
    .RESETN(net796),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35271_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03028_),
    .QN(_00479_),
    .RESETN(net797),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35272_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03029_),
    .QN(_00509_),
    .RESETN(net798),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35273_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03030_),
    .QN(_00539_),
    .RESETN(net799),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35274_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03031_),
    .QN(_00569_),
    .RESETN(net800),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35275_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03032_),
    .QN(_00599_),
    .RESETN(net801),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35276_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03033_),
    .QN(_00629_),
    .RESETN(net802),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35277_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03034_),
    .QN(_00328_),
    .RESETN(net803),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35278_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03035_),
    .QN(_00691_),
    .RESETN(net804),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35279_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03036_),
    .QN(_00723_),
    .RESETN(net805),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35280_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03037_),
    .QN(_00756_),
    .RESETN(net806),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35281_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03038_),
    .QN(_00789_),
    .RESETN(net807),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35282_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03039_),
    .QN(_00822_),
    .RESETN(net808),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35283_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03040_),
    .QN(_00854_),
    .RESETN(net809),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35284_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03041_),
    .QN(_00887_),
    .RESETN(net810),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35285_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03042_),
    .QN(_00919_),
    .RESETN(net811),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35286_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03043_),
    .QN(_00952_),
    .RESETN(net812),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35287_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03044_),
    .QN(_00984_),
    .RESETN(net813),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35288_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03045_),
    .QN(_01018_),
    .RESETN(net814),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35289_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03046_),
    .QN(_01050_),
    .RESETN(net815),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35290_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03047_),
    .QN(_01083_),
    .RESETN(net816),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35291_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03048_),
    .QN(_01115_),
    .RESETN(net817),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35292_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03049_),
    .QN(_01149_),
    .RESETN(net818),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35293_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03050_),
    .QN(_01181_),
    .RESETN(net819),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35294_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03051_),
    .QN(_01215_),
    .RESETN(net820),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35295_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03052_),
    .QN(_01247_),
    .RESETN(net821),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35296_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03053_),
    .QN(_01281_),
    .RESETN(net822),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35297_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03054_),
    .QN(_00297_),
    .RESETN(net823),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35298_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03055_),
    .QN(_00251_),
    .RESETN(net824),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35299_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03056_),
    .QN(_00359_),
    .RESETN(net825),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35300_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03057_),
    .QN(_00390_),
    .RESETN(net826),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35301_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03058_),
    .QN(_00420_),
    .RESETN(net827),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35302_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03059_),
    .QN(_00450_),
    .RESETN(net828),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35303_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03060_),
    .QN(_00480_),
    .RESETN(net829),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35304_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03061_),
    .QN(_00510_),
    .RESETN(net830),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35305_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03062_),
    .QN(_00540_),
    .RESETN(net831),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35306_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03063_),
    .QN(_00570_),
    .RESETN(net832),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35307_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03064_),
    .QN(_00600_),
    .RESETN(net833),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35308_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03065_),
    .QN(_00630_),
    .RESETN(net834),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35309_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03066_),
    .QN(_00329_),
    .RESETN(net835),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35310_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03067_),
    .QN(_00692_),
    .RESETN(net836),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35311_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03068_),
    .QN(_00724_),
    .RESETN(net837),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35312_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03069_),
    .QN(_00757_),
    .RESETN(net838),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35313_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03070_),
    .QN(_00790_),
    .RESETN(net839),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35314_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03071_),
    .QN(_00823_),
    .RESETN(net840),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35315_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03072_),
    .QN(_00855_),
    .RESETN(net841),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35316_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03073_),
    .QN(_00888_),
    .RESETN(net842),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35317_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03074_),
    .QN(_00920_),
    .RESETN(net843),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35318_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03075_),
    .QN(_00953_),
    .RESETN(net844),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35319_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03076_),
    .QN(_00985_),
    .RESETN(net845),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35320_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03077_),
    .QN(_01019_),
    .RESETN(net846),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35321_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03078_),
    .QN(_01051_),
    .RESETN(net847),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35322_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03079_),
    .QN(_01084_),
    .RESETN(net848),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35323_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03080_),
    .QN(_01116_),
    .RESETN(net849),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35324_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03081_),
    .QN(_01150_),
    .RESETN(net850),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35325_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03082_),
    .QN(_01182_),
    .RESETN(net851),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35326_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03083_),
    .QN(_01216_),
    .RESETN(net852),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35327_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03084_),
    .QN(_01248_),
    .RESETN(net853),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35328_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03085_),
    .QN(_01282_),
    .RESETN(net854),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35329_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03086_),
    .QN(_00298_),
    .RESETN(net855),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35330_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03087_),
    .QN(_00252_),
    .RESETN(net856),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35331_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03088_),
    .QN(_00360_),
    .RESETN(net857),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35332_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03089_),
    .QN(_00391_),
    .RESETN(net858),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35333_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03090_),
    .QN(_00421_),
    .RESETN(net859),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35334_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03091_),
    .QN(_00451_),
    .RESETN(net860),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35335_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03092_),
    .QN(_00481_),
    .RESETN(net861),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35336_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03093_),
    .QN(_00511_),
    .RESETN(net862),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35337_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03094_),
    .QN(_00541_),
    .RESETN(net863),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35338_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03095_),
    .QN(_00571_),
    .RESETN(net864),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35339_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03096_),
    .QN(_00601_),
    .RESETN(net865),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35340_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03097_),
    .QN(_00631_),
    .RESETN(net866),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35341_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03098_),
    .QN(_00330_),
    .RESETN(net867),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35342_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03099_),
    .QN(_00693_),
    .RESETN(net868),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35343_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03100_),
    .QN(_00725_),
    .RESETN(net869),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35344_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03101_),
    .QN(_00758_),
    .RESETN(net870),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35345_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03102_),
    .QN(_00791_),
    .RESETN(net871),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35346_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03103_),
    .QN(_00824_),
    .RESETN(net872),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35347_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03104_),
    .QN(_00856_),
    .RESETN(net873),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35348_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03105_),
    .QN(_00889_),
    .RESETN(net874),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35349_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03106_),
    .QN(_00921_),
    .RESETN(net875),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35350_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03107_),
    .QN(_00954_),
    .RESETN(net876),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35351_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03108_),
    .QN(_00986_),
    .RESETN(net877),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35352_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03109_),
    .QN(_01020_),
    .RESETN(net878),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35353_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03110_),
    .QN(_01052_),
    .RESETN(net879),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35354_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03111_),
    .QN(_01085_),
    .RESETN(net880),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35355_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03112_),
    .QN(_01117_),
    .RESETN(net881),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35356_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03113_),
    .QN(_01151_),
    .RESETN(net882),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35357_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03114_),
    .QN(_01183_),
    .RESETN(net883),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35358_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03115_),
    .QN(_01217_),
    .RESETN(net884),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35359_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03116_),
    .QN(_01249_),
    .RESETN(net885),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35360_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03117_),
    .QN(_01283_),
    .RESETN(net886),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35361_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03118_),
    .QN(_00299_),
    .RESETN(net887),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35362_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03119_),
    .QN(_00253_),
    .RESETN(net888),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35363_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03120_),
    .QN(_00361_),
    .RESETN(net889),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35364_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03121_),
    .QN(_00392_),
    .RESETN(net890),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35365_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03122_),
    .QN(_00422_),
    .RESETN(net891),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35366_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03123_),
    .QN(_00452_),
    .RESETN(net892),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35367_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03124_),
    .QN(_00482_),
    .RESETN(net893),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35368_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03125_),
    .QN(_00512_),
    .RESETN(net894),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35369_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03126_),
    .QN(_00542_),
    .RESETN(net895),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35370_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03127_),
    .QN(_00572_),
    .RESETN(net896),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35371_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03128_),
    .QN(_00602_),
    .RESETN(net897),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35372_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03129_),
    .QN(_00632_),
    .RESETN(net898),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35373_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03130_),
    .QN(_00331_),
    .RESETN(net899),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35374_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03131_),
    .QN(_00694_),
    .RESETN(net900),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35375_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03132_),
    .QN(_00726_),
    .RESETN(net901),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35376_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03133_),
    .QN(_00759_),
    .RESETN(net902),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35377_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03134_),
    .QN(_00792_),
    .RESETN(net903),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35378_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03135_),
    .QN(_00825_),
    .RESETN(net904),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35379_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03136_),
    .QN(_00857_),
    .RESETN(net905),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35380_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03137_),
    .QN(_00890_),
    .RESETN(net906),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35381_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03138_),
    .QN(_00922_),
    .RESETN(net907),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35382_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03139_),
    .QN(_00955_),
    .RESETN(net908),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35383_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03140_),
    .QN(_00987_),
    .RESETN(net909),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35384_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03141_),
    .QN(_01021_),
    .RESETN(net910),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35385_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03142_),
    .QN(_01053_),
    .RESETN(net911),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35386_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03143_),
    .QN(_01086_),
    .RESETN(net912),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35387_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03144_),
    .QN(_01118_),
    .RESETN(net913),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35388_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03145_),
    .QN(_01152_),
    .RESETN(net914),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35389_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03146_),
    .QN(_01184_),
    .RESETN(net915),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35390_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03147_),
    .QN(_01218_),
    .RESETN(net916),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35391_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03148_),
    .QN(_01250_),
    .RESETN(net917),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35392_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03149_),
    .QN(_01284_),
    .RESETN(net918),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35393_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03150_),
    .QN(_00300_),
    .RESETN(net919),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35394_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03151_),
    .QN(_00254_),
    .RESETN(net920),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35395_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03152_),
    .QN(_00362_),
    .RESETN(net921),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35396_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03153_),
    .QN(_00393_),
    .RESETN(net922),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35397_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03154_),
    .QN(_00423_),
    .RESETN(net923),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35398_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03155_),
    .QN(_00453_),
    .RESETN(net924),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35399_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03156_),
    .QN(_00483_),
    .RESETN(net925),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35400_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03157_),
    .QN(_00513_),
    .RESETN(net926),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35401_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03158_),
    .QN(_00543_),
    .RESETN(net927),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35402_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03159_),
    .QN(_00573_),
    .RESETN(net928),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35403_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03160_),
    .QN(_00603_),
    .RESETN(net929),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35404_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03161_),
    .QN(_00633_),
    .RESETN(net930),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35405_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03162_),
    .QN(_00332_),
    .RESETN(net931),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35406_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03163_),
    .QN(_00695_),
    .RESETN(net932),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35407_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03164_),
    .QN(_00727_),
    .RESETN(net933),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35408_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03165_),
    .QN(_00760_),
    .RESETN(net934),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35409_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03166_),
    .QN(_00793_),
    .RESETN(net935),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35410_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03167_),
    .QN(_00826_),
    .RESETN(net936),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35411_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03168_),
    .QN(_00858_),
    .RESETN(net937),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35412_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03169_),
    .QN(_00891_),
    .RESETN(net938),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35413_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03170_),
    .QN(_00923_),
    .RESETN(net939),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35414_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03171_),
    .QN(_00956_),
    .RESETN(net940),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35415_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03172_),
    .QN(_00988_),
    .RESETN(net941),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35416_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03173_),
    .QN(_01022_),
    .RESETN(net942),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35417_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03174_),
    .QN(_01054_),
    .RESETN(net943),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35418_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03175_),
    .QN(_01087_),
    .RESETN(net944),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35419_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03176_),
    .QN(_01119_),
    .RESETN(net945),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35420_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03177_),
    .QN(_01153_),
    .RESETN(net946),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35421_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03178_),
    .QN(_01185_),
    .RESETN(net947),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35422_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03179_),
    .QN(_01219_),
    .RESETN(net948),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35423_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03180_),
    .QN(_01251_),
    .RESETN(net949),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35424_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03181_),
    .QN(_01285_),
    .RESETN(net950),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35425_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03182_),
    .QN(_00301_),
    .RESETN(net951),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35426_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03183_),
    .QN(_00255_),
    .RESETN(net952),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35427_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03184_),
    .QN(_00363_),
    .RESETN(net953),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35428_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03185_),
    .QN(_00394_),
    .RESETN(net954),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35429_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03186_),
    .QN(_00424_),
    .RESETN(net955),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35430_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03187_),
    .QN(_00454_),
    .RESETN(net956),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35431_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03188_),
    .QN(_00484_),
    .RESETN(net957),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35432_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03189_),
    .QN(_00514_),
    .RESETN(net958),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35433_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03190_),
    .QN(_00544_),
    .RESETN(net959),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35434_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03191_),
    .QN(_00574_),
    .RESETN(net960),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35435_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03192_),
    .QN(_00604_),
    .RESETN(net961),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35436_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03193_),
    .QN(_00634_),
    .RESETN(net962),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35437_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03194_),
    .QN(_00333_),
    .RESETN(net963),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35438_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03195_),
    .QN(_00696_),
    .RESETN(net964),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35439_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03196_),
    .QN(_00728_),
    .RESETN(net965),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35440_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03197_),
    .QN(_00761_),
    .RESETN(net966),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35441_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03198_),
    .QN(_00794_),
    .RESETN(net967),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35442_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03199_),
    .QN(_00827_),
    .RESETN(net968),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35443_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03200_),
    .QN(_00859_),
    .RESETN(net969),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35444_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03201_),
    .QN(_00892_),
    .RESETN(net970),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35445_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03202_),
    .QN(_00924_),
    .RESETN(net971),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35446_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03203_),
    .QN(_00957_),
    .RESETN(net972),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35447_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03204_),
    .QN(_00989_),
    .RESETN(net973),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35448_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03205_),
    .QN(_01023_),
    .RESETN(net974),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35449_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03206_),
    .QN(_01055_),
    .RESETN(net975),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35450_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03207_),
    .QN(_01088_),
    .RESETN(net976),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35451_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03208_),
    .QN(_01120_),
    .RESETN(net977),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35452_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03209_),
    .QN(_01154_),
    .RESETN(net978),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35453_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03210_),
    .QN(_01186_),
    .RESETN(net979),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35454_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03211_),
    .QN(_01220_),
    .RESETN(net980),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35455_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03212_),
    .QN(_01252_),
    .RESETN(net981),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35456_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03213_),
    .QN(_01286_),
    .RESETN(net982),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35457_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03214_),
    .QN(_00302_),
    .RESETN(net983),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35458_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03215_),
    .QN(_00256_),
    .RESETN(net984),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35459_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03216_),
    .QN(_00364_),
    .RESETN(net985),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35460_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03217_),
    .QN(_00395_),
    .RESETN(net986),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35461_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03218_),
    .QN(_00425_),
    .RESETN(net987),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35462_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03219_),
    .QN(_00455_),
    .RESETN(net988),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35463_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03220_),
    .QN(_00485_),
    .RESETN(net989),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35464_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03221_),
    .QN(_00515_),
    .RESETN(net990),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35465_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03222_),
    .QN(_00545_),
    .RESETN(net991),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35466_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03223_),
    .QN(_00575_),
    .RESETN(net992),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35467_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03224_),
    .QN(_00605_),
    .RESETN(net993),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35468_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03225_),
    .QN(_00635_),
    .RESETN(net994),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35469_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03226_),
    .QN(_00334_),
    .RESETN(net995),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35470_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03227_),
    .QN(_00697_),
    .RESETN(net996),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35471_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03228_),
    .QN(_00729_),
    .RESETN(net997),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35472_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03229_),
    .QN(_00762_),
    .RESETN(net998),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35473_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03230_),
    .QN(_00795_),
    .RESETN(net999),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35474_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03231_),
    .QN(_00828_),
    .RESETN(net1000),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35475_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03232_),
    .QN(_00860_),
    .RESETN(net1001),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35476_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03233_),
    .QN(_00893_),
    .RESETN(net1002),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35477_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03234_),
    .QN(_00925_),
    .RESETN(net1003),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35478_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03235_),
    .QN(_00958_),
    .RESETN(net1004),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35479_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03236_),
    .QN(_00990_),
    .RESETN(net1005),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35480_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03237_),
    .QN(_01024_),
    .RESETN(net1006),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35481_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03238_),
    .QN(_01056_),
    .RESETN(net1007),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35482_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03239_),
    .QN(_01089_),
    .RESETN(net1008),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35483_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03240_),
    .QN(_01121_),
    .RESETN(net1009),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35484_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03241_),
    .QN(_01155_),
    .RESETN(net1010),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35485_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03242_),
    .QN(_01187_),
    .RESETN(net1011),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35486_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03243_),
    .QN(_01221_),
    .RESETN(net1012),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35487_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03244_),
    .QN(_01253_),
    .RESETN(net1013),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35488_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03245_),
    .QN(_01287_),
    .RESETN(net1014),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35489_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03246_),
    .QN(_00303_),
    .RESETN(net1015),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35490_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03247_),
    .QN(_00257_),
    .RESETN(net1016),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35491_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03248_),
    .QN(_00365_),
    .RESETN(net1017),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35492_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03249_),
    .QN(_00396_),
    .RESETN(net1018),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35493_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03250_),
    .QN(_00426_),
    .RESETN(net1019),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35494_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03251_),
    .QN(_00456_),
    .RESETN(net1020),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35495_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03252_),
    .QN(_00486_),
    .RESETN(net1021),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35496_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03253_),
    .QN(_00516_),
    .RESETN(net1022),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35497_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03254_),
    .QN(_00546_),
    .RESETN(net1023),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35498_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03255_),
    .QN(_00576_),
    .RESETN(net1024),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35499_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03256_),
    .QN(_00606_),
    .RESETN(net1025),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35500_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03257_),
    .QN(_00636_),
    .RESETN(net1026),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35501_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03258_),
    .QN(_00335_),
    .RESETN(net1027),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35502_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03259_),
    .QN(_00698_),
    .RESETN(net1028),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35503_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03260_),
    .QN(_00730_),
    .RESETN(net1029),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35504_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03261_),
    .QN(_00763_),
    .RESETN(net1030),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35505_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03262_),
    .QN(_00796_),
    .RESETN(net1031),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35506_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03263_),
    .QN(_00829_),
    .RESETN(net1032),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35507_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03264_),
    .QN(_00861_),
    .RESETN(net1033),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35508_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03265_),
    .QN(_00894_),
    .RESETN(net1034),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35509_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03266_),
    .QN(_00926_),
    .RESETN(net1035),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35510_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03267_),
    .QN(_00959_),
    .RESETN(net1036),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35511_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03268_),
    .QN(_00991_),
    .RESETN(net1037),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35512_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03269_),
    .QN(_01025_),
    .RESETN(net1038),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35513_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03270_),
    .QN(_01057_),
    .RESETN(net1039),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35514_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03271_),
    .QN(_01090_),
    .RESETN(net1040),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35515_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03272_),
    .QN(_01122_),
    .RESETN(net1041),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35516_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03273_),
    .QN(_01156_),
    .RESETN(net1042),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35517_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03274_),
    .QN(_01188_),
    .RESETN(net1043),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35518_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03275_),
    .QN(_01222_),
    .RESETN(net1044),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35519_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03276_),
    .QN(_01254_),
    .RESETN(net1045),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35520_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03277_),
    .QN(_01288_),
    .RESETN(net1046),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35521_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03278_),
    .QN(_00304_),
    .RESETN(net1047),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35522_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03279_),
    .QN(_00258_),
    .RESETN(net1048),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35523_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03280_),
    .QN(_00366_),
    .RESETN(net1049),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35524_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03281_),
    .QN(_00397_),
    .RESETN(net1050),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35525_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03282_),
    .QN(_00427_),
    .RESETN(net1051),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35526_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03283_),
    .QN(_00457_),
    .RESETN(net1052),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35527_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03284_),
    .QN(_00487_),
    .RESETN(net1053),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35528_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03285_),
    .QN(_00517_),
    .RESETN(net1054),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35529_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03286_),
    .QN(_00547_),
    .RESETN(net1055),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35530_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03287_),
    .QN(_00577_),
    .RESETN(net1056),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35531_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03288_),
    .QN(_00607_),
    .RESETN(net1057),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35532_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03289_),
    .QN(_00637_),
    .RESETN(net1058),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35533_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03290_),
    .QN(_00336_),
    .RESETN(net1059),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35534_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03291_),
    .QN(_00699_),
    .RESETN(net1060),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35535_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03292_),
    .QN(_00731_),
    .RESETN(net1061),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35536_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03293_),
    .QN(_00764_),
    .RESETN(net1062),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35537_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03294_),
    .QN(_00797_),
    .RESETN(net1063),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35538_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03295_),
    .QN(_00830_),
    .RESETN(net1064),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35539_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03296_),
    .QN(_00862_),
    .RESETN(net1065),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35540_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03297_),
    .QN(_00895_),
    .RESETN(net1066),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35541_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03298_),
    .QN(_00927_),
    .RESETN(net1067),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35542_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03299_),
    .QN(_00960_),
    .RESETN(net1068),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35543_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03300_),
    .QN(_00992_),
    .RESETN(net1069),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35544_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03301_),
    .QN(_01026_),
    .RESETN(net1070),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35545_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03302_),
    .QN(_01058_),
    .RESETN(net1071),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35546_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03303_),
    .QN(_01091_),
    .RESETN(net1072),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35547_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03304_),
    .QN(_01123_),
    .RESETN(net1073),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35548_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03305_),
    .QN(_01157_),
    .RESETN(net1074),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35549_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03306_),
    .QN(_01189_),
    .RESETN(net1075),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35550_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03307_),
    .QN(_01223_),
    .RESETN(net1076),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35551_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03308_),
    .QN(_01255_),
    .RESETN(net1077),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35552_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03309_),
    .QN(_01289_),
    .RESETN(net1078),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35553_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03310_),
    .QN(_00305_),
    .RESETN(net1079),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35554_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03311_),
    .QN(_00259_),
    .RESETN(net1080),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35555_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03312_),
    .QN(_00367_),
    .RESETN(net1081),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35556_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03313_),
    .QN(_00398_),
    .RESETN(net1082),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35557_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03314_),
    .QN(_00428_),
    .RESETN(net1083),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35558_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03315_),
    .QN(_00458_),
    .RESETN(net1084),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35559_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03316_),
    .QN(_00488_),
    .RESETN(net1085),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35560_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03317_),
    .QN(_00518_),
    .RESETN(net1086),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35561_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03318_),
    .QN(_00548_),
    .RESETN(net1087),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35562_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03319_),
    .QN(_00578_),
    .RESETN(net1088),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35563_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03320_),
    .QN(_00608_),
    .RESETN(net1089),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35564_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03321_),
    .QN(_00638_),
    .RESETN(net1090),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35565_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03322_),
    .QN(_00337_),
    .RESETN(net1091),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35566_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03323_),
    .QN(_00700_),
    .RESETN(net1092),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35567_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03324_),
    .QN(_00732_),
    .RESETN(net1093),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35568_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03325_),
    .QN(_00765_),
    .RESETN(net1094),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35569_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03326_),
    .QN(_00798_),
    .RESETN(net1095),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35570_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03327_),
    .QN(_00831_),
    .RESETN(net1096),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35571_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03328_),
    .QN(_00863_),
    .RESETN(net1097),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35572_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03329_),
    .QN(_00896_),
    .RESETN(net1098),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35573_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03330_),
    .QN(_00928_),
    .RESETN(net1099),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35574_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03331_),
    .QN(_00961_),
    .RESETN(net1100),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35575_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03332_),
    .QN(_00993_),
    .RESETN(net1101),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35576_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03333_),
    .QN(_01027_),
    .RESETN(net1102),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35577_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03334_),
    .QN(_01059_),
    .RESETN(net1103),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35578_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03335_),
    .QN(_01092_),
    .RESETN(net1104),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35579_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03336_),
    .QN(_01124_),
    .RESETN(net1105),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35580_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03337_),
    .QN(_01158_),
    .RESETN(net1106),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35581_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03338_),
    .QN(_01190_),
    .RESETN(net1107),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35582_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03339_),
    .QN(_01224_),
    .RESETN(net1108),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35583_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03340_),
    .QN(_01256_),
    .RESETN(net1109),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35584_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03341_),
    .QN(_01290_),
    .RESETN(net1110),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35585_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03342_),
    .QN(_00306_),
    .RESETN(net1111),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35586_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03343_),
    .QN(_00260_),
    .RESETN(net1112),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35587_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03344_),
    .QN(_00368_),
    .RESETN(net1113),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35588_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03345_),
    .QN(_00399_),
    .RESETN(net1114),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35589_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03346_),
    .QN(_00429_),
    .RESETN(net1115),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35590_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03347_),
    .QN(_00459_),
    .RESETN(net1116),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35591_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03348_),
    .QN(_00489_),
    .RESETN(net1117),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35592_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03349_),
    .QN(_00519_),
    .RESETN(net1118),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35593_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03350_),
    .QN(_00549_),
    .RESETN(net1119),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35594_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03351_),
    .QN(_00579_),
    .RESETN(net1120),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35595_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03352_),
    .QN(_00609_),
    .RESETN(net1121),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35596_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03353_),
    .QN(_00639_),
    .RESETN(net1122),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35597_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03354_),
    .QN(_00338_),
    .RESETN(net1123),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35598_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03355_),
    .QN(_00701_),
    .RESETN(net1124),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35599_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03356_),
    .QN(_00733_),
    .RESETN(net1125),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35600_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03357_),
    .QN(_00766_),
    .RESETN(net1126),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35601_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03358_),
    .QN(_00799_),
    .RESETN(net1127),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35602_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03359_),
    .QN(_00832_),
    .RESETN(net1128),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35603_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03360_),
    .QN(_00864_),
    .RESETN(net1129),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35604_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03361_),
    .QN(_00897_),
    .RESETN(net1130),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35605_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03362_),
    .QN(_00929_),
    .RESETN(net1131),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35606_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03363_),
    .QN(_00962_),
    .RESETN(net1132),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35607_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03364_),
    .QN(_00994_),
    .RESETN(net1133),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35608_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03365_),
    .QN(_01028_),
    .RESETN(net1134),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35609_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03366_),
    .QN(_01060_),
    .RESETN(net1135),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35610_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03367_),
    .QN(_01093_),
    .RESETN(net1136),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35611_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03368_),
    .QN(_01125_),
    .RESETN(net1137),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35612_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03369_),
    .QN(_01159_),
    .RESETN(net1138),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35613_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03370_),
    .QN(_01191_),
    .RESETN(net1139),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35614_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03371_),
    .QN(_01225_),
    .RESETN(net1140),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35615_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03372_),
    .QN(_01257_),
    .RESETN(net1141),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35616_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03373_),
    .QN(_01291_),
    .RESETN(net1142),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35617_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03374_),
    .QN(_00307_),
    .RESETN(net1143),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35618_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03375_),
    .QN(_00261_),
    .RESETN(net1144),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35619_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03376_),
    .QN(_00369_),
    .RESETN(net1145),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35620_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03377_),
    .QN(_00400_),
    .RESETN(net1146),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35621_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03378_),
    .QN(_00430_),
    .RESETN(net1147),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35622_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03379_),
    .QN(_00460_),
    .RESETN(net1148),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35623_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03380_),
    .QN(_00490_),
    .RESETN(net1149),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35624_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03381_),
    .QN(_00520_),
    .RESETN(net1150),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35625_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03382_),
    .QN(_00550_),
    .RESETN(net1151),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35626_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03383_),
    .QN(_00580_),
    .RESETN(net1152),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35627_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03384_),
    .QN(_00610_),
    .RESETN(net1153),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35628_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03385_),
    .QN(_00640_),
    .RESETN(net1154),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35629_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03386_),
    .QN(_00339_),
    .RESETN(net1155),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35630_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03387_),
    .QN(_00702_),
    .RESETN(net1156),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35631_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03388_),
    .QN(_00734_),
    .RESETN(net1157),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35632_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03389_),
    .QN(_00767_),
    .RESETN(net1158),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35633_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03390_),
    .QN(_00800_),
    .RESETN(net1159),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35634_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03391_),
    .QN(_00833_),
    .RESETN(net1160),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35635_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03392_),
    .QN(_00865_),
    .RESETN(net1161),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35636_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03393_),
    .QN(_00898_),
    .RESETN(net1162),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35637_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03394_),
    .QN(_00930_),
    .RESETN(net1163),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35638_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03395_),
    .QN(_00963_),
    .RESETN(net1164),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35639_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03396_),
    .QN(_00995_),
    .RESETN(net1165),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35640_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03397_),
    .QN(_01029_),
    .RESETN(net1166),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35641_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03398_),
    .QN(_01061_),
    .RESETN(net1167),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35642_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03399_),
    .QN(_01094_),
    .RESETN(net1168),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35643_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03400_),
    .QN(_01126_),
    .RESETN(net1169),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35644_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03401_),
    .QN(_01160_),
    .RESETN(net1170),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35645_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03402_),
    .QN(_01192_),
    .RESETN(net1171),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35646_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03403_),
    .QN(_01226_),
    .RESETN(net1172),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35647_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03404_),
    .QN(_01258_),
    .RESETN(net1173),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35648_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03405_),
    .QN(_01292_),
    .RESETN(net1174),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35649_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03406_),
    .QN(_00308_),
    .RESETN(net1175),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35650_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03407_),
    .QN(_00262_),
    .RESETN(net1176),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35651_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03408_),
    .QN(_00370_),
    .RESETN(net1177),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35652_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03409_),
    .QN(_00401_),
    .RESETN(net1178),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35653_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03410_),
    .QN(_00431_),
    .RESETN(net1179),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35654_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03411_),
    .QN(_00461_),
    .RESETN(net1180),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35655_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03412_),
    .QN(_00491_),
    .RESETN(net1181),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35656_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03413_),
    .QN(_00521_),
    .RESETN(net1182),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35657_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03414_),
    .QN(_00551_),
    .RESETN(net1183),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35658_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03415_),
    .QN(_00581_),
    .RESETN(net1184),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35659_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03416_),
    .QN(_00611_),
    .RESETN(net1185),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35660_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03417_),
    .QN(_00641_),
    .RESETN(net1186),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35661_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03418_),
    .QN(_00340_),
    .RESETN(net1187),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35662_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03419_),
    .QN(_00703_),
    .RESETN(net1188),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35663_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03420_),
    .QN(_00735_),
    .RESETN(net1189),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35664_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03421_),
    .QN(_00768_),
    .RESETN(net1190),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35665_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03422_),
    .QN(_00801_),
    .RESETN(net1191),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35666_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03423_),
    .QN(_00834_),
    .RESETN(net1192),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35667_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03424_),
    .QN(_00866_),
    .RESETN(net1193),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35668_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03425_),
    .QN(_00899_),
    .RESETN(net1194),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35669_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03426_),
    .QN(_00931_),
    .RESETN(net1195),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35670_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03427_),
    .QN(_00964_),
    .RESETN(net1196),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35671_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03428_),
    .QN(_00996_),
    .RESETN(net1197),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35672_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03429_),
    .QN(_01030_),
    .RESETN(net1198),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35673_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03430_),
    .QN(_01062_),
    .RESETN(net1199),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35674_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03431_),
    .QN(_01095_),
    .RESETN(net1200),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35675_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03432_),
    .QN(_01127_),
    .RESETN(net1201),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35676_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03433_),
    .QN(_01161_),
    .RESETN(net1202),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35677_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03434_),
    .QN(_01193_),
    .RESETN(net1203),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35678_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03435_),
    .QN(_01227_),
    .RESETN(net1204),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35679_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03436_),
    .QN(_01259_),
    .RESETN(net1205),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35680_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03437_),
    .QN(_01293_),
    .RESETN(net1206),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35681_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03438_),
    .QN(_00309_),
    .RESETN(net1207),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35682_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03439_),
    .QN(_00263_),
    .RESETN(net1208),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35683_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03440_),
    .QN(_00371_),
    .RESETN(net1209),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35684_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03441_),
    .QN(_00402_),
    .RESETN(net1210),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35685_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03442_),
    .QN(_00432_),
    .RESETN(net1211),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35686_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03443_),
    .QN(_00462_),
    .RESETN(net1212),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35687_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03444_),
    .QN(_00492_),
    .RESETN(net1213),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35688_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03445_),
    .QN(_00522_),
    .RESETN(net1214),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35689_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03446_),
    .QN(_00552_),
    .RESETN(net1215),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35690_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03447_),
    .QN(_00582_),
    .RESETN(net1216),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35691_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03448_),
    .QN(_00612_),
    .RESETN(net1217),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35692_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03449_),
    .QN(_00642_),
    .RESETN(net1218),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35693_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03450_),
    .QN(_00341_),
    .RESETN(net1219),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35694_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03451_),
    .QN(_00704_),
    .RESETN(net1220),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35695_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03452_),
    .QN(_00736_),
    .RESETN(net1221),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35696_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03453_),
    .QN(_00769_),
    .RESETN(net1222),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35697_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03454_),
    .QN(_00802_),
    .RESETN(net1223),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35698_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03455_),
    .QN(_00835_),
    .RESETN(net1224),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35699_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03456_),
    .QN(_00867_),
    .RESETN(net1225),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35700_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03457_),
    .QN(_00900_),
    .RESETN(net1226),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35701_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03458_),
    .QN(_00932_),
    .RESETN(net1227),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35702_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03459_),
    .QN(_00965_),
    .RESETN(net1228),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35703_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03460_),
    .QN(_00997_),
    .RESETN(net1229),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35704_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03461_),
    .QN(_01031_),
    .RESETN(net1230),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35705_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03462_),
    .QN(_01063_),
    .RESETN(net1231),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35706_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03463_),
    .QN(_01096_),
    .RESETN(net1232),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35707_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03464_),
    .QN(_01128_),
    .RESETN(net1233),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35708_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03465_),
    .QN(_01162_),
    .RESETN(net1234),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35709_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03466_),
    .QN(_01194_),
    .RESETN(net1235),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35710_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03467_),
    .QN(_01228_),
    .RESETN(net1236),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35711_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03468_),
    .QN(_01260_),
    .RESETN(net1237),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35712_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03469_),
    .QN(_01294_),
    .RESETN(net1238),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35713_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03470_),
    .QN(_00310_),
    .RESETN(net1239),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35714_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03471_),
    .QN(_00264_),
    .RESETN(net1240),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35715_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03472_),
    .QN(_00372_),
    .RESETN(net1241),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35716_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03473_),
    .QN(_00403_),
    .RESETN(net1242),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35717_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03474_),
    .QN(_00433_),
    .RESETN(net1243),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35718_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03475_),
    .QN(_00463_),
    .RESETN(net1244),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35719_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03476_),
    .QN(_00493_),
    .RESETN(net1245),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35720_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03477_),
    .QN(_00523_),
    .RESETN(net1246),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35721_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03478_),
    .QN(_00553_),
    .RESETN(net1247),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35722_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03479_),
    .QN(_00583_),
    .RESETN(net1248),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35723_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03480_),
    .QN(_00613_),
    .RESETN(net1249),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35724_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03481_),
    .QN(_00643_),
    .RESETN(net1250),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35725_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03482_),
    .QN(_00342_),
    .RESETN(net1251),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35726_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03483_),
    .QN(_00705_),
    .RESETN(net1252),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35727_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03484_),
    .QN(_00737_),
    .RESETN(net1253),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35728_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03485_),
    .QN(_00770_),
    .RESETN(net1254),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35729_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03486_),
    .QN(_00803_),
    .RESETN(net1255),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35730_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03487_),
    .QN(_00836_),
    .RESETN(net1256),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35731_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03488_),
    .QN(_00868_),
    .RESETN(net1257),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35732_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03489_),
    .QN(_00901_),
    .RESETN(net1258),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35733_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03490_),
    .QN(_00933_),
    .RESETN(net1259),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35734_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03491_),
    .QN(_00966_),
    .RESETN(net1260),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35735_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03492_),
    .QN(_00998_),
    .RESETN(net1261),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35736_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03493_),
    .QN(_01032_),
    .RESETN(net1262),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35737_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03494_),
    .QN(_01064_),
    .RESETN(net1263),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35738_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03495_),
    .QN(_01097_),
    .RESETN(net1264),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35739_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03496_),
    .QN(_01129_),
    .RESETN(net1265),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35740_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03497_),
    .QN(_01163_),
    .RESETN(net1266),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35741_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03498_),
    .QN(_01195_),
    .RESETN(net1267),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35742_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03499_),
    .QN(_01229_),
    .RESETN(net1268),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35743_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03500_),
    .QN(_01261_),
    .RESETN(net1269),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35744_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03501_),
    .QN(_01295_),
    .RESETN(net1270),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35745_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03502_),
    .QN(_00311_),
    .RESETN(net1271),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35746_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03503_),
    .QN(_00265_),
    .RESETN(net1272),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35747_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03504_),
    .QN(_00373_),
    .RESETN(net1273),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35748_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03505_),
    .QN(_00404_),
    .RESETN(net1274),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35749_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03506_),
    .QN(_00434_),
    .RESETN(net1275),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35750_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03507_),
    .QN(_00464_),
    .RESETN(net1276),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35751_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03508_),
    .QN(_00494_),
    .RESETN(net1277),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35752_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03509_),
    .QN(_00524_),
    .RESETN(net1278),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35753_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03510_),
    .QN(_00554_),
    .RESETN(net1279),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35754_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03511_),
    .QN(_00584_),
    .RESETN(net1280),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35755_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03512_),
    .QN(_00614_),
    .RESETN(net1281),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35756_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03513_),
    .QN(_00644_),
    .RESETN(net1282),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35757_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03514_),
    .QN(_00343_),
    .RESETN(net1283),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35758_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03515_),
    .QN(_00706_),
    .RESETN(net1284),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35759_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03516_),
    .QN(_00738_),
    .RESETN(net1285),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35760_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03517_),
    .QN(_00771_),
    .RESETN(net1286),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35761_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03518_),
    .QN(_00804_),
    .RESETN(net1287),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35762_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03519_),
    .QN(_00837_),
    .RESETN(net1288),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35763_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03520_),
    .QN(_00869_),
    .RESETN(net1289),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35764_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03521_),
    .QN(_00902_),
    .RESETN(net1290),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35765_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03522_),
    .QN(_00934_),
    .RESETN(net1291),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35766_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03523_),
    .QN(_00967_),
    .RESETN(net1292),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35767_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03524_),
    .QN(_00999_),
    .RESETN(net1293),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35768_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03525_),
    .QN(_01033_),
    .RESETN(net1294),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35769_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03526_),
    .QN(_01065_),
    .RESETN(net1295),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35770_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03527_),
    .QN(_01098_),
    .RESETN(net1296),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35771_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03528_),
    .QN(_01130_),
    .RESETN(net1297),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35772_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03529_),
    .QN(_01164_),
    .RESETN(net1298),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35773_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03530_),
    .QN(_01196_),
    .RESETN(net1299),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35774_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03531_),
    .QN(_01230_),
    .RESETN(net1300),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35775_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03532_),
    .QN(_01262_),
    .RESETN(net1301),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35776_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03533_),
    .QN(_01296_),
    .RESETN(net1302),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35777_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03534_),
    .QN(_00312_),
    .RESETN(net1303),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35778_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03535_),
    .QN(_00266_),
    .RESETN(net1304),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35779_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03536_),
    .QN(_00374_),
    .RESETN(net1305),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35780_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03537_),
    .QN(_00405_),
    .RESETN(net1306),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35781_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03538_),
    .QN(_00435_),
    .RESETN(net1307),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35782_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03539_),
    .QN(_00465_),
    .RESETN(net1308),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35783_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03540_),
    .QN(_00495_),
    .RESETN(net1309),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35784_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03541_),
    .QN(_00525_),
    .RESETN(net1310),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35785_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03542_),
    .QN(_00555_),
    .RESETN(net1311),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35786_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03543_),
    .QN(_00585_),
    .RESETN(net1312),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35787_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03544_),
    .QN(_00615_),
    .RESETN(net1313),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35788_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03545_),
    .QN(_00645_),
    .RESETN(net1314),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35789_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03546_),
    .QN(_00344_),
    .RESETN(net1315),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35790_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03547_),
    .QN(_00707_),
    .RESETN(net1316),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35791_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03548_),
    .QN(_00739_),
    .RESETN(net1317),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35792_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03549_),
    .QN(_00772_),
    .RESETN(net1318),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35793_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03550_),
    .QN(_00805_),
    .RESETN(net1319),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35794_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03551_),
    .QN(_00838_),
    .RESETN(net1320),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35795_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03552_),
    .QN(_00870_),
    .RESETN(net1321),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35796_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03553_),
    .QN(_00903_),
    .RESETN(net1322),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35797_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03554_),
    .QN(_00935_),
    .RESETN(net1323),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35798_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03555_),
    .QN(_00968_),
    .RESETN(net1324),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35799_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03556_),
    .QN(_01000_),
    .RESETN(net1325),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35800_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03557_),
    .QN(_01034_),
    .RESETN(net1326),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35801_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03558_),
    .QN(_01066_),
    .RESETN(net1327),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35802_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03559_),
    .QN(_01099_),
    .RESETN(net1328),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35803_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03560_),
    .QN(_01131_),
    .RESETN(net1329),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35804_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03561_),
    .QN(_01165_),
    .RESETN(net1330),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35805_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03562_),
    .QN(_01197_),
    .RESETN(net1331),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35806_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03563_),
    .QN(_01231_),
    .RESETN(net1332),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35807_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03564_),
    .QN(_01263_),
    .RESETN(net1333),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35808_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03565_),
    .QN(_01297_),
    .RESETN(net1334),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35809_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03566_),
    .QN(_00313_),
    .RESETN(net1335),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35810_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03567_),
    .QN(_00267_),
    .RESETN(net1336),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35811_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03568_),
    .QN(_00375_),
    .RESETN(net1337),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35812_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03569_),
    .QN(_00406_),
    .RESETN(net1338),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35813_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03570_),
    .QN(_00436_),
    .RESETN(net1339),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35814_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03571_),
    .QN(_00466_),
    .RESETN(net1340),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35815_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03572_),
    .QN(_00496_),
    .RESETN(net1341),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35816_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03573_),
    .QN(_00526_),
    .RESETN(net1342),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35817_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03574_),
    .QN(_00556_),
    .RESETN(net1343),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35818_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03575_),
    .QN(_00586_),
    .RESETN(net1344),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35819_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03576_),
    .QN(_00616_),
    .RESETN(net1345),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35820_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03577_),
    .QN(_00646_),
    .RESETN(net1346),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35821_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03578_),
    .QN(_00345_),
    .RESETN(net1347),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35822_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03579_),
    .QN(_00708_),
    .RESETN(net1348),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35823_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03580_),
    .QN(_00740_),
    .RESETN(net1349),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35824_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03581_),
    .QN(_00773_),
    .RESETN(net1350),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35825_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03582_),
    .QN(_00806_),
    .RESETN(net1351),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35826_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03583_),
    .QN(_00839_),
    .RESETN(net1352),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35827_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03584_),
    .QN(_00871_),
    .RESETN(net1353),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35828_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03585_),
    .QN(_00904_),
    .RESETN(net1354),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35829_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03586_),
    .QN(_00936_),
    .RESETN(net1355),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35830_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03587_),
    .QN(_00969_),
    .RESETN(net1356),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35831_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03588_),
    .QN(_01001_),
    .RESETN(net1357),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35832_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03589_),
    .QN(_01035_),
    .RESETN(net1358),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35833_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03590_),
    .QN(_01067_),
    .RESETN(net1359),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35834_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03591_),
    .QN(_01100_),
    .RESETN(net1360),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35835_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03592_),
    .QN(_01132_),
    .RESETN(net1361),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35836_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03593_),
    .QN(_01166_),
    .RESETN(net1362),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35837_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03594_),
    .QN(_01198_),
    .RESETN(net1363),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35838_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03595_),
    .QN(_01232_),
    .RESETN(net1364),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35839_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03596_),
    .QN(_01264_),
    .RESETN(net1365),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35840_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03597_),
    .QN(_01298_),
    .RESETN(net1366),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35841_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03598_),
    .QN(_00314_),
    .RESETN(net1367),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35842_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03599_),
    .QN(_00268_),
    .RESETN(net1368),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35843_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03600_),
    .QN(_00376_),
    .RESETN(net1369),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35844_ (.CLK(clknet_level_3_1_31123_clk_i),
    .D(_03601_),
    .QN(_00407_),
    .RESETN(net1370),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35845_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03602_),
    .QN(_00437_),
    .RESETN(net1371),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35846_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03603_),
    .QN(_00467_),
    .RESETN(net1372),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35847_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03604_),
    .QN(_00497_),
    .RESETN(net1373),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35848_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03605_),
    .QN(_00527_),
    .RESETN(net1374),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35849_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03606_),
    .QN(_00557_),
    .RESETN(net1375),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35850_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03607_),
    .QN(_00587_),
    .RESETN(net1376),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35851_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03608_),
    .QN(_00617_),
    .RESETN(net1377),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35852_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03609_),
    .QN(_00647_),
    .RESETN(net1378),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35853_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03610_),
    .QN(_00346_),
    .RESETN(net1379),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35854_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03611_),
    .QN(_00709_),
    .RESETN(net1380),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35855_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03612_),
    .QN(_00741_),
    .RESETN(net1381),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35856_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03613_),
    .QN(_00774_),
    .RESETN(net1382),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35857_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03614_),
    .QN(_00807_),
    .RESETN(net1383),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35858_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03615_),
    .QN(_00840_),
    .RESETN(net1384),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35859_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03616_),
    .QN(_00872_),
    .RESETN(net1385),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35860_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03617_),
    .QN(_00905_),
    .RESETN(net1386),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35861_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03618_),
    .QN(_00937_),
    .RESETN(net1387),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35862_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03619_),
    .QN(_00970_),
    .RESETN(net1388),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35863_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03620_),
    .QN(_01002_),
    .RESETN(net1389),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35864_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03621_),
    .QN(_01036_),
    .RESETN(net1390),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35865_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03622_),
    .QN(_01068_),
    .RESETN(net1391),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35866_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03623_),
    .QN(_01101_),
    .RESETN(net1392),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35867_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03624_),
    .QN(_01133_),
    .RESETN(net1393),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35868_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03625_),
    .QN(_01167_),
    .RESETN(net1394),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35869_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03626_),
    .QN(_01199_),
    .RESETN(net1395),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35870_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03627_),
    .QN(_01233_),
    .RESETN(net1396),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35871_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03628_),
    .QN(_01265_),
    .RESETN(net1397),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35872_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03629_),
    .QN(_01299_),
    .RESETN(net1398),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35873_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03630_),
    .QN(_00315_),
    .RESETN(net1399),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35874_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03631_),
    .QN(_00269_),
    .RESETN(net1400),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35875_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03632_),
    .QN(_00377_),
    .RESETN(net1401),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35876_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03633_),
    .QN(_00408_),
    .RESETN(net1402),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35877_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03634_),
    .QN(_00438_),
    .RESETN(net1403),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35878_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03635_),
    .QN(_00468_),
    .RESETN(net1404),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35879_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03636_),
    .QN(_00498_),
    .RESETN(net1405),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35880_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03637_),
    .QN(_00528_),
    .RESETN(net1406),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35881_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03638_),
    .QN(_00558_),
    .RESETN(net1407),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35882_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03639_),
    .QN(_00588_),
    .RESETN(net1408),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35883_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03640_),
    .QN(_00618_),
    .RESETN(net1409),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35884_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03641_),
    .QN(_00648_),
    .RESETN(net1410),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35885_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03642_),
    .QN(_00347_),
    .RESETN(net1411),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35886_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03643_),
    .QN(_00710_),
    .RESETN(net1412),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35887_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03644_),
    .QN(_00742_),
    .RESETN(net1413),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35888_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03645_),
    .QN(_00775_),
    .RESETN(net1414),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35889_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03646_),
    .QN(_00808_),
    .RESETN(net1415),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35890_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03647_),
    .QN(_00841_),
    .RESETN(net1416),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35891_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03648_),
    .QN(_00873_),
    .RESETN(net1417),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35892_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03649_),
    .QN(_00906_),
    .RESETN(net1418),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35893_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03650_),
    .QN(_00938_),
    .RESETN(net1419),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35894_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03651_),
    .QN(_00971_),
    .RESETN(net1420),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35895_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03652_),
    .QN(_01003_),
    .RESETN(net1421),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35896_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03653_),
    .QN(_01037_),
    .RESETN(net1422),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35897_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03654_),
    .QN(_01069_),
    .RESETN(net1423),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35898_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03655_),
    .QN(_01102_),
    .RESETN(net1424),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35899_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03656_),
    .QN(_01134_),
    .RESETN(net1425),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35900_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03657_),
    .QN(_01168_),
    .RESETN(net1426),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35901_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03658_),
    .QN(_01200_),
    .RESETN(net1427),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35902_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03659_),
    .QN(_01234_),
    .RESETN(net1428),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35903_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03660_),
    .QN(_01266_),
    .RESETN(net1429),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35904_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03661_),
    .QN(_01300_),
    .RESETN(net1430),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35905_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03662_),
    .QN(_00316_),
    .RESETN(net1431),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35906_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03663_),
    .QN(_00270_),
    .RESETN(net1432),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35907_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03664_),
    .QN(_00378_),
    .RESETN(net1433),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35908_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03665_),
    .QN(_00409_),
    .RESETN(net1434),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35909_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03666_),
    .QN(_00439_),
    .RESETN(net1435),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35910_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03667_),
    .QN(_00469_),
    .RESETN(net1436),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35911_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03668_),
    .QN(_00499_),
    .RESETN(net1437),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35912_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03669_),
    .QN(_00529_),
    .RESETN(net1438),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _35913_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03670_),
    .QN(_00559_),
    .RESETN(net1439),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35914_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03671_),
    .QN(_00589_),
    .RESETN(net1440),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35915_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03672_),
    .QN(_00619_),
    .RESETN(net1441),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35916_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03673_),
    .QN(_00649_),
    .RESETN(net1442),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35917_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03674_),
    .QN(_00348_),
    .RESETN(net1443),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35918_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03675_),
    .QN(_00711_),
    .RESETN(net1444),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35919_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03676_),
    .QN(_00743_),
    .RESETN(net1445),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35920_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03677_),
    .QN(_00776_),
    .RESETN(net1446),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35921_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03678_),
    .QN(_00809_),
    .RESETN(net1447),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35922_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03679_),
    .QN(_00842_),
    .RESETN(net1448),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35923_ (.CLK(clknet_level_3_1_27_clk_i),
    .D(_03680_),
    .QN(_00874_),
    .RESETN(net1449),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35924_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03681_),
    .QN(_00907_),
    .RESETN(net1450),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35925_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03682_),
    .QN(_00939_),
    .RESETN(net1451),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35926_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03683_),
    .QN(_00972_),
    .RESETN(net1452),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35927_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03684_),
    .QN(_01004_),
    .RESETN(net1453),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35928_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03685_),
    .QN(_01038_),
    .RESETN(net1454),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35929_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03686_),
    .QN(_01070_),
    .RESETN(net1455),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35930_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03687_),
    .QN(_01103_),
    .RESETN(net1456),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35931_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03688_),
    .QN(_01135_),
    .RESETN(net1457),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35932_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03689_),
    .QN(_01169_),
    .RESETN(net1458),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35933_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03690_),
    .QN(_01201_),
    .RESETN(net1459),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35934_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03691_),
    .QN(_01235_),
    .RESETN(net1460),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _35935_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03692_),
    .QN(_01267_),
    .RESETN(net1461),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35936_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03693_),
    .QN(_01301_),
    .RESETN(net1462),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _35937_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03694_),
    .QN(_00317_),
    .RESETN(net1463),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35938_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03695_),
    .QN(_00271_),
    .RESETN(net1464),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35939_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03696_),
    .QN(_00379_),
    .RESETN(net1465),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35940_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03697_),
    .QN(_00410_),
    .RESETN(net1466),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35941_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03698_),
    .QN(_00440_),
    .RESETN(net1467),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35942_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03699_),
    .QN(_00470_),
    .RESETN(net1468),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35943_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03700_),
    .QN(_00500_),
    .RESETN(net1469),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35944_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03701_),
    .QN(_00530_),
    .RESETN(net1470),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35945_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03702_),
    .QN(_00560_),
    .RESETN(net1471),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35946_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03703_),
    .QN(_00590_),
    .RESETN(net1472),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35947_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03704_),
    .QN(_00620_),
    .RESETN(net1473),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35948_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03705_),
    .QN(_00650_),
    .RESETN(net1474),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35949_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03706_),
    .QN(_00349_),
    .RESETN(net1475),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35950_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03707_),
    .QN(_00712_),
    .RESETN(net1476),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35951_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03708_),
    .QN(_00744_),
    .RESETN(net1477),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35952_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03709_),
    .QN(_00777_),
    .RESETN(net1478),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35953_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03710_),
    .QN(_00810_),
    .RESETN(net1479),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35954_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03711_),
    .QN(_00843_),
    .RESETN(net1480),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35955_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03712_),
    .QN(_00875_),
    .RESETN(net1481),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35956_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03713_),
    .QN(_00908_),
    .RESETN(net1482),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35957_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03714_),
    .QN(_00940_),
    .RESETN(net1483),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35958_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03715_),
    .QN(_00973_),
    .RESETN(net1484),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35959_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03716_),
    .QN(_01005_),
    .RESETN(net1485),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35960_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03717_),
    .QN(_01039_),
    .RESETN(net1486),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35961_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03718_),
    .QN(_01071_),
    .RESETN(net1487),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35962_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03719_),
    .QN(_01104_),
    .RESETN(net1488),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35963_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03720_),
    .QN(_01136_),
    .RESETN(net1489),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35964_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03721_),
    .QN(_01170_),
    .RESETN(net1490),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35965_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03722_),
    .QN(_01202_),
    .RESETN(net1491),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35966_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03723_),
    .QN(_01236_),
    .RESETN(net1492),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35967_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03724_),
    .QN(_01268_),
    .RESETN(net1493),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35968_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03725_),
    .QN(_01302_),
    .RESETN(net1494),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _35969_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03726_),
    .QN(_00318_),
    .RESETN(net1495),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _35970_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03727_),
    .QN(_00272_),
    .RESETN(net1496),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35971_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03728_),
    .QN(_00380_),
    .RESETN(net1497),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _35972_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03729_),
    .QN(_00411_),
    .RESETN(net1498),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _35973_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03730_),
    .QN(_00441_),
    .RESETN(net1499),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35974_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03731_),
    .QN(_00471_),
    .RESETN(net1500),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35975_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03732_),
    .QN(_00501_),
    .RESETN(net1501),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _35976_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03733_),
    .QN(_00531_),
    .RESETN(net1502),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _35977_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03734_),
    .QN(_00561_),
    .RESETN(net1503),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35978_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03735_),
    .QN(_00591_),
    .RESETN(net1504),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _35979_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03736_),
    .QN(_00621_),
    .RESETN(net1505),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35980_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03737_),
    .QN(_00651_),
    .RESETN(net1506),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _35981_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03738_),
    .QN(_00350_),
    .RESETN(net1507),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35982_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03739_),
    .QN(_00713_),
    .RESETN(net1508),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35983_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03740_),
    .QN(_00745_),
    .RESETN(net1509),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35984_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03741_),
    .QN(_00778_),
    .RESETN(net1510),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35985_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03742_),
    .QN(_00811_),
    .RESETN(net1511),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35986_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03743_),
    .QN(_00844_),
    .RESETN(net1512),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _35987_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03744_),
    .QN(_00876_),
    .RESETN(net1513),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35988_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03745_),
    .QN(_00909_),
    .RESETN(net1514),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35989_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03746_),
    .QN(_00941_),
    .RESETN(net1515),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35990_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03747_),
    .QN(_00974_),
    .RESETN(net1516),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _35991_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03748_),
    .QN(_01006_),
    .RESETN(net1517),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _35992_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03749_),
    .QN(_01040_),
    .RESETN(net1518),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35993_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03750_),
    .QN(_01072_),
    .RESETN(net1519),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _35994_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03751_),
    .QN(_01105_),
    .RESETN(net1520),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35995_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03752_),
    .QN(_01137_),
    .RESETN(net1521),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _35996_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03753_),
    .QN(_01171_),
    .RESETN(net1522),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _35997_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03754_),
    .QN(_01203_),
    .RESETN(net1523),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _35998_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03755_),
    .QN(_01237_),
    .RESETN(net1524),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _35999_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03756_),
    .QN(_01269_),
    .RESETN(net1525),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _36000_ (.CLK(clknet_level_3_1_28111_clk_i),
    .D(_03757_),
    .QN(_01303_),
    .RESETN(net1526),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36001_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03758_),
    .QN(_00319_),
    .RESETN(net1527),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36002_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03759_),
    .QN(_00273_),
    .RESETN(net1528),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36003_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03760_),
    .QN(_00381_),
    .RESETN(net1529),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36004_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03761_),
    .QN(_00412_),
    .RESETN(net1530),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36005_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03762_),
    .QN(_00442_),
    .RESETN(net1531),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36006_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03763_),
    .QN(_00472_),
    .RESETN(net1532),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36007_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03764_),
    .QN(_00502_),
    .RESETN(net1533),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36008_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03765_),
    .QN(_00532_),
    .RESETN(net1534),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36009_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03766_),
    .QN(_00562_),
    .RESETN(net1535),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36010_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03767_),
    .QN(_00592_),
    .RESETN(net1536),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36011_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03768_),
    .QN(_00622_),
    .RESETN(net1537),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36012_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03769_),
    .QN(_00652_),
    .RESETN(net1538),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36013_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03770_),
    .QN(_00351_),
    .RESETN(net1539),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36014_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03771_),
    .QN(_00714_),
    .RESETN(net1540),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36015_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03772_),
    .QN(_00746_),
    .RESETN(net1541),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36016_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03773_),
    .QN(_00779_),
    .RESETN(net1542),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36017_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03774_),
    .QN(_00812_),
    .RESETN(net1543),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36018_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03775_),
    .QN(_00845_),
    .RESETN(net1544),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36019_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03776_),
    .QN(_00877_),
    .RESETN(net1545),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36020_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03777_),
    .QN(_00910_),
    .RESETN(net1546),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36021_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03778_),
    .QN(_00942_),
    .RESETN(net1547),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36022_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03779_),
    .QN(_00975_),
    .RESETN(net1548),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36023_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03780_),
    .QN(_01007_),
    .RESETN(net1549),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36024_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03781_),
    .QN(_01041_),
    .RESETN(net1550),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36025_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03782_),
    .QN(_01073_),
    .RESETN(net1551),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36026_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03783_),
    .QN(_01106_),
    .RESETN(net1552),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36027_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03784_),
    .QN(_01138_),
    .RESETN(net1553),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36028_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03785_),
    .QN(_01172_),
    .RESETN(net1554),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36029_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03786_),
    .QN(_01204_),
    .RESETN(net1555),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36030_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03787_),
    .QN(_01238_),
    .RESETN(net1556),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36031_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03788_),
    .QN(_01270_),
    .RESETN(net1557),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36032_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03789_),
    .QN(_01304_),
    .RESETN(net1558),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36033_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03790_),
    .QN(_00320_),
    .RESETN(net1559),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36034_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03791_),
    .QN(_00274_),
    .RESETN(net1560),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36035_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03792_),
    .QN(_00382_),
    .RESETN(net1561),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36036_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03793_),
    .QN(_00413_),
    .RESETN(net1562),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _36037_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03794_),
    .QN(_00443_),
    .RESETN(net1563),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36038_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03795_),
    .QN(_00473_),
    .RESETN(net1564),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36039_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03796_),
    .QN(_00503_),
    .RESETN(net1565),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36040_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03797_),
    .QN(_00533_),
    .RESETN(net1566),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36041_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03798_),
    .QN(_00563_),
    .RESETN(net1567),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36042_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03799_),
    .QN(_00593_),
    .RESETN(net1568),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36043_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03800_),
    .QN(_00623_),
    .RESETN(net1569),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36044_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03801_),
    .QN(_00653_),
    .RESETN(net1570),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36045_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03802_),
    .QN(_00352_),
    .RESETN(net1571),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36046_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03803_),
    .QN(_00715_),
    .RESETN(net1572),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _36047_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03804_),
    .QN(_00747_),
    .RESETN(net1573),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36048_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03805_),
    .QN(_00780_),
    .RESETN(net1574),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _36049_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03806_),
    .QN(_00813_),
    .RESETN(net1575),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36050_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03807_),
    .QN(_00846_),
    .RESETN(net1576),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36051_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03808_),
    .QN(_00878_),
    .RESETN(net1577),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _36052_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03809_),
    .QN(_00911_),
    .RESETN(net1578),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36053_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03810_),
    .QN(_00943_),
    .RESETN(net1579),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36054_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03811_),
    .QN(_00976_),
    .RESETN(net1580),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36055_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03812_),
    .QN(_01008_),
    .RESETN(net1581),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36056_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03813_),
    .QN(_01042_),
    .RESETN(net1582),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36057_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03814_),
    .QN(_01074_),
    .RESETN(net1583),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36058_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03815_),
    .QN(_01107_),
    .RESETN(net1584),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36059_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03816_),
    .QN(_01139_),
    .RESETN(net1585),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36060_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03817_),
    .QN(_01173_),
    .RESETN(net1586),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36061_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03818_),
    .QN(_01205_),
    .RESETN(net1587),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36062_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03819_),
    .QN(_01239_),
    .RESETN(net1588),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36063_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03820_),
    .QN(_01271_),
    .RESETN(net1589),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36064_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03821_),
    .QN(_01305_),
    .RESETN(net1590),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36065_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03822_),
    .QN(_00321_),
    .RESETN(net1591),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36066_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03823_),
    .QN(_00275_),
    .RESETN(net1592),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36067_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03824_),
    .QN(_00383_),
    .RESETN(net1593),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36068_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03825_),
    .QN(_00414_),
    .RESETN(net1594),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36069_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03826_),
    .QN(_00444_),
    .RESETN(net1595),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36070_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03827_),
    .QN(_00474_),
    .RESETN(net1596),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36071_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03828_),
    .QN(_00504_),
    .RESETN(net1597),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36072_ (.CLK(clknet_level_3_1_1039_clk_i),
    .D(_03829_),
    .QN(_00534_),
    .RESETN(net1598),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36073_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03830_),
    .QN(_00564_),
    .RESETN(net1599),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36074_ (.CLK(clknet_level_3_1_935_clk_i),
    .D(_03831_),
    .QN(_00594_),
    .RESETN(net1600),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36075_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03832_),
    .QN(_00624_),
    .RESETN(net1601),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36076_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03833_),
    .QN(_00654_),
    .RESETN(net1602),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36077_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03834_),
    .QN(_00353_),
    .RESETN(net1603),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36078_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03835_),
    .QN(_00716_),
    .RESETN(net1604),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36079_ (.CLK(clknet_level_3_1_1559_clk_i),
    .D(_03836_),
    .QN(_00748_),
    .RESETN(net1605),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36080_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03837_),
    .QN(_00781_),
    .RESETN(net1606),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36081_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03838_),
    .QN(_00814_),
    .RESETN(net1607),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36082_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03839_),
    .QN(_00847_),
    .RESETN(net1608),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36083_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03840_),
    .QN(_00879_),
    .RESETN(net1609),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36084_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03841_),
    .QN(_00912_),
    .RESETN(net1610),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36085_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03842_),
    .QN(_00944_),
    .RESETN(net1611),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36086_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03843_),
    .QN(_00977_),
    .RESETN(net1612),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36087_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03844_),
    .QN(_01009_),
    .RESETN(net1613),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36088_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03845_),
    .QN(_01043_),
    .RESETN(net1614),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36089_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03846_),
    .QN(_01075_),
    .RESETN(net1615),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36090_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03847_),
    .QN(_01108_),
    .RESETN(net1616),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36091_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03848_),
    .QN(_01140_),
    .RESETN(net1617),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36092_ (.CLK(clknet_level_3_1_519_clk_i),
    .D(_03849_),
    .QN(_01174_),
    .RESETN(net1618),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36093_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03850_),
    .QN(_01206_),
    .RESETN(net1619),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36094_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03851_),
    .QN(_01240_),
    .RESETN(net1620),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36095_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03852_),
    .QN(_01272_),
    .RESETN(net1621),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36096_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03853_),
    .QN(_01306_),
    .RESETN(net1622),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36097_ (.CLK(clknet_level_3_1_29115_clk_i),
    .D(_03854_),
    .QN(_00322_),
    .RESETN(net1623),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36098_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03855_),
    .QN(_00276_),
    .RESETN(net1624),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36099_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03856_),
    .QN(_00384_),
    .RESETN(net1625),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36100_ (.CLK(clknet_level_3_1_30119_clk_i),
    .D(_03857_),
    .QN(_00415_),
    .RESETN(net1626),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _36101_ (.CLK(clknet_level_3_1_2391_clk_i),
    .D(_03858_),
    .QN(_00445_),
    .RESETN(net1627),
    .SETN(net440));
 DFFASRHQNx1_ASAP7_75t_R _36102_ (.CLK(clknet_level_3_1_2495_clk_i),
    .D(_03859_),
    .QN(_00475_),
    .RESETN(net1628),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36103_ (.CLK(clknet_level_3_1_26103_clk_i),
    .D(_03860_),
    .QN(_00505_),
    .RESETN(net1629),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36104_ (.CLK(clknet_level_3_1_1143_clk_i),
    .D(_03861_),
    .QN(_00535_),
    .RESETN(net1630),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36105_ (.CLK(clknet_level_3_1_1351_clk_i),
    .D(_03862_),
    .QN(_00565_),
    .RESETN(net1631),
    .SETN(net439));
 DFFASRHQNx1_ASAP7_75t_R _36106_ (.CLK(clknet_level_3_1_831_clk_i),
    .D(_03863_),
    .QN(_00595_),
    .RESETN(net1632),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36107_ (.CLK(clknet_level_3_1_2599_clk_i),
    .D(_03864_),
    .QN(_00625_),
    .RESETN(net1633),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36108_ (.CLK(clknet_level_3_1_1247_clk_i),
    .D(_03865_),
    .QN(_00655_),
    .RESETN(net1634),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36109_ (.CLK(clknet_level_3_1_2183_clk_i),
    .D(_03866_),
    .QN(_00354_),
    .RESETN(net1635),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36110_ (.CLK(clknet_level_3_1_415_clk_i),
    .D(_03867_),
    .QN(_00717_),
    .RESETN(net1636),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _36111_ (.CLK(clknet_level_3_1_1663_clk_i),
    .D(_03868_),
    .QN(_00749_),
    .RESETN(net1637),
    .SETN(net436));
 DFFASRHQNx1_ASAP7_75t_R _36112_ (.CLK(clknet_level_3_1_32127_clk_i),
    .D(_03869_),
    .QN(_00782_),
    .RESETN(net1638),
    .SETN(net443));
 DFFASRHQNx1_ASAP7_75t_R _36113_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03870_),
    .QN(_00815_),
    .RESETN(net1639),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36114_ (.CLK(clknet_level_3_1_1975_clk_i),
    .D(_03871_),
    .QN(_00848_),
    .RESETN(net1640),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36115_ (.CLK(clknet_level_3_1_13_clk_i),
    .D(_03872_),
    .QN(_00880_),
    .RESETN(net1641),
    .SETN(net445));
 DFFASRHQNx1_ASAP7_75t_R _36116_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03873_),
    .QN(_00913_),
    .RESETN(net1642),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36117_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03874_),
    .QN(_00945_),
    .RESETN(net1643),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36118_ (.CLK(clknet_level_3_1_2079_clk_i),
    .D(_03875_),
    .QN(_00978_),
    .RESETN(net1644),
    .SETN(net435));
 DFFASRHQNx1_ASAP7_75t_R _36119_ (.CLK(clknet_level_3_1_33131_clk_i),
    .D(_03876_),
    .QN(_01010_),
    .RESETN(net1645),
    .SETN(net442));
 DFFASRHQNx1_ASAP7_75t_R _36120_ (.CLK(clknet_level_3_1_1455_clk_i),
    .D(_03877_),
    .QN(_01044_),
    .RESETN(net1646),
    .SETN(net447));
 DFFASRHQNx1_ASAP7_75t_R _36121_ (.CLK(clknet_level_3_1_34135_clk_i),
    .D(_03878_),
    .QN(_01076_),
    .RESETN(net1647),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36122_ (.CLK(clknet_level_3_1_1871_clk_i),
    .D(_03879_),
    .QN(_01109_),
    .RESETN(net1648),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36123_ (.CLK(clknet_level_3_1_1767_clk_i),
    .D(_03880_),
    .QN(_01141_),
    .RESETN(net1649),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36124_ (.CLK(clknet_level_3_1_623_clk_i),
    .D(_03881_),
    .QN(_01175_),
    .RESETN(net1650),
    .SETN(net438));
 DFFASRHQNx1_ASAP7_75t_R _36125_ (.CLK(clknet_level_3_1_727_clk_i),
    .D(_03882_),
    .QN(_01207_),
    .RESETN(net1651),
    .SETN(net446));
 DFFASRHQNx1_ASAP7_75t_R _36126_ (.CLK(clknet_level_3_1_2287_clk_i),
    .D(_03883_),
    .QN(_01241_),
    .RESETN(net1652),
    .SETN(net437));
 DFFASRHQNx1_ASAP7_75t_R _36127_ (.CLK(clknet_level_3_1_311_clk_i),
    .D(_03884_),
    .QN(_01273_),
    .RESETN(net1653),
    .SETN(net444));
 DFFASRHQNx1_ASAP7_75t_R _36128_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(_03885_),
    .QN(_01307_),
    .RESETN(net1654),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36129_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03886_),
    .QN(_01519_),
    .RESETN(net1655),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36130_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03887_),
    .QN(_00659_),
    .RESETN(net1656),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36131_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03888_),
    .QN(_01518_),
    .RESETN(net1657),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36132_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03889_),
    .QN(_01517_),
    .RESETN(net1658),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36133_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03890_),
    .QN(_01516_),
    .RESETN(net1659),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36134_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03891_),
    .QN(_01515_),
    .RESETN(net1660),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36135_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03892_),
    .QN(_01514_),
    .RESETN(net1661),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36136_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03893_),
    .QN(_01513_),
    .RESETN(net1662),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36137_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03894_),
    .QN(_01512_),
    .RESETN(net1663),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36138_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03895_),
    .QN(_01511_),
    .RESETN(net1664),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36139_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03896_),
    .QN(_01510_),
    .RESETN(net1665),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36140_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03897_),
    .QN(_01509_),
    .RESETN(net1666),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36141_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03898_),
    .QN(_01508_),
    .RESETN(net1667),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36142_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03899_),
    .QN(_01507_),
    .RESETN(net1668),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36143_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03900_),
    .QN(_01506_),
    .RESETN(net1669),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36144_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03901_),
    .QN(_01505_),
    .RESETN(net1670),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36145_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03902_),
    .QN(_01504_),
    .RESETN(net1671),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36146_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03903_),
    .QN(_01503_),
    .RESETN(net1672),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36147_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03904_),
    .QN(_01502_),
    .RESETN(net1673),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36148_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03905_),
    .QN(_01501_),
    .RESETN(net1674),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36149_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03906_),
    .QN(_01500_),
    .RESETN(net1675),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36150_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03907_),
    .QN(_01499_),
    .RESETN(net1676),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36151_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03908_),
    .QN(_01498_),
    .RESETN(net1677),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36152_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03909_),
    .QN(_01497_),
    .RESETN(net1678),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36153_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03910_),
    .QN(_01496_),
    .RESETN(net1679),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36154_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03911_),
    .QN(_01495_),
    .RESETN(net1680),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36155_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03912_),
    .QN(_01494_),
    .RESETN(net1681),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36156_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03913_),
    .QN(_01493_),
    .RESETN(net1682),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36157_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03914_),
    .QN(_01492_),
    .RESETN(net1683),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36158_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_03915_),
    .QN(_01491_),
    .RESETN(net1684),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36159_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_03916_),
    .QN(_01490_),
    .RESETN(net1685),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36160_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03917_),
    .QN(_01489_),
    .RESETN(net1686),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36161_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_03918_),
    .QN(_01488_),
    .RESETN(net1687),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36162_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03919_),
    .QN(_00660_),
    .RESETN(net1688),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36163_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03920_),
    .QN(_01487_),
    .RESETN(net1689),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36164_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03921_),
    .QN(_01486_),
    .RESETN(net1690),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36165_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03922_),
    .QN(_01485_),
    .RESETN(net1691),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36166_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03923_),
    .QN(_01484_),
    .RESETN(net1692),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36167_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03924_),
    .QN(_01483_),
    .RESETN(net1693),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36168_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03925_),
    .QN(_01482_),
    .RESETN(net1694),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36169_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03926_),
    .QN(_01481_),
    .RESETN(net1695),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36170_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03927_),
    .QN(_01480_),
    .RESETN(net1696),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36171_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03928_),
    .QN(_01479_),
    .RESETN(net1697),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36172_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03929_),
    .QN(_01478_),
    .RESETN(net1698),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36173_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03930_),
    .QN(_01477_),
    .RESETN(net1699),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36174_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03931_),
    .QN(_01476_),
    .RESETN(net1700),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36175_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03932_),
    .QN(_01475_),
    .RESETN(net1701),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36176_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03933_),
    .QN(_01474_),
    .RESETN(net1702),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36177_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03934_),
    .QN(_01473_),
    .RESETN(net1703),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36178_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03935_),
    .QN(_01472_),
    .RESETN(net1704),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36179_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03936_),
    .QN(_01471_),
    .RESETN(net1705),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36180_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03937_),
    .QN(_01470_),
    .RESETN(net1706),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36181_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03938_),
    .QN(_01469_),
    .RESETN(net1707),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36182_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03939_),
    .QN(_01468_),
    .RESETN(net1708),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36183_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03940_),
    .QN(_01467_),
    .RESETN(net1709),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36184_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_03941_),
    .QN(_01466_),
    .RESETN(net1710),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36185_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03942_),
    .QN(_01465_),
    .RESETN(net1711),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36186_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_03943_),
    .QN(_01464_),
    .RESETN(net1712),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36187_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03944_),
    .QN(_01463_),
    .RESETN(net1713),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36188_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03945_),
    .QN(_01462_),
    .RESETN(net1714),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36189_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_03946_),
    .QN(_01461_),
    .RESETN(net1715),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36190_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03947_),
    .QN(_01460_),
    .RESETN(net1716),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36191_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03948_),
    .QN(_01459_),
    .RESETN(net1717),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36192_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_03949_),
    .QN(_01458_),
    .RESETN(net1718),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36193_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_03950_),
    .QN(_01457_),
    .RESETN(net1719),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36194_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_03951_),
    .QN(_01456_),
    .RESETN(net1720),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36195_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_03952_),
    .QN(_01455_),
    .RESETN(net1721),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36196_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_03953_),
    .QN(_01454_),
    .RESETN(net453),
    .SETN(net1722));
 DFFASRHQNx1_ASAP7_75t_R _36197_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_03954_),
    .QN(_01453_),
    .RESETN(net1723),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36198_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03955_),
    .QN(_01452_),
    .RESETN(net1724),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36199_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03956_),
    .QN(_01451_),
    .RESETN(net1725),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36200_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03957_),
    .QN(_01450_),
    .RESETN(net1726),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36201_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03958_),
    .QN(_01449_),
    .RESETN(net1727),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36202_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03959_),
    .QN(_01448_),
    .RESETN(net1728),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36203_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03960_),
    .QN(_01447_),
    .RESETN(net1729),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36204_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03961_),
    .QN(_01446_),
    .RESETN(net1730),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36205_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03962_),
    .QN(_01445_),
    .RESETN(net1731),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36206_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03963_),
    .QN(_01444_),
    .RESETN(net1732),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36207_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03964_),
    .QN(_01443_),
    .RESETN(net1733),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36208_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03965_),
    .QN(_01442_),
    .RESETN(net1734),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36209_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03966_),
    .QN(_01441_),
    .RESETN(net1735),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36210_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03967_),
    .QN(_02221_),
    .RESETN(net1736),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36211_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03968_),
    .QN(_02220_),
    .RESETN(net1737),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36212_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03969_),
    .QN(_02219_),
    .RESETN(net1738),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36213_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03970_),
    .QN(_02218_),
    .RESETN(net1739),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36214_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03971_),
    .QN(_02217_),
    .RESETN(net1740),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36215_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03972_),
    .QN(_02216_),
    .RESETN(net1741),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36216_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03973_),
    .QN(_02215_),
    .RESETN(net1742),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36217_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03974_),
    .QN(_02214_),
    .RESETN(net1743),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36218_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03975_),
    .QN(_02213_),
    .RESETN(net1744),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36219_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03976_),
    .QN(_02212_),
    .RESETN(net1745),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36220_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03977_),
    .QN(_02211_),
    .RESETN(net1746),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36221_ (.CLK(\clknet_leaf_4_core_clock_gate_i.clk_o ),
    .D(_03978_),
    .QN(_02210_),
    .RESETN(net1747),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36222_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03979_),
    .QN(_02209_),
    .RESETN(net1748),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36223_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03980_),
    .QN(_02208_),
    .RESETN(net1749),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36224_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03981_),
    .QN(_02207_),
    .RESETN(net1750),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36225_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_03982_),
    .QN(_02206_),
    .RESETN(net1751),
    .SETN(net451));
 DFFASRHQNx1_ASAP7_75t_R _36226_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03983_),
    .QN(_02205_),
    .RESETN(net1752),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36227_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_03984_),
    .QN(_02204_),
    .RESETN(net1753),
    .SETN(net448));
 DFFASRHQNx1_ASAP7_75t_R _36228_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03985_),
    .QN(_02203_),
    .RESETN(net1754),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36229_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_03986_),
    .QN(_02202_),
    .RESETN(net1755),
    .SETN(net450));
 DFFHQNx1_ASAP7_75t_R _36230_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03987_),
    .QN(_02201_));
 DFFHQNx1_ASAP7_75t_R _36231_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03988_),
    .QN(_02200_));
 DFFHQNx1_ASAP7_75t_R _36232_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03989_),
    .QN(_02199_));
 DFFHQNx1_ASAP7_75t_R _36233_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03990_),
    .QN(_02198_));
 DFFHQNx1_ASAP7_75t_R _36234_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03991_),
    .QN(_02197_));
 DFFHQNx1_ASAP7_75t_R _36235_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03992_),
    .QN(_02196_));
 DFFHQNx1_ASAP7_75t_R _36236_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03993_),
    .QN(_02195_));
 DFFHQNx1_ASAP7_75t_R _36237_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_03994_),
    .QN(_02194_));
 DFFHQNx1_ASAP7_75t_R _36238_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03995_),
    .QN(_02193_));
 DFFHQNx1_ASAP7_75t_R _36239_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03996_),
    .QN(_02192_));
 DFFHQNx1_ASAP7_75t_R _36240_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03997_),
    .QN(_02191_));
 DFFHQNx1_ASAP7_75t_R _36241_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03998_),
    .QN(_02190_));
 DFFHQNx1_ASAP7_75t_R _36242_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_03999_),
    .QN(_02189_));
 DFFHQNx1_ASAP7_75t_R _36243_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04000_),
    .QN(_02188_));
 DFFHQNx1_ASAP7_75t_R _36244_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04001_),
    .QN(_02187_));
 DFFHQNx1_ASAP7_75t_R _36245_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04002_),
    .QN(_02186_));
 DFFHQNx1_ASAP7_75t_R _36246_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04003_),
    .QN(_02185_));
 DFFHQNx1_ASAP7_75t_R _36247_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04004_),
    .QN(_02184_));
 DFFHQNx1_ASAP7_75t_R _36248_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04005_),
    .QN(_02183_));
 DFFHQNx1_ASAP7_75t_R _36249_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04006_),
    .QN(_02182_));
 DFFHQNx1_ASAP7_75t_R _36250_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04007_),
    .QN(_02181_));
 DFFHQNx1_ASAP7_75t_R _36251_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04008_),
    .QN(_02180_));
 DFFHQNx1_ASAP7_75t_R _36252_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04009_),
    .QN(_02179_));
 DFFHQNx1_ASAP7_75t_R _36253_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04010_),
    .QN(_02178_));
 DFFHQNx1_ASAP7_75t_R _36254_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04011_),
    .QN(_02177_));
 DFFHQNx1_ASAP7_75t_R _36255_ (.CLK(\clknet_leaf_22_core_clock_gate_i.clk_o ),
    .D(_04012_),
    .QN(_02176_));
 DFFHQNx1_ASAP7_75t_R _36256_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04013_),
    .QN(_02175_));
 DFFHQNx1_ASAP7_75t_R _36257_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04014_),
    .QN(_02174_));
 DFFHQNx1_ASAP7_75t_R _36258_ (.CLK(\clknet_leaf_20_core_clock_gate_i.clk_o ),
    .D(_04015_),
    .QN(_02173_));
 DFFHQNx1_ASAP7_75t_R _36259_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(_04016_),
    .QN(_01729_));
 DFFASRHQNx1_ASAP7_75t_R _36260_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_00006_),
    .QN(_01730_),
    .RESETN(net1756),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36261_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(_00007_),
    .QN(_01731_),
    .RESETN(net1757),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36262_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_00000_),
    .QN(_01732_),
    .RESETN(net452),
    .SETN(net1758));
 DFFASRHQNx1_ASAP7_75t_R _36263_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_00001_),
    .QN(_01314_),
    .RESETN(net1759),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36264_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04017_),
    .QN(_02172_),
    .RESETN(net1760),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36265_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04018_),
    .QN(_02171_),
    .RESETN(net1761),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36266_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04019_),
    .QN(_02170_),
    .RESETN(net1762),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36267_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04020_),
    .QN(_02169_),
    .RESETN(net1763),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36268_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04021_),
    .QN(_02168_),
    .RESETN(net1764),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36269_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04022_),
    .QN(_02167_),
    .RESETN(net1765),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36270_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04023_),
    .QN(_02166_),
    .RESETN(net1766),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36271_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04024_),
    .QN(_02165_),
    .RESETN(net1767),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36272_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04025_),
    .QN(_02164_),
    .RESETN(net1768),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36273_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04026_),
    .QN(_02163_),
    .RESETN(net1769),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36274_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04027_),
    .QN(_02162_),
    .RESETN(net1770),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36275_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04028_),
    .QN(_02161_),
    .RESETN(net1771),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36276_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04029_),
    .QN(_02160_),
    .RESETN(net1772),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36277_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04030_),
    .QN(_02159_),
    .RESETN(net1773),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36278_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04031_),
    .QN(_02158_),
    .RESETN(net1774),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36279_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04032_),
    .QN(_02157_),
    .RESETN(net1775),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36280_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04033_),
    .QN(_02156_),
    .RESETN(net1776),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36281_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04034_),
    .QN(_02155_),
    .RESETN(net1777),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36282_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04035_),
    .QN(_02154_),
    .RESETN(net1778),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36283_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04036_),
    .QN(_02153_),
    .RESETN(net1779),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36284_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04037_),
    .QN(_02152_),
    .RESETN(net1780),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36285_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04038_),
    .QN(_02151_),
    .RESETN(net1781),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36286_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04039_),
    .QN(_02150_),
    .RESETN(net1782),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36287_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04040_),
    .QN(_02149_),
    .RESETN(net1783),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36288_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04041_),
    .QN(_02148_),
    .RESETN(net1784),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36289_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04042_),
    .QN(_02147_),
    .RESETN(net1785),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36290_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04043_),
    .QN(_02146_),
    .RESETN(net1786),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36291_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04044_),
    .QN(_02145_),
    .RESETN(net1787),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36292_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04045_),
    .QN(_02144_),
    .RESETN(net1788),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36293_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04046_),
    .QN(_02143_),
    .RESETN(net1789),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36294_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04047_),
    .QN(_02142_),
    .RESETN(net1790),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36295_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04048_),
    .QN(_02141_),
    .RESETN(net1791),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36296_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04049_),
    .QN(_02140_),
    .RESETN(net457),
    .SETN(net1792));
 DFFASRHQNx1_ASAP7_75t_R _36297_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04050_),
    .QN(_17810_),
    .RESETN(net457),
    .SETN(net1793));
 DFFASRHQNx1_ASAP7_75t_R _36298_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04051_),
    .QN(_02139_),
    .RESETN(net1794),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36299_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04052_),
    .QN(_02138_),
    .RESETN(net1795),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36300_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04053_),
    .QN(_02137_),
    .RESETN(net1796),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36301_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04054_),
    .QN(_02136_),
    .RESETN(net1797),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36302_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04055_),
    .QN(_02135_),
    .RESETN(net1798),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36303_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04056_),
    .QN(_02134_),
    .RESETN(net1799),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36304_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04057_),
    .QN(_02133_),
    .RESETN(net1800),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36305_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04058_),
    .QN(_02132_),
    .RESETN(net1801),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36306_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04059_),
    .QN(_02131_),
    .RESETN(net1802),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36307_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04060_),
    .QN(_02130_),
    .RESETN(net1803),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36308_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04061_),
    .QN(_02129_),
    .RESETN(net1804),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36309_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04062_),
    .QN(_02128_),
    .RESETN(net1805),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36310_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04063_),
    .QN(_02127_),
    .RESETN(net1806),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36311_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04064_),
    .QN(_02126_),
    .RESETN(net1807),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36312_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04065_),
    .QN(_02125_),
    .RESETN(net1808),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36313_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04066_),
    .QN(_02124_),
    .RESETN(net1809),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36314_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04067_),
    .QN(_02123_),
    .RESETN(net1810),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36315_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04068_),
    .QN(_02122_),
    .RESETN(net1811),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36316_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04069_),
    .QN(_02121_),
    .RESETN(net1812),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36317_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04070_),
    .QN(_02120_),
    .RESETN(net1813),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36318_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04071_),
    .QN(_02119_),
    .RESETN(net1814),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36319_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04072_),
    .QN(_02118_),
    .RESETN(net1815),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36320_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04073_),
    .QN(_02117_),
    .RESETN(net1816),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36321_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04074_),
    .QN(_02116_),
    .RESETN(net1817),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36322_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04075_),
    .QN(_02115_),
    .RESETN(net1818),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36323_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04076_),
    .QN(_02114_),
    .RESETN(net1819),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36324_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04077_),
    .QN(_02113_),
    .RESETN(net1820),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36325_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04078_),
    .QN(_02112_),
    .RESETN(net1821),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36326_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04079_),
    .QN(_02111_),
    .RESETN(net1822),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36327_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04080_),
    .QN(_02110_),
    .RESETN(net1823),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36328_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04081_),
    .QN(_02109_),
    .RESETN(net1824),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36329_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04082_),
    .QN(_02108_),
    .RESETN(net1825),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36330_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04083_),
    .QN(_02107_),
    .RESETN(net1826),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36331_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04084_),
    .QN(_02106_),
    .RESETN(net1827),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36332_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04085_),
    .QN(_02105_),
    .RESETN(net453),
    .SETN(net1828));
 DFFASRHQNx1_ASAP7_75t_R _36333_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04086_),
    .QN(_02104_),
    .RESETN(net1829),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36334_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04087_),
    .QN(_02103_),
    .RESETN(net1830),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36335_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04088_),
    .QN(_02102_),
    .RESETN(net1831),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36336_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04089_),
    .QN(_02101_),
    .RESETN(net1832),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36337_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04090_),
    .QN(_02100_),
    .RESETN(net1833),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36338_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04091_),
    .QN(_02099_),
    .RESETN(net1834),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36339_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04092_),
    .QN(_02098_),
    .RESETN(net1835),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36340_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(net3648),
    .QN(_02097_),
    .RESETN(net1836),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36341_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04094_),
    .QN(_02096_),
    .RESETN(net1837),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36342_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04095_),
    .QN(_02095_),
    .RESETN(net1838),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36343_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(net3380),
    .QN(_02094_),
    .RESETN(net1839),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36344_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04097_),
    .QN(_02093_),
    .RESETN(net1840),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36345_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04098_),
    .QN(_02092_),
    .RESETN(net1841),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36346_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04099_),
    .QN(_02091_),
    .RESETN(net1842),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36347_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04100_),
    .QN(_02090_),
    .RESETN(net1843),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36348_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04101_),
    .QN(_02089_),
    .RESETN(net1844),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36349_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04102_),
    .QN(_02088_),
    .RESETN(net1845),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36350_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04103_),
    .QN(_02087_),
    .RESETN(net1846),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36351_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04104_),
    .QN(_02086_),
    .RESETN(net1847),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36352_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04105_),
    .QN(_02085_),
    .RESETN(net1848),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36353_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04106_),
    .QN(_02084_),
    .RESETN(net1849),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36354_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04107_),
    .QN(_02083_),
    .RESETN(net1850),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36355_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04108_),
    .QN(_02082_),
    .RESETN(net1851),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36356_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04109_),
    .QN(_02081_),
    .RESETN(net1852),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36357_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04110_),
    .QN(_02080_),
    .RESETN(net1853),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36358_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04111_),
    .QN(_02079_),
    .RESETN(net1854),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36359_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04112_),
    .QN(_02078_),
    .RESETN(net1855),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36360_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04113_),
    .QN(_02077_),
    .RESETN(net1856),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36361_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04114_),
    .QN(_02076_),
    .RESETN(net1857),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36362_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04115_),
    .QN(_02075_),
    .RESETN(net1858),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36363_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04116_),
    .QN(_02074_),
    .RESETN(net1859),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36364_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04117_),
    .QN(_02073_),
    .RESETN(net1860),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36365_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04118_),
    .QN(_02072_),
    .RESETN(net1861),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36366_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04119_),
    .QN(_02071_),
    .RESETN(net1862),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36367_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04120_),
    .QN(_02070_),
    .RESETN(net1863),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36368_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04121_),
    .QN(_02069_),
    .RESETN(net1864),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36369_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04122_),
    .QN(_02068_),
    .RESETN(net1865),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36370_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04123_),
    .QN(_02067_),
    .RESETN(net1866),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36371_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04124_),
    .QN(_00095_),
    .RESETN(net1867),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36372_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04125_),
    .QN(_00098_),
    .RESETN(net1868),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36373_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04126_),
    .QN(_00101_),
    .RESETN(net1869),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36374_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04127_),
    .QN(_00657_),
    .RESETN(net1870),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36375_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04128_),
    .QN(_00656_),
    .RESETN(net1871),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36376_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04129_),
    .QN(_00108_),
    .RESETN(net1872),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36377_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04130_),
    .QN(_00111_),
    .RESETN(net1873),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36378_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04131_),
    .QN(_00114_),
    .RESETN(net1874),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36379_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04132_),
    .QN(_00117_),
    .RESETN(net1875),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36380_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04133_),
    .QN(_00120_),
    .RESETN(net1876),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36381_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04134_),
    .QN(_00123_),
    .RESETN(net1877),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36382_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04135_),
    .QN(_00126_),
    .RESETN(net1878),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36383_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04136_),
    .QN(_00129_),
    .RESETN(net1879),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36384_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04137_),
    .QN(_00132_),
    .RESETN(net1880),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36385_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04138_),
    .QN(_00135_),
    .RESETN(net1881),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36386_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04139_),
    .QN(_00138_),
    .RESETN(net1882),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36387_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04140_),
    .QN(_00141_),
    .RESETN(net1883),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36388_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04141_),
    .QN(_00144_),
    .RESETN(net1884),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36389_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04142_),
    .QN(_00147_),
    .RESETN(net1885),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36390_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04143_),
    .QN(_00150_),
    .RESETN(net1886),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36391_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04144_),
    .QN(_00153_),
    .RESETN(net1887),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36392_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04145_),
    .QN(_00156_),
    .RESETN(net1888),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36393_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04146_),
    .QN(_00159_),
    .RESETN(net1889),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36394_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04147_),
    .QN(_00161_),
    .RESETN(net1890),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36395_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04148_),
    .QN(_02066_),
    .RESETN(net1891),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36396_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04149_),
    .QN(_02065_),
    .RESETN(net1892),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36397_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04150_),
    .QN(_02064_),
    .RESETN(net1893),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36398_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04151_),
    .QN(_02063_),
    .RESETN(net1894),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36399_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04152_),
    .QN(_02062_),
    .RESETN(net1895),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36400_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04153_),
    .QN(_02061_),
    .RESETN(net1896),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36401_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04154_),
    .QN(_02060_),
    .RESETN(net1897),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36402_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04155_),
    .QN(_02059_),
    .RESETN(net1898),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36403_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04156_),
    .QN(_02058_),
    .RESETN(net1899),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36404_ (.CLK(\clknet_leaf_7_core_clock_gate_i.clk_o ),
    .D(_04157_),
    .QN(_02057_),
    .RESETN(net1900),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36405_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04158_),
    .QN(_02056_),
    .RESETN(net1901),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36406_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04159_),
    .QN(_02055_),
    .RESETN(net1902),
    .SETN(net2385));
 DFFASRHQNx1_ASAP7_75t_R _36407_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04160_),
    .QN(_02054_),
    .RESETN(net1903),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36408_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04161_),
    .QN(_02053_),
    .RESETN(net1904),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36409_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04162_),
    .QN(_02052_),
    .RESETN(net1905),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36410_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04163_),
    .QN(_02051_),
    .RESETN(net1906),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36411_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04164_),
    .QN(_02050_),
    .RESETN(net1907),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36412_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04165_),
    .QN(_02049_),
    .RESETN(net1908),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36413_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04166_),
    .QN(_02048_),
    .RESETN(net1909),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36414_ (.CLK(\clknet_leaf_8_core_clock_gate_i.clk_o ),
    .D(_04167_),
    .QN(_02047_),
    .RESETN(net1910),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36415_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04168_),
    .QN(_02046_),
    .RESETN(net1911),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36416_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04169_),
    .QN(_02045_),
    .RESETN(net1912),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36417_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04170_),
    .QN(_02044_),
    .RESETN(net1913),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36418_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04171_),
    .QN(_02043_),
    .RESETN(net1914),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36419_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04172_),
    .QN(_02042_),
    .RESETN(net1915),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36420_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04173_),
    .QN(_02041_),
    .RESETN(net1916),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36421_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04174_),
    .QN(_02040_),
    .RESETN(net1917),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36422_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04175_),
    .QN(_02039_),
    .RESETN(net1918),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36423_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04176_),
    .QN(_02038_),
    .RESETN(net1919),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36424_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04177_),
    .QN(_02037_),
    .RESETN(net1920),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36425_ (.CLK(\clknet_leaf_9_core_clock_gate_i.clk_o ),
    .D(_04178_),
    .QN(_02036_),
    .RESETN(net1921),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36426_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04179_),
    .QN(_02035_),
    .RESETN(net1922),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36427_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04180_),
    .QN(_02034_),
    .RESETN(net1923),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36428_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04181_),
    .QN(_02033_),
    .RESETN(net1924),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36429_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04182_),
    .QN(_02032_),
    .RESETN(net1925),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36430_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04183_),
    .QN(_02031_),
    .RESETN(net1926),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36431_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04184_),
    .QN(_02030_),
    .RESETN(net1927),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36432_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04185_),
    .QN(_02029_),
    .RESETN(net1928),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36433_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04186_),
    .QN(_02028_),
    .RESETN(net1929),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36434_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04187_),
    .QN(_02027_),
    .RESETN(net1930),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36435_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04188_),
    .QN(_02026_),
    .RESETN(net1931),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36436_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04189_),
    .QN(_02025_),
    .RESETN(net1932),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36437_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04190_),
    .QN(_02024_),
    .RESETN(net1933),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36438_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04191_),
    .QN(_02023_),
    .RESETN(net1934),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36439_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04192_),
    .QN(_02022_),
    .RESETN(net1935),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36440_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04193_),
    .QN(_02021_),
    .RESETN(net1936),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36441_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04194_),
    .QN(_02020_),
    .RESETN(net1937),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36442_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04195_),
    .QN(_02019_),
    .RESETN(net1938),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36443_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04196_),
    .QN(_02018_),
    .RESETN(net1939),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36444_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04197_),
    .QN(_02017_),
    .RESETN(net1940),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36445_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04198_),
    .QN(_02016_),
    .RESETN(net1941),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36446_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04199_),
    .QN(_02015_),
    .RESETN(net1942),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36447_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04200_),
    .QN(_02014_),
    .RESETN(net1943),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36448_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04201_),
    .QN(_02013_),
    .RESETN(net1944),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36449_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04202_),
    .QN(_02012_),
    .RESETN(net1945),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36450_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04203_),
    .QN(_02011_),
    .RESETN(net1946),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36451_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04204_),
    .QN(_02010_),
    .RESETN(net1947),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36452_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04205_),
    .QN(_02009_),
    .RESETN(net1948),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36453_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04206_),
    .QN(_02008_),
    .RESETN(net1949),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36454_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04207_),
    .QN(_02007_),
    .RESETN(net1950),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36455_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(net3582),
    .QN(_02006_),
    .RESETN(net1951),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36456_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04209_),
    .QN(_02005_),
    .RESETN(net1952),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36457_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(net3640),
    .QN(_02004_),
    .RESETN(net1953),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36458_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04211_),
    .QN(_02003_),
    .RESETN(net1954),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36459_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04212_),
    .QN(_02002_),
    .RESETN(net1955),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36460_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04213_),
    .QN(_02001_),
    .RESETN(net1956),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36461_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04214_),
    .QN(_02000_),
    .RESETN(net1957),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36462_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04215_),
    .QN(_01999_),
    .RESETN(net1958),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36463_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04216_),
    .QN(_01998_),
    .RESETN(net1959),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36464_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04217_),
    .QN(_01997_),
    .RESETN(net1960),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36465_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04218_),
    .QN(_01996_),
    .RESETN(net1961),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36466_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04219_),
    .QN(_01995_),
    .RESETN(net1962),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36467_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04220_),
    .QN(_01994_),
    .RESETN(net1963),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36468_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04221_),
    .QN(_01993_),
    .RESETN(net1964),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36469_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04222_),
    .QN(_01992_),
    .RESETN(net1965),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36470_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04223_),
    .QN(_01991_),
    .RESETN(net1966),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36471_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04224_),
    .QN(_01990_),
    .RESETN(net1967),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36472_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04225_),
    .QN(_01989_),
    .RESETN(net1968),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36473_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04226_),
    .QN(_01988_),
    .RESETN(net1969),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36474_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04227_),
    .QN(_01987_),
    .RESETN(net1970),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36475_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04228_),
    .QN(_01986_),
    .RESETN(net1971),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36476_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04229_),
    .QN(_01985_),
    .RESETN(net1972),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36477_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04230_),
    .QN(_01984_),
    .RESETN(net1973),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36478_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04231_),
    .QN(_01983_),
    .RESETN(net1974),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36479_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04232_),
    .QN(_01982_),
    .RESETN(net1975),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36480_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04233_),
    .QN(_01981_),
    .RESETN(net1976),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36481_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04234_),
    .QN(_01980_),
    .RESETN(net1977),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36482_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04235_),
    .QN(_01979_),
    .RESETN(net1978),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36483_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04236_),
    .QN(_01978_),
    .RESETN(net1979),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36484_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04237_),
    .QN(_01977_),
    .RESETN(net1980),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36485_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04238_),
    .QN(_01976_),
    .RESETN(net1981),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36486_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04239_),
    .QN(_01975_),
    .RESETN(net1982),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36487_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04240_),
    .QN(_01974_),
    .RESETN(net1983),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36488_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04241_),
    .QN(_01973_),
    .RESETN(net1984),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36489_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04242_),
    .QN(_01972_),
    .RESETN(net1985),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36490_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04243_),
    .QN(_01971_),
    .RESETN(net1986),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36491_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04244_),
    .QN(_01970_),
    .RESETN(net1987),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36492_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04245_),
    .QN(_01969_),
    .RESETN(net1988),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36493_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04246_),
    .QN(_01968_),
    .RESETN(net1989),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36494_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04247_),
    .QN(_01967_),
    .RESETN(net1990),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36495_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04248_),
    .QN(_01966_),
    .RESETN(net1991),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36496_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04249_),
    .QN(_01965_),
    .RESETN(net1992),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36497_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04250_),
    .QN(_01964_),
    .RESETN(net1993),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36498_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(net3605),
    .QN(_01963_),
    .RESETN(net1994),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36499_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(net3661),
    .QN(_01962_),
    .RESETN(net1995),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36500_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(net3558),
    .QN(_01961_),
    .RESETN(net1996),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36501_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(net3712),
    .QN(_01960_),
    .RESETN(net1997),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36502_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04255_),
    .QN(_01959_),
    .RESETN(net1998),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36503_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04256_),
    .QN(_01958_),
    .RESETN(net1999),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36504_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04257_),
    .QN(_01957_),
    .RESETN(net2000),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36505_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04258_),
    .QN(_01956_),
    .RESETN(net2001),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36506_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04259_),
    .QN(_01955_),
    .RESETN(net2002),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36507_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04260_),
    .QN(_01954_),
    .RESETN(net2003),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36508_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(_04261_),
    .QN(_01953_),
    .RESETN(net2004),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36509_ (.CLK(\clknet_leaf_10_core_clock_gate_i.clk_o ),
    .D(net3595),
    .QN(_01952_),
    .RESETN(net2005),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36510_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04263_),
    .QN(_01951_),
    .RESETN(net2006),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36511_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04264_),
    .QN(_01950_),
    .RESETN(net2007),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36512_ (.CLK(\clknet_leaf_11_core_clock_gate_i.clk_o ),
    .D(_04265_),
    .QN(_01949_),
    .RESETN(net2008),
    .SETN(net459));
 DFFASRHQNx1_ASAP7_75t_R _36513_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(_04266_),
    .QN(_01948_),
    .RESETN(net2009),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36514_ (.CLK(\clknet_leaf_12_core_clock_gate_i.clk_o ),
    .D(net3655),
    .QN(_01947_),
    .RESETN(net2010),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36515_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(net3545),
    .QN(_01946_),
    .RESETN(net2011),
    .SETN(net458));
 DFFASRHQNx1_ASAP7_75t_R _36516_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04269_),
    .QN(_01945_),
    .RESETN(net2012),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36517_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04270_),
    .QN(_01944_),
    .RESETN(net2013),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36518_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04271_),
    .QN(_01943_),
    .RESETN(net2014),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36519_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04272_),
    .QN(_01942_),
    .RESETN(net2015),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36520_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04273_),
    .QN(_01941_),
    .RESETN(net2016),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36521_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04274_),
    .QN(_01940_),
    .RESETN(net2017),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36522_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04275_),
    .QN(_01939_),
    .RESETN(net2018),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36523_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04276_),
    .QN(_01938_),
    .RESETN(net2019),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36524_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04277_),
    .QN(_01937_),
    .RESETN(net2020),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36525_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04278_),
    .QN(_01936_),
    .RESETN(net2021),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36526_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04279_),
    .QN(_01935_),
    .RESETN(net2022),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36527_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04280_),
    .QN(_01934_),
    .RESETN(net2023),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36528_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04281_),
    .QN(_01933_),
    .RESETN(net2024),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36529_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04282_),
    .QN(_01932_),
    .RESETN(net2025),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36530_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04283_),
    .QN(_01931_),
    .RESETN(net2026),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36531_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04284_),
    .QN(_01930_),
    .RESETN(net2027),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36532_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04285_),
    .QN(_01929_),
    .RESETN(net2028),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36533_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04286_),
    .QN(_01928_),
    .RESETN(net2029),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36534_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04287_),
    .QN(_01927_),
    .RESETN(net2030),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36535_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04288_),
    .QN(_01926_),
    .RESETN(net2031),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36536_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04289_),
    .QN(_01925_),
    .RESETN(net2032),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36537_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04290_),
    .QN(_01924_),
    .RESETN(net2033),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36538_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04291_),
    .QN(_01923_),
    .RESETN(net2034),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36539_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04292_),
    .QN(_01922_),
    .RESETN(net2035),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36540_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04293_),
    .QN(_01921_),
    .RESETN(net2036),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36541_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04294_),
    .QN(_01920_),
    .RESETN(net2037),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36542_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04295_),
    .QN(_01919_),
    .RESETN(net2038),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36543_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04296_),
    .QN(_01918_),
    .RESETN(net2039),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36544_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04297_),
    .QN(_01917_),
    .RESETN(net2040),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36545_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04298_),
    .QN(_01916_),
    .RESETN(net2041),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36546_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04299_),
    .QN(_01915_),
    .RESETN(net2042),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36547_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04300_),
    .QN(_01914_),
    .RESETN(net2043),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36548_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(net3519),
    .QN(_01913_),
    .RESETN(net2044),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36549_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04302_),
    .QN(_01912_),
    .RESETN(net2045),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36550_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04303_),
    .QN(_01911_),
    .RESETN(net2046),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36551_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04304_),
    .QN(_01910_),
    .RESETN(net2047),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36552_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04305_),
    .QN(_01909_),
    .RESETN(net2048),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36553_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04306_),
    .QN(_01908_),
    .RESETN(net2049),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36554_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04307_),
    .QN(_01907_),
    .RESETN(net2050),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36555_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04308_),
    .QN(_01906_),
    .RESETN(net2051),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36556_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04309_),
    .QN(_01905_),
    .RESETN(net2052),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36557_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04310_),
    .QN(_01904_),
    .RESETN(net2053),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36558_ (.CLK(\clknet_leaf_13_core_clock_gate_i.clk_o ),
    .D(_04311_),
    .QN(_01903_),
    .RESETN(net2054),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36559_ (.CLK(\clknet_leaf_14_core_clock_gate_i.clk_o ),
    .D(_04312_),
    .QN(_01902_),
    .RESETN(net2055),
    .SETN(net453));
 DFFASRHQNx1_ASAP7_75t_R _36560_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04313_),
    .QN(_01901_),
    .RESETN(net2056),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36561_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04314_),
    .QN(_01900_),
    .RESETN(net2057),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36562_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04315_),
    .QN(_01899_),
    .RESETN(net2058),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36563_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04316_),
    .QN(_01898_),
    .RESETN(net2059),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36564_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04317_),
    .QN(_01897_),
    .RESETN(net2060),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36565_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04318_),
    .QN(_01896_),
    .RESETN(net2061),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36566_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04319_),
    .QN(_01895_),
    .RESETN(net2062),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36567_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04320_),
    .QN(_01894_),
    .RESETN(net2063),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36568_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04321_),
    .QN(_01893_),
    .RESETN(net2064),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36569_ (.CLK(\clknet_leaf_21_core_clock_gate_i.clk_o ),
    .D(_04322_),
    .QN(_01892_),
    .RESETN(net2065),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36570_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04323_),
    .QN(_01891_),
    .RESETN(net2066),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36571_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04324_),
    .QN(_01890_),
    .RESETN(net2067),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36572_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04325_),
    .QN(_01889_),
    .RESETN(net2068),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36573_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04326_),
    .QN(_01888_),
    .RESETN(net2069),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36574_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04327_),
    .QN(_01887_),
    .RESETN(net2070),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36575_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04328_),
    .QN(_01886_),
    .RESETN(net2071),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36576_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04329_),
    .QN(_01885_),
    .RESETN(net2072),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36577_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04330_),
    .QN(_01884_),
    .RESETN(net2073),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36578_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04331_),
    .QN(_01883_),
    .RESETN(net2074),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36579_ (.CLK(\clknet_leaf_18_core_clock_gate_i.clk_o ),
    .D(_04332_),
    .QN(_01882_),
    .RESETN(net2075),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36580_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04333_),
    .QN(_01881_),
    .RESETN(net2076),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36581_ (.CLK(\clknet_leaf_17_core_clock_gate_i.clk_o ),
    .D(_04334_),
    .QN(_01880_),
    .RESETN(net2077),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36582_ (.CLK(\clknet_leaf_19_core_clock_gate_i.clk_o ),
    .D(_04335_),
    .QN(_01879_),
    .RESETN(net2078),
    .SETN(net455));
 DFFASRHQNx1_ASAP7_75t_R _36583_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04336_),
    .QN(_01878_),
    .RESETN(net2079),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36584_ (.CLK(\clknet_leaf_16_core_clock_gate_i.clk_o ),
    .D(_04337_),
    .QN(_01877_),
    .RESETN(net2080),
    .SETN(net456));
 DFFASRHQNx1_ASAP7_75t_R _36585_ (.CLK(\clknet_leaf_15_core_clock_gate_i.clk_o ),
    .D(_04338_),
    .QN(_01876_),
    .RESETN(net2081),
    .SETN(net457));
 DFFASRHQNx1_ASAP7_75t_R _36586_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04339_),
    .QN(_00661_),
    .RESETN(net2082),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36587_ (.CLK(\clknet_leaf_6_core_clock_gate_i.clk_o ),
    .D(_04340_),
    .QN(_01315_),
    .RESETN(net2083),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36588_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_04341_),
    .QN(_01875_),
    .RESETN(net2084),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36589_ (.CLK(\clknet_leaf_3_core_clock_gate_i.clk_o ),
    .D(_04342_),
    .QN(_01874_),
    .RESETN(net2085),
    .SETN(net452));
 DFFASRHQNx1_ASAP7_75t_R _36590_ (.CLK(\clknet_leaf_1_core_clock_gate_i.clk_o ),
    .D(_04343_),
    .QN(_00285_),
    .RESETN(net2086),
    .SETN(net450));
 DFFASRHQNx1_ASAP7_75t_R _36591_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04344_),
    .QN(_01873_),
    .RESETN(net2087),
    .SETN(net449));
 DFFASRHQNx1_ASAP7_75t_R _36592_ (.CLK(\clknet_leaf_2_core_clock_gate_i.clk_o ),
    .D(_04345_),
    .QN(_01872_),
    .RESETN(net450),
    .SETN(net2088));
 DFFASRHQNx1_ASAP7_75t_R _36593_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3819),
    .QN(_01871_),
    .RESETN(net2089),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36594_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3873),
    .QN(_01870_),
    .RESETN(net2090),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36595_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3825),
    .QN(_01869_),
    .RESETN(net2091),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36596_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3879),
    .QN(_01868_),
    .RESETN(net2092),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36597_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3807),
    .QN(_01867_),
    .RESETN(net2093),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36598_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net2435),
    .QN(_01866_),
    .RESETN(net2094),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36599_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3831),
    .QN(_01865_),
    .RESETN(net2095),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36600_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3891),
    .QN(_01864_),
    .RESETN(net2096),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36601_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3861),
    .QN(_01863_),
    .RESETN(net2097),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36602_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3897),
    .QN(_01862_),
    .RESETN(net2098),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36603_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3849),
    .QN(_01861_),
    .RESETN(net2099),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36604_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3903),
    .QN(_01860_),
    .RESETN(net2100),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36605_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net2489),
    .QN(_01859_),
    .RESETN(net2101),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36606_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3855),
    .QN(_01858_),
    .RESETN(net2102),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36607_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3885),
    .QN(_01857_),
    .RESETN(net2103),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36608_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net2567),
    .QN(_01856_),
    .RESETN(net2104),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36609_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net2393),
    .QN(_01855_),
    .RESETN(net2105),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36610_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3837),
    .QN(_01854_),
    .RESETN(net2106),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36611_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3801),
    .QN(_01853_),
    .RESETN(net2107),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36612_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3843),
    .QN(_01852_),
    .RESETN(net2108),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36613_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3912),
    .QN(_01851_),
    .RESETN(net2109),
    .SETN(net460));
 DFFASRHQNx1_ASAP7_75t_R _36614_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net2477),
    .QN(_01850_),
    .RESETN(net2110),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36615_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3813),
    .QN(_01849_),
    .RESETN(net2111),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36616_ (.CLK(\clknet_leaf_5_core_clock_gate_i.clk_o ),
    .D(net3867),
    .QN(_01733_),
    .RESETN(net2112),
    .SETN(net441));
 DFFASRHQNx1_ASAP7_75t_R _36617_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(core_busy_d),
    .QN(_01734_),
    .RESETN(net2113),
    .SETN(net454));
 DLLx1_ASAP7_75t_R _36618_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(net3142),
    .Q(\core_clock_gate_i.en_latch ));
 DFFASRHQNx1_ASAP7_75t_R _36619_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(net2760),
    .QN(_00237_),
    .RESETN(net2114),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36620_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .QN(_01735_),
    .RESETN(net2115),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36621_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(net2462),
    .QN(_01736_),
    .RESETN(net2116),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36622_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(net2716),
    .QN(_00238_),
    .RESETN(net2117),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36623_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(net2978),
    .QN(_01737_),
    .RESETN(net2118),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36624_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(net2742),
    .QN(_01848_),
    .RESETN(net2119),
    .SETN(net454));
 DFFHQNx1_ASAP7_75t_R _36625_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04370_),
    .QN(_01847_));
 DFFHQNx1_ASAP7_75t_R _36626_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04371_),
    .QN(_01846_));
 DFFHQNx1_ASAP7_75t_R _36627_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04372_),
    .QN(_01845_));
 DFFHQNx1_ASAP7_75t_R _36628_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04373_),
    .QN(_01844_));
 DFFHQNx1_ASAP7_75t_R _36629_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04374_),
    .QN(_01843_));
 DFFHQNx1_ASAP7_75t_R _36630_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04375_),
    .QN(_01842_));
 DFFHQNx1_ASAP7_75t_R _36631_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04376_),
    .QN(_01841_));
 DFFHQNx1_ASAP7_75t_R _36632_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04377_),
    .QN(_01840_));
 DFFHQNx1_ASAP7_75t_R _36633_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04378_),
    .QN(_01839_));
 DFFHQNx1_ASAP7_75t_R _36634_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04379_),
    .QN(_01838_));
 DFFHQNx1_ASAP7_75t_R _36635_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04380_),
    .QN(_01837_));
 DFFHQNx1_ASAP7_75t_R _36636_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04381_),
    .QN(_01836_));
 DFFHQNx1_ASAP7_75t_R _36637_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04382_),
    .QN(_01835_));
 DFFHQNx1_ASAP7_75t_R _36638_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04383_),
    .QN(_01834_));
 DFFHQNx1_ASAP7_75t_R _36639_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04384_),
    .QN(_01833_));
 DFFHQNx1_ASAP7_75t_R _36640_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04385_),
    .QN(_01832_));
 DFFHQNx1_ASAP7_75t_R _36641_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04386_),
    .QN(_01831_));
 DFFHQNx1_ASAP7_75t_R _36642_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04387_),
    .QN(_01830_));
 DFFHQNx1_ASAP7_75t_R _36643_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04388_),
    .QN(_01829_));
 DFFHQNx1_ASAP7_75t_R _36644_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04389_),
    .QN(_01828_));
 DFFHQNx1_ASAP7_75t_R _36645_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04390_),
    .QN(_01827_));
 DFFHQNx1_ASAP7_75t_R _36646_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04391_),
    .QN(_01826_));
 DFFHQNx1_ASAP7_75t_R _36647_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04392_),
    .QN(_01825_));
 DFFHQNx1_ASAP7_75t_R _36648_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04393_),
    .QN(_01824_));
 DFFHQNx1_ASAP7_75t_R _36649_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04394_),
    .QN(_01823_));
 DFFHQNx1_ASAP7_75t_R _36650_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04395_),
    .QN(_01822_));
 DFFHQNx1_ASAP7_75t_R _36651_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04396_),
    .QN(_01821_));
 DFFHQNx1_ASAP7_75t_R _36652_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04397_),
    .QN(_01820_));
 DFFHQNx1_ASAP7_75t_R _36653_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04398_),
    .QN(_01819_));
 DFFHQNx1_ASAP7_75t_R _36654_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04399_),
    .QN(_01818_));
 DFFHQNx1_ASAP7_75t_R _36655_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04400_),
    .QN(_01817_));
 DFFHQNx1_ASAP7_75t_R _36656_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04401_),
    .QN(_01816_));
 DFFHQNx1_ASAP7_75t_R _36657_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04402_),
    .QN(_01738_));
 DFFASRHQNx1_ASAP7_75t_R _36658_ (.CLK(\clknet_leaf_23_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .QN(_00240_),
    .RESETN(net2120),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36659_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .QN(_00239_),
    .RESETN(net2121),
    .SETN(net454));
 DFFASRHQNx1_ASAP7_75t_R _36660_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .QN(_01815_),
    .RESETN(net2122),
    .SETN(net454));
 DFFHQNx1_ASAP7_75t_R _36661_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04403_),
    .QN(_01814_));
 DFFHQNx1_ASAP7_75t_R _36662_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04404_),
    .QN(_01813_));
 DFFHQNx1_ASAP7_75t_R _36663_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04405_),
    .QN(_01812_));
 DFFHQNx1_ASAP7_75t_R _36664_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04406_),
    .QN(_01811_));
 DFFHQNx1_ASAP7_75t_R _36665_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04407_),
    .QN(_01810_));
 DFFHQNx1_ASAP7_75t_R _36666_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04408_),
    .QN(_01809_));
 DFFHQNx1_ASAP7_75t_R _36667_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04409_),
    .QN(_01808_));
 DFFHQNx1_ASAP7_75t_R _36668_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04410_),
    .QN(_01807_));
 DFFHQNx1_ASAP7_75t_R _36669_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04411_),
    .QN(_01806_));
 DFFHQNx1_ASAP7_75t_R _36670_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04412_),
    .QN(_01805_));
 DFFHQNx1_ASAP7_75t_R _36671_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04413_),
    .QN(_01804_));
 DFFHQNx1_ASAP7_75t_R _36672_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04414_),
    .QN(_01803_));
 DFFHQNx1_ASAP7_75t_R _36673_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04415_),
    .QN(_01802_));
 DFFHQNx1_ASAP7_75t_R _36674_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04416_),
    .QN(_01801_));
 DFFHQNx1_ASAP7_75t_R _36675_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04417_),
    .QN(_01800_));
 DFFHQNx1_ASAP7_75t_R _36676_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04418_),
    .QN(_01799_));
 DFFHQNx1_ASAP7_75t_R _36677_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04419_),
    .QN(_01798_));
 DFFHQNx1_ASAP7_75t_R _36678_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04420_),
    .QN(_01797_));
 DFFHQNx1_ASAP7_75t_R _36679_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04421_),
    .QN(_01796_));
 DFFHQNx1_ASAP7_75t_R _36680_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04422_),
    .QN(_01795_));
 DFFHQNx1_ASAP7_75t_R _36681_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04423_),
    .QN(_01794_));
 DFFHQNx1_ASAP7_75t_R _36682_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04424_),
    .QN(_01793_));
 DFFHQNx1_ASAP7_75t_R _36683_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04425_),
    .QN(_01792_));
 DFFHQNx1_ASAP7_75t_R _36684_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04426_),
    .QN(_01791_));
 DFFHQNx1_ASAP7_75t_R _36685_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04427_),
    .QN(_01790_));
 DFFHQNx1_ASAP7_75t_R _36686_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(_04428_),
    .QN(_01789_));
 DFFHQNx1_ASAP7_75t_R _36687_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04429_),
    .QN(_01788_));
 DFFHQNx1_ASAP7_75t_R _36688_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04430_),
    .QN(_01787_));
 DFFHQNx1_ASAP7_75t_R _36689_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04431_),
    .QN(_01786_));
 DFFHQNx1_ASAP7_75t_R _36690_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04432_),
    .QN(_01785_));
 DFFHQNx1_ASAP7_75t_R _36691_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(_04433_),
    .QN(_01784_));
 DFFHQNx1_ASAP7_75t_R _36692_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04434_),
    .QN(_01783_));
 DFFHQNx1_ASAP7_75t_R _36693_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(_04435_),
    .QN(_01782_));
 DFFHQNx1_ASAP7_75t_R _36694_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(_04436_),
    .QN(_01781_));
 DFFHQNx1_ASAP7_75t_R _36695_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2576),
    .QN(_01780_));
 DFFHQNx1_ASAP7_75t_R _36696_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2554),
    .QN(_01779_));
 DFFHQNx1_ASAP7_75t_R _36697_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2426),
    .QN(_01778_));
 DFFHQNx1_ASAP7_75t_R _36698_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2544),
    .QN(_01777_));
 DFFHQNx1_ASAP7_75t_R _36699_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(net2802),
    .QN(_01776_));
 DFFHQNx1_ASAP7_75t_R _36700_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2453),
    .QN(_01775_));
 DFFHQNx1_ASAP7_75t_R _36701_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2468),
    .QN(_01774_));
 DFFHQNx1_ASAP7_75t_R _36702_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2471),
    .QN(_01773_));
 DFFHQNx1_ASAP7_75t_R _36703_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(net2561),
    .QN(_01772_));
 DFFHQNx1_ASAP7_75t_R _36704_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2450),
    .QN(_01771_));
 DFFHQNx1_ASAP7_75t_R _36705_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2517),
    .QN(_01770_));
 DFFHQNx1_ASAP7_75t_R _36706_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2432),
    .QN(_01769_));
 DFFHQNx1_ASAP7_75t_R _36707_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(net2408),
    .QN(_01768_));
 DFFHQNx1_ASAP7_75t_R _36708_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2501),
    .QN(_01767_));
 DFFHQNx1_ASAP7_75t_R _36709_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(net2429),
    .QN(_01766_));
 DFFHQNx1_ASAP7_75t_R _36710_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(net2402),
    .QN(_01765_));
 DFFHQNx1_ASAP7_75t_R _36711_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(net2610),
    .QN(_01764_));
 DFFHQNx1_ASAP7_75t_R _36712_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2474),
    .QN(_01763_));
 DFFHQNx1_ASAP7_75t_R _36713_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2465),
    .QN(_01762_));
 DFFHQNx1_ASAP7_75t_R _36714_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(net2587),
    .QN(_01761_));
 DFFHQNx1_ASAP7_75t_R _36715_ (.CLK(\clknet_leaf_31_core_clock_gate_i.clk_o ),
    .D(net2773),
    .QN(_01760_));
 DFFHQNx1_ASAP7_75t_R _36716_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2447),
    .QN(_01759_));
 DFFHQNx1_ASAP7_75t_R _36717_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2480),
    .QN(_01758_));
 DFFHQNx1_ASAP7_75t_R _36718_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2508),
    .QN(_01757_));
 DFFHQNx1_ASAP7_75t_R _36719_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2520),
    .QN(_01756_));
 DFFHQNx1_ASAP7_75t_R _36720_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2486),
    .QN(_01755_));
 DFFHQNx1_ASAP7_75t_R _36721_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2514),
    .QN(_01754_));
 DFFHQNx1_ASAP7_75t_R _36722_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2456),
    .QN(_01753_));
 DFFHQNx1_ASAP7_75t_R _36723_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(net2405),
    .QN(_01752_));
 DFFHQNx1_ASAP7_75t_R _36724_ (.CLK(\clknet_leaf_28_core_clock_gate_i.clk_o ),
    .D(net2492),
    .QN(_01751_));
 DFFHQNx1_ASAP7_75t_R _36725_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(net2411),
    .QN(_01750_));
 DFFHQNx1_ASAP7_75t_R _36726_ (.CLK(\clknet_leaf_30_core_clock_gate_i.clk_o ),
    .D(net2444),
    .QN(_01749_));
 DFFHQNx1_ASAP7_75t_R _36727_ (.CLK(\clknet_leaf_27_core_clock_gate_i.clk_o ),
    .D(net2530),
    .QN(_01748_));
 DFFASRHQNx1_ASAP7_75t_R _36728_ (.CLK(clknet_level_3_1_27107_clk_i),
    .D(net3952),
    .QN(_01747_),
    .RESETN(net2123),
    .SETN(net455));
 DFFHQNx1_ASAP7_75t_R _36729_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04471_),
    .QN(_01746_));
 DFFHQNx1_ASAP7_75t_R _36730_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04472_),
    .QN(_00163_));
 DFFHQNx1_ASAP7_75t_R _36731_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04473_),
    .QN(_00165_));
 DFFHQNx1_ASAP7_75t_R _36732_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04474_),
    .QN(_00168_));
 DFFHQNx1_ASAP7_75t_R _36733_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04475_),
    .QN(_00172_));
 DFFHQNx1_ASAP7_75t_R _36734_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04476_),
    .QN(_00175_));
 DFFHQNx1_ASAP7_75t_R _36735_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04477_),
    .QN(_00278_));
 DFFHQNx1_ASAP7_75t_R _36736_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04478_),
    .QN(_00323_));
 DFFHQNx1_ASAP7_75t_R _36737_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04479_),
    .QN(_00184_));
 DFFHQNx1_ASAP7_75t_R _36738_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04480_),
    .QN(_00187_));
 DFFHQNx1_ASAP7_75t_R _36739_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04481_),
    .QN(_00191_));
 DFFHQNx1_ASAP7_75t_R _36740_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04482_),
    .QN(_00194_));
 DFFHQNx1_ASAP7_75t_R _36741_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04483_),
    .QN(_00281_));
 DFFHQNx1_ASAP7_75t_R _36742_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04484_),
    .QN(_00282_));
 DFFHQNx1_ASAP7_75t_R _36743_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04485_),
    .QN(_00279_));
 DFFHQNx1_ASAP7_75t_R _36744_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04486_),
    .QN(_00290_));
 DFFHQNx1_ASAP7_75t_R _36745_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04487_),
    .QN(_00289_));
 DFFHQNx1_ASAP7_75t_R _36746_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04488_),
    .QN(_00288_));
 DFFHQNx1_ASAP7_75t_R _36747_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04489_),
    .QN(_00287_));
 DFFHQNx1_ASAP7_75t_R _36748_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04490_),
    .QN(_00286_));
 DFFHQNx1_ASAP7_75t_R _36749_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04491_),
    .QN(_00246_));
 DFFHQNx1_ASAP7_75t_R _36750_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04492_),
    .QN(_01745_));
 DFFHQNx1_ASAP7_75t_R _36751_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04493_),
    .QN(_01744_));
 DFFHQNx1_ASAP7_75t_R _36752_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04494_),
    .QN(_00245_));
 DFFHQNx1_ASAP7_75t_R _36753_ (.CLK(\clknet_leaf_0_core_clock_gate_i.clk_o ),
    .D(_04495_),
    .QN(_00244_));
 DFFHQNx1_ASAP7_75t_R _36754_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04496_),
    .QN(_01743_));
 DFFHQNx1_ASAP7_75t_R _36755_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04497_),
    .QN(_00283_));
 DFFHQNx1_ASAP7_75t_R _36756_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04498_),
    .QN(_01742_));
 DFFHQNx1_ASAP7_75t_R _36757_ (.CLK(\clknet_leaf_25_core_clock_gate_i.clk_o ),
    .D(_04499_),
    .QN(_01741_));
 DFFHQNx1_ASAP7_75t_R _36758_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04500_),
    .QN(_01740_));
 DFFHQNx1_ASAP7_75t_R _36759_ (.CLK(\clknet_leaf_26_core_clock_gate_i.clk_o ),
    .D(_04501_),
    .QN(_01739_));
 DFFHQNx1_ASAP7_75t_R _36760_ (.CLK(\clknet_leaf_29_core_clock_gate_i.clk_o ),
    .D(_04502_),
    .QN(_00280_));
 DFFASRHQNx1_ASAP7_75t_R _36761_ (.CLK(\clknet_leaf_24_core_clock_gate_i.clk_o ),
    .D(_04503_),
    .QN(_01311_),
    .RESETN(net2124),
    .SETN(net454));
 BUFx4_ASAP7_75t_R clkbuf_leaf_0_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_0_clk_i));
 TIEHIx1_ASAP7_75t_R _34880__467 (.H(net467));
 TAPCELL_ASAP7_75t_R PHY_30 ();
 BUFx2_ASAP7_75t_R _36765_ (.A(net462),
    .Y(alert_minor_o));
 BUFx2_ASAP7_75t_R _36766_ (.A(net463),
    .Y(data_addr_o[0]));
 BUFx2_ASAP7_75t_R _36767_ (.A(net464),
    .Y(data_addr_o[1]));
 TAPCELL_ASAP7_75t_R PHY_29 ();
 TAPCELL_ASAP7_75t_R PHY_28 ();
 TAPCELL_ASAP7_75t_R PHY_27 ();
 TAPCELL_ASAP7_75t_R PHY_26 ();
 TAPCELL_ASAP7_75t_R PHY_25 ();
 TAPCELL_ASAP7_75t_R PHY_24 ();
 TAPCELL_ASAP7_75t_R PHY_23 ();
 TAPCELL_ASAP7_75t_R PHY_22 ();
 TAPCELL_ASAP7_75t_R PHY_21 ();
 TAPCELL_ASAP7_75t_R PHY_20 ();
 TAPCELL_ASAP7_75t_R PHY_19 ();
 TAPCELL_ASAP7_75t_R PHY_18 ();
 TAPCELL_ASAP7_75t_R PHY_17 ();
 TAPCELL_ASAP7_75t_R PHY_16 ();
 TAPCELL_ASAP7_75t_R PHY_15 ();
 TAPCELL_ASAP7_75t_R PHY_14 ();
 TAPCELL_ASAP7_75t_R PHY_13 ();
 TAPCELL_ASAP7_75t_R PHY_12 ();
 TAPCELL_ASAP7_75t_R PHY_11 ();
 TAPCELL_ASAP7_75t_R PHY_10 ();
 TAPCELL_ASAP7_75t_R PHY_9 ();
 TAPCELL_ASAP7_75t_R PHY_8 ();
 TAPCELL_ASAP7_75t_R PHY_7 ();
 TAPCELL_ASAP7_75t_R PHY_6 ();
 TAPCELL_ASAP7_75t_R PHY_5 ();
 TAPCELL_ASAP7_75t_R PHY_4 ();
 TAPCELL_ASAP7_75t_R PHY_3 ();
 TAPCELL_ASAP7_75t_R PHY_2 ();
 TAPCELL_ASAP7_75t_R PHY_1 ();
 TAPCELL_ASAP7_75t_R PHY_0 ();
 BUFx2_ASAP7_75t_R _36798_ (.A(net465),
    .Y(instr_addr_o[0]));
 BUFx2_ASAP7_75t_R _36799_ (.A(net466),
    .Y(instr_addr_o[1]));
 TIEHIx1_ASAP7_75t_R _34952__539 (.H(net539));
 TIEHIx1_ASAP7_75t_R _34953__540 (.H(net540));
 TIEHIx1_ASAP7_75t_R _34954__541 (.H(net541));
 TIEHIx1_ASAP7_75t_R _34955__542 (.H(net542));
 TIEHIx1_ASAP7_75t_R _34956__543 (.H(net543));
 TIEHIx1_ASAP7_75t_R _34957__544 (.H(net544));
 TIEHIx1_ASAP7_75t_R _34958__545 (.H(net545));
 TIEHIx1_ASAP7_75t_R _34959__546 (.H(net546));
 TIEHIx1_ASAP7_75t_R _34960__547 (.H(net547));
 TIEHIx1_ASAP7_75t_R _34961__548 (.H(net548));
 TIEHIx1_ASAP7_75t_R _34962__549 (.H(net549));
 TIEHIx1_ASAP7_75t_R _34963__550 (.H(net550));
 TIEHIx1_ASAP7_75t_R _34964__551 (.H(net551));
 TIEHIx1_ASAP7_75t_R _34965__552 (.H(net552));
 TIEHIx1_ASAP7_75t_R _34966__553 (.H(net553));
 TIEHIx1_ASAP7_75t_R _34967__554 (.H(net554));
 TIEHIx1_ASAP7_75t_R _34968__555 (.H(net555));
 TIEHIx1_ASAP7_75t_R _34969__556 (.H(net556));
 TIEHIx1_ASAP7_75t_R _34970__557 (.H(net557));
 TIEHIx1_ASAP7_75t_R _34971__558 (.H(net558));
 TIEHIx1_ASAP7_75t_R _34972__559 (.H(net559));
 TIEHIx1_ASAP7_75t_R _34973__560 (.H(net560));
 TIEHIx1_ASAP7_75t_R _34974__561 (.H(net561));
 TIEHIx1_ASAP7_75t_R _34975__562 (.H(net562));
 TIEHIx1_ASAP7_75t_R _34976__563 (.H(net563));
 TIEHIx1_ASAP7_75t_R _34977__564 (.H(net564));
 TIEHIx1_ASAP7_75t_R _34978__565 (.H(net565));
 TIEHIx1_ASAP7_75t_R _34979__566 (.H(net566));
 TIEHIx1_ASAP7_75t_R _34980__567 (.H(net567));
 TIEHIx1_ASAP7_75t_R _34981__568 (.H(net568));
 TIEHIx1_ASAP7_75t_R _34982__569 (.H(net569));
 TIEHIx1_ASAP7_75t_R _34983__570 (.H(net570));
 TIEHIx1_ASAP7_75t_R _34984__571 (.H(net571));
 TIEHIx1_ASAP7_75t_R _34985__572 (.H(net572));
 TIEHIx1_ASAP7_75t_R _34986__573 (.H(net573));
 TIEHIx1_ASAP7_75t_R _34987__574 (.H(net574));
 TIEHIx1_ASAP7_75t_R _34988__575 (.H(net575));
 TIEHIx1_ASAP7_75t_R _34989__576 (.H(net576));
 TIEHIx1_ASAP7_75t_R _34990__577 (.H(net577));
 TIEHIx1_ASAP7_75t_R _34991__578 (.H(net578));
 TIEHIx1_ASAP7_75t_R _34992__579 (.H(net579));
 TIEHIx1_ASAP7_75t_R _34993__580 (.H(net580));
 TIEHIx1_ASAP7_75t_R _34994__581 (.H(net581));
 TIEHIx1_ASAP7_75t_R _34995__582 (.H(net582));
 TIEHIx1_ASAP7_75t_R _34996__583 (.H(net583));
 TIEHIx1_ASAP7_75t_R _34997__584 (.H(net584));
 TIEHIx1_ASAP7_75t_R _34998__585 (.H(net585));
 TIEHIx1_ASAP7_75t_R _34999__586 (.H(net586));
 TIEHIx1_ASAP7_75t_R _35000__587 (.H(net587));
 TIEHIx1_ASAP7_75t_R _35001__588 (.H(net588));
 TIEHIx1_ASAP7_75t_R _35002__589 (.H(net589));
 TIEHIx1_ASAP7_75t_R _35003__590 (.H(net590));
 TIEHIx1_ASAP7_75t_R _35004__591 (.H(net591));
 TIEHIx1_ASAP7_75t_R _35005__592 (.H(net592));
 TIEHIx1_ASAP7_75t_R _35006__593 (.H(net593));
 TIEHIx1_ASAP7_75t_R _35007__594 (.H(net594));
 TIEHIx1_ASAP7_75t_R _35008__595 (.H(net595));
 TIEHIx1_ASAP7_75t_R _35009__596 (.H(net596));
 TIEHIx1_ASAP7_75t_R _35010__597 (.H(net597));
 TIEHIx1_ASAP7_75t_R _35011__598 (.H(net598));
 TIEHIx1_ASAP7_75t_R _35012__599 (.H(net599));
 TIEHIx1_ASAP7_75t_R _35013__600 (.H(net600));
 TIEHIx1_ASAP7_75t_R _35014__601 (.H(net601));
 TIEHIx1_ASAP7_75t_R _35015__602 (.H(net602));
 TIEHIx1_ASAP7_75t_R _35016__603 (.H(net603));
 TIEHIx1_ASAP7_75t_R _35017__604 (.H(net604));
 TIEHIx1_ASAP7_75t_R _35018__605 (.H(net605));
 TIEHIx1_ASAP7_75t_R _35019__606 (.H(net606));
 TIEHIx1_ASAP7_75t_R _35020__607 (.H(net607));
 TIEHIx1_ASAP7_75t_R _35021__608 (.H(net608));
 TIEHIx1_ASAP7_75t_R _35022__609 (.H(net609));
 TIEHIx1_ASAP7_75t_R _35023__610 (.H(net610));
 TIEHIx1_ASAP7_75t_R _35024__611 (.H(net611));
 TIEHIx1_ASAP7_75t_R _35025__612 (.H(net612));
 TIEHIx1_ASAP7_75t_R _35026__613 (.H(net613));
 TIEHIx1_ASAP7_75t_R _35027__614 (.H(net614));
 TIEHIx1_ASAP7_75t_R _35028__615 (.H(net615));
 TIEHIx1_ASAP7_75t_R _35029__616 (.H(net616));
 TIEHIx1_ASAP7_75t_R _35030__617 (.H(net617));
 TIEHIx1_ASAP7_75t_R _35031__618 (.H(net618));
 TIEHIx1_ASAP7_75t_R _35032__619 (.H(net619));
 TIEHIx1_ASAP7_75t_R _35033__620 (.H(net620));
 TIEHIx1_ASAP7_75t_R _35034__621 (.H(net621));
 TIEHIx1_ASAP7_75t_R _35035__622 (.H(net622));
 TIEHIx1_ASAP7_75t_R _35036__623 (.H(net623));
 TIEHIx1_ASAP7_75t_R _35037__624 (.H(net624));
 TIEHIx1_ASAP7_75t_R _35038__625 (.H(net625));
 TIEHIx1_ASAP7_75t_R _35039__626 (.H(net626));
 TIEHIx1_ASAP7_75t_R _35040__627 (.H(net627));
 TIEHIx1_ASAP7_75t_R _35041__628 (.H(net628));
 TIEHIx1_ASAP7_75t_R _35042__629 (.H(net629));
 TIEHIx1_ASAP7_75t_R _35043__630 (.H(net630));
 TIEHIx1_ASAP7_75t_R _35044__631 (.H(net631));
 TIEHIx1_ASAP7_75t_R _35045__632 (.H(net632));
 TIEHIx1_ASAP7_75t_R _35046__633 (.H(net633));
 TIEHIx1_ASAP7_75t_R _35047__634 (.H(net634));
 TIEHIx1_ASAP7_75t_R _35048__635 (.H(net635));
 TIEHIx1_ASAP7_75t_R _35049__636 (.H(net636));
 TIEHIx1_ASAP7_75t_R _35050__637 (.H(net637));
 TIEHIx1_ASAP7_75t_R _35051__638 (.H(net638));
 TIEHIx1_ASAP7_75t_R _35052__639 (.H(net639));
 TIEHIx1_ASAP7_75t_R _35053__640 (.H(net640));
 TIEHIx1_ASAP7_75t_R _35054__641 (.H(net641));
 TIEHIx1_ASAP7_75t_R _35055__642 (.H(net642));
 TIEHIx1_ASAP7_75t_R _35056__643 (.H(net643));
 TIEHIx1_ASAP7_75t_R _35057__644 (.H(net644));
 TIEHIx1_ASAP7_75t_R _35058__645 (.H(net645));
 TIEHIx1_ASAP7_75t_R _35059__646 (.H(net646));
 TIEHIx1_ASAP7_75t_R _35060__647 (.H(net647));
 TIEHIx1_ASAP7_75t_R _35061__648 (.H(net648));
 TIEHIx1_ASAP7_75t_R _35062__649 (.H(net649));
 TIEHIx1_ASAP7_75t_R _35063__650 (.H(net650));
 TIEHIx1_ASAP7_75t_R _35064__651 (.H(net651));
 TIEHIx1_ASAP7_75t_R _35065__652 (.H(net652));
 TIEHIx1_ASAP7_75t_R _35066__653 (.H(net653));
 TIEHIx1_ASAP7_75t_R _35067__654 (.H(net654));
 TIEHIx1_ASAP7_75t_R _35068__655 (.H(net655));
 TIEHIx1_ASAP7_75t_R _35069__656 (.H(net656));
 TIEHIx1_ASAP7_75t_R _35070__657 (.H(net657));
 TIEHIx1_ASAP7_75t_R _35071__658 (.H(net658));
 TIEHIx1_ASAP7_75t_R _35072__659 (.H(net659));
 TIEHIx1_ASAP7_75t_R _35073__660 (.H(net660));
 TIEHIx1_ASAP7_75t_R _35074__661 (.H(net661));
 TIEHIx1_ASAP7_75t_R _35106__662 (.H(net662));
 TIEHIx1_ASAP7_75t_R _35107__663 (.H(net663));
 TIEHIx1_ASAP7_75t_R _35108__664 (.H(net664));
 TIEHIx1_ASAP7_75t_R _35109__665 (.H(net665));
 TIEHIx1_ASAP7_75t_R _35110__666 (.H(net666));
 TIEHIx1_ASAP7_75t_R _35111__667 (.H(net667));
 TIEHIx1_ASAP7_75t_R _35112__668 (.H(net668));
 TIEHIx1_ASAP7_75t_R _35113__669 (.H(net669));
 TIEHIx1_ASAP7_75t_R _35114__670 (.H(net670));
 TIEHIx1_ASAP7_75t_R _35115__671 (.H(net671));
 TIEHIx1_ASAP7_75t_R _35116__672 (.H(net672));
 TIEHIx1_ASAP7_75t_R _35117__673 (.H(net673));
 TIEHIx1_ASAP7_75t_R _35118__674 (.H(net674));
 TIEHIx1_ASAP7_75t_R _35119__675 (.H(net675));
 TIEHIx1_ASAP7_75t_R _35120__676 (.H(net676));
 TIEHIx1_ASAP7_75t_R _35121__677 (.H(net677));
 TIEHIx1_ASAP7_75t_R _35122__678 (.H(net678));
 TIEHIx1_ASAP7_75t_R _35123__679 (.H(net679));
 TIEHIx1_ASAP7_75t_R _35124__680 (.H(net680));
 TIEHIx1_ASAP7_75t_R _35125__681 (.H(net681));
 TIEHIx1_ASAP7_75t_R _35126__682 (.H(net682));
 TIEHIx1_ASAP7_75t_R _35127__683 (.H(net683));
 TIEHIx1_ASAP7_75t_R _35128__684 (.H(net684));
 TIEHIx1_ASAP7_75t_R _35129__685 (.H(net685));
 TIEHIx1_ASAP7_75t_R _35130__686 (.H(net686));
 TIEHIx1_ASAP7_75t_R _35131__687 (.H(net687));
 TIEHIx1_ASAP7_75t_R _35132__688 (.H(net688));
 TIEHIx1_ASAP7_75t_R _35133__689 (.H(net689));
 TIEHIx1_ASAP7_75t_R _35134__690 (.H(net690));
 TIEHIx1_ASAP7_75t_R _35135__691 (.H(net691));
 TIEHIx1_ASAP7_75t_R _35136__692 (.H(net692));
 TIEHIx1_ASAP7_75t_R _35137__693 (.H(net693));
 TIEHIx1_ASAP7_75t_R _35138__694 (.H(net694));
 TIEHIx1_ASAP7_75t_R _35169__695 (.H(net695));
 TIEHIx1_ASAP7_75t_R _35170__696 (.H(net696));
 TIEHIx1_ASAP7_75t_R _35171__697 (.H(net697));
 TIEHIx1_ASAP7_75t_R _35172__698 (.H(net698));
 TIEHIx1_ASAP7_75t_R _35173__699 (.H(net699));
 TIEHIx1_ASAP7_75t_R _35174__700 (.H(net700));
 TIEHIx1_ASAP7_75t_R _35175__701 (.H(net701));
 TIEHIx1_ASAP7_75t_R _35176__702 (.H(net702));
 TIEHIx1_ASAP7_75t_R _35177__703 (.H(net703));
 TIEHIx1_ASAP7_75t_R _35178__704 (.H(net704));
 TIEHIx1_ASAP7_75t_R _35179__705 (.H(net705));
 TIEHIx1_ASAP7_75t_R _35180__706 (.H(net706));
 TIEHIx1_ASAP7_75t_R _35181__707 (.H(net707));
 TIEHIx1_ASAP7_75t_R _35182__708 (.H(net708));
 TIEHIx1_ASAP7_75t_R _35183__709 (.H(net709));
 TIEHIx1_ASAP7_75t_R _35184__710 (.H(net710));
 TIEHIx1_ASAP7_75t_R _35185__711 (.H(net711));
 TIEHIx1_ASAP7_75t_R _35186__712 (.H(net712));
 TIEHIx1_ASAP7_75t_R _35187__713 (.H(net713));
 TIEHIx1_ASAP7_75t_R _35188__714 (.H(net714));
 TIEHIx1_ASAP7_75t_R _35189__715 (.H(net715));
 TIEHIx1_ASAP7_75t_R _35190__716 (.H(net716));
 TIEHIx1_ASAP7_75t_R _35191__717 (.H(net717));
 TIEHIx1_ASAP7_75t_R _35192__718 (.H(net718));
 TIEHIx1_ASAP7_75t_R _35193__719 (.H(net719));
 TIEHIx1_ASAP7_75t_R _35194__720 (.H(net720));
 TIEHIx1_ASAP7_75t_R _35195__721 (.H(net721));
 TIEHIx1_ASAP7_75t_R _35196__722 (.H(net722));
 TIEHIx1_ASAP7_75t_R _35197__723 (.H(net723));
 TIEHIx1_ASAP7_75t_R _35198__724 (.H(net724));
 TIEHIx1_ASAP7_75t_R _35199__725 (.H(net725));
 TIEHIx1_ASAP7_75t_R _35200__726 (.H(net726));
 TIEHIx1_ASAP7_75t_R _35201__727 (.H(net727));
 TIEHIx1_ASAP7_75t_R _35202__728 (.H(net728));
 TIEHIx1_ASAP7_75t_R _35203__729 (.H(net729));
 TIEHIx1_ASAP7_75t_R _35204__730 (.H(net730));
 TIEHIx1_ASAP7_75t_R _35205__731 (.H(net731));
 TIEHIx1_ASAP7_75t_R _35206__732 (.H(net732));
 TIEHIx1_ASAP7_75t_R _35207__733 (.H(net733));
 TIEHIx1_ASAP7_75t_R _35208__734 (.H(net734));
 TIEHIx1_ASAP7_75t_R _35209__735 (.H(net735));
 TIEHIx1_ASAP7_75t_R _35210__736 (.H(net736));
 TIEHIx1_ASAP7_75t_R _35211__737 (.H(net737));
 TIEHIx1_ASAP7_75t_R _35212__738 (.H(net738));
 TIEHIx1_ASAP7_75t_R _35213__739 (.H(net739));
 TIEHIx1_ASAP7_75t_R _35214__740 (.H(net740));
 TIEHIx1_ASAP7_75t_R _35215__741 (.H(net741));
 TIEHIx1_ASAP7_75t_R _35216__742 (.H(net742));
 TIEHIx1_ASAP7_75t_R _35217__743 (.H(net743));
 TIEHIx1_ASAP7_75t_R _35218__744 (.H(net744));
 TIEHIx1_ASAP7_75t_R _35219__745 (.H(net745));
 TIEHIx1_ASAP7_75t_R _35220__746 (.H(net746));
 TIEHIx1_ASAP7_75t_R _35221__747 (.H(net747));
 TIEHIx1_ASAP7_75t_R _35222__748 (.H(net748));
 TIEHIx1_ASAP7_75t_R _35223__749 (.H(net749));
 TIEHIx1_ASAP7_75t_R _35224__750 (.H(net750));
 TIEHIx1_ASAP7_75t_R _35225__751 (.H(net751));
 TIEHIx1_ASAP7_75t_R _35226__752 (.H(net752));
 TIEHIx1_ASAP7_75t_R _35227__753 (.H(net753));
 TIEHIx1_ASAP7_75t_R _35228__754 (.H(net754));
 TIEHIx1_ASAP7_75t_R _35229__755 (.H(net755));
 TIEHIx1_ASAP7_75t_R _35230__756 (.H(net756));
 TIEHIx1_ASAP7_75t_R _35231__757 (.H(net757));
 TIEHIx1_ASAP7_75t_R _35232__758 (.H(net758));
 TIEHIx1_ASAP7_75t_R _35233__759 (.H(net759));
 TIEHIx1_ASAP7_75t_R _35234__760 (.H(net760));
 TIEHIx1_ASAP7_75t_R _35235__761 (.H(net761));
 TIEHIx1_ASAP7_75t_R _35236__762 (.H(net762));
 TIEHIx1_ASAP7_75t_R _35237__763 (.H(net763));
 TIEHIx1_ASAP7_75t_R _35238__764 (.H(net764));
 TIEHIx1_ASAP7_75t_R _35239__765 (.H(net765));
 TIEHIx1_ASAP7_75t_R _35240__766 (.H(net766));
 TIEHIx1_ASAP7_75t_R _35241__767 (.H(net767));
 TIEHIx1_ASAP7_75t_R _35242__768 (.H(net768));
 TIEHIx1_ASAP7_75t_R _35243__769 (.H(net769));
 TIEHIx1_ASAP7_75t_R _35244__770 (.H(net770));
 TIEHIx1_ASAP7_75t_R _35245__771 (.H(net771));
 TIEHIx1_ASAP7_75t_R _35246__772 (.H(net772));
 TIEHIx1_ASAP7_75t_R _35247__773 (.H(net773));
 TIEHIx1_ASAP7_75t_R _35248__774 (.H(net774));
 TIEHIx1_ASAP7_75t_R _35249__775 (.H(net775));
 TIEHIx1_ASAP7_75t_R _35250__776 (.H(net776));
 TIEHIx1_ASAP7_75t_R _35251__777 (.H(net777));
 TIEHIx1_ASAP7_75t_R _35252__778 (.H(net778));
 TIEHIx1_ASAP7_75t_R _35253__779 (.H(net779));
 TIEHIx1_ASAP7_75t_R _35254__780 (.H(net780));
 TIEHIx1_ASAP7_75t_R _35255__781 (.H(net781));
 TIEHIx1_ASAP7_75t_R _35256__782 (.H(net782));
 TIEHIx1_ASAP7_75t_R _35257__783 (.H(net783));
 TIEHIx1_ASAP7_75t_R _35258__784 (.H(net784));
 TIEHIx1_ASAP7_75t_R _35259__785 (.H(net785));
 TIEHIx1_ASAP7_75t_R _35260__786 (.H(net786));
 TIEHIx1_ASAP7_75t_R _35261__787 (.H(net787));
 TIEHIx1_ASAP7_75t_R _35262__788 (.H(net788));
 TIEHIx1_ASAP7_75t_R _35263__789 (.H(net789));
 TIEHIx1_ASAP7_75t_R _35264__790 (.H(net790));
 TIEHIx1_ASAP7_75t_R _35265__791 (.H(net791));
 TIEHIx1_ASAP7_75t_R _35266__792 (.H(net792));
 TIEHIx1_ASAP7_75t_R _35267__793 (.H(net793));
 TIEHIx1_ASAP7_75t_R _35268__794 (.H(net794));
 TIEHIx1_ASAP7_75t_R _35269__795 (.H(net795));
 TIEHIx1_ASAP7_75t_R _35270__796 (.H(net796));
 TIEHIx1_ASAP7_75t_R _35271__797 (.H(net797));
 TIEHIx1_ASAP7_75t_R _35272__798 (.H(net798));
 TIEHIx1_ASAP7_75t_R _35273__799 (.H(net799));
 TIEHIx1_ASAP7_75t_R _35274__800 (.H(net800));
 TIEHIx1_ASAP7_75t_R _35275__801 (.H(net801));
 TIEHIx1_ASAP7_75t_R _35276__802 (.H(net802));
 TIEHIx1_ASAP7_75t_R _35277__803 (.H(net803));
 TIEHIx1_ASAP7_75t_R _35278__804 (.H(net804));
 TIEHIx1_ASAP7_75t_R _35279__805 (.H(net805));
 TIEHIx1_ASAP7_75t_R _35280__806 (.H(net806));
 TIEHIx1_ASAP7_75t_R _35281__807 (.H(net807));
 TIEHIx1_ASAP7_75t_R _35282__808 (.H(net808));
 TIEHIx1_ASAP7_75t_R _35283__809 (.H(net809));
 TIEHIx1_ASAP7_75t_R _35284__810 (.H(net810));
 TIEHIx1_ASAP7_75t_R _35285__811 (.H(net811));
 TIEHIx1_ASAP7_75t_R _35286__812 (.H(net812));
 TIEHIx1_ASAP7_75t_R _35287__813 (.H(net813));
 TIEHIx1_ASAP7_75t_R _35288__814 (.H(net814));
 TIEHIx1_ASAP7_75t_R _35289__815 (.H(net815));
 TIEHIx1_ASAP7_75t_R _35290__816 (.H(net816));
 TIEHIx1_ASAP7_75t_R _35291__817 (.H(net817));
 TIEHIx1_ASAP7_75t_R _35292__818 (.H(net818));
 TIEHIx1_ASAP7_75t_R _35293__819 (.H(net819));
 TIEHIx1_ASAP7_75t_R _35294__820 (.H(net820));
 TIEHIx1_ASAP7_75t_R _35295__821 (.H(net821));
 TIEHIx1_ASAP7_75t_R _35296__822 (.H(net822));
 TIEHIx1_ASAP7_75t_R _35297__823 (.H(net823));
 TIEHIx1_ASAP7_75t_R _35298__824 (.H(net824));
 TIEHIx1_ASAP7_75t_R _35299__825 (.H(net825));
 TIEHIx1_ASAP7_75t_R _35300__826 (.H(net826));
 TIEHIx1_ASAP7_75t_R _35301__827 (.H(net827));
 TIEHIx1_ASAP7_75t_R _35302__828 (.H(net828));
 TIEHIx1_ASAP7_75t_R _35303__829 (.H(net829));
 TIEHIx1_ASAP7_75t_R _35304__830 (.H(net830));
 TIEHIx1_ASAP7_75t_R _35305__831 (.H(net831));
 TIEHIx1_ASAP7_75t_R _35306__832 (.H(net832));
 TIEHIx1_ASAP7_75t_R _35307__833 (.H(net833));
 TIEHIx1_ASAP7_75t_R _35308__834 (.H(net834));
 TIEHIx1_ASAP7_75t_R _35309__835 (.H(net835));
 TIEHIx1_ASAP7_75t_R _35310__836 (.H(net836));
 TIEHIx1_ASAP7_75t_R _35311__837 (.H(net837));
 TIEHIx1_ASAP7_75t_R _35312__838 (.H(net838));
 TIEHIx1_ASAP7_75t_R _35313__839 (.H(net839));
 TIEHIx1_ASAP7_75t_R _35314__840 (.H(net840));
 TIEHIx1_ASAP7_75t_R _35315__841 (.H(net841));
 TIEHIx1_ASAP7_75t_R _35316__842 (.H(net842));
 TIEHIx1_ASAP7_75t_R _35317__843 (.H(net843));
 TIEHIx1_ASAP7_75t_R _35318__844 (.H(net844));
 TIEHIx1_ASAP7_75t_R _35319__845 (.H(net845));
 TIEHIx1_ASAP7_75t_R _35320__846 (.H(net846));
 TIEHIx1_ASAP7_75t_R _35321__847 (.H(net847));
 TIEHIx1_ASAP7_75t_R _35322__848 (.H(net848));
 TIEHIx1_ASAP7_75t_R _35323__849 (.H(net849));
 TIEHIx1_ASAP7_75t_R _35324__850 (.H(net850));
 TIEHIx1_ASAP7_75t_R _35325__851 (.H(net851));
 TIEHIx1_ASAP7_75t_R _35326__852 (.H(net852));
 TIEHIx1_ASAP7_75t_R _35327__853 (.H(net853));
 TIEHIx1_ASAP7_75t_R _35328__854 (.H(net854));
 TIEHIx1_ASAP7_75t_R _35329__855 (.H(net855));
 TIEHIx1_ASAP7_75t_R _35330__856 (.H(net856));
 TIEHIx1_ASAP7_75t_R _35331__857 (.H(net857));
 TIEHIx1_ASAP7_75t_R _35332__858 (.H(net858));
 TIEHIx1_ASAP7_75t_R _35333__859 (.H(net859));
 TIEHIx1_ASAP7_75t_R _35334__860 (.H(net860));
 TIEHIx1_ASAP7_75t_R _35335__861 (.H(net861));
 TIEHIx1_ASAP7_75t_R _35336__862 (.H(net862));
 TIEHIx1_ASAP7_75t_R _35337__863 (.H(net863));
 TIEHIx1_ASAP7_75t_R _35338__864 (.H(net864));
 TIEHIx1_ASAP7_75t_R _35339__865 (.H(net865));
 TIEHIx1_ASAP7_75t_R _35340__866 (.H(net866));
 TIEHIx1_ASAP7_75t_R _35341__867 (.H(net867));
 TIEHIx1_ASAP7_75t_R _35342__868 (.H(net868));
 TIEHIx1_ASAP7_75t_R _35343__869 (.H(net869));
 TIEHIx1_ASAP7_75t_R _35344__870 (.H(net870));
 TIEHIx1_ASAP7_75t_R _35345__871 (.H(net871));
 TIEHIx1_ASAP7_75t_R _35346__872 (.H(net872));
 TIEHIx1_ASAP7_75t_R _35347__873 (.H(net873));
 TIEHIx1_ASAP7_75t_R _35348__874 (.H(net874));
 TIEHIx1_ASAP7_75t_R _35349__875 (.H(net875));
 TIEHIx1_ASAP7_75t_R _35350__876 (.H(net876));
 TIEHIx1_ASAP7_75t_R _35351__877 (.H(net877));
 TIEHIx1_ASAP7_75t_R _35352__878 (.H(net878));
 TIEHIx1_ASAP7_75t_R _35353__879 (.H(net879));
 TIEHIx1_ASAP7_75t_R _35354__880 (.H(net880));
 TIEHIx1_ASAP7_75t_R _35355__881 (.H(net881));
 TIEHIx1_ASAP7_75t_R _35356__882 (.H(net882));
 TIEHIx1_ASAP7_75t_R _35357__883 (.H(net883));
 TIEHIx1_ASAP7_75t_R _35358__884 (.H(net884));
 TIEHIx1_ASAP7_75t_R _35359__885 (.H(net885));
 TIEHIx1_ASAP7_75t_R _35360__886 (.H(net886));
 TIEHIx1_ASAP7_75t_R _35361__887 (.H(net887));
 TIEHIx1_ASAP7_75t_R _35362__888 (.H(net888));
 TIEHIx1_ASAP7_75t_R _35363__889 (.H(net889));
 TIEHIx1_ASAP7_75t_R _35364__890 (.H(net890));
 TIEHIx1_ASAP7_75t_R _35365__891 (.H(net891));
 TIEHIx1_ASAP7_75t_R _35366__892 (.H(net892));
 TIEHIx1_ASAP7_75t_R _35367__893 (.H(net893));
 TIEHIx1_ASAP7_75t_R _35368__894 (.H(net894));
 TIEHIx1_ASAP7_75t_R _35369__895 (.H(net895));
 TIEHIx1_ASAP7_75t_R _35370__896 (.H(net896));
 TIEHIx1_ASAP7_75t_R _35371__897 (.H(net897));
 TIEHIx1_ASAP7_75t_R _35372__898 (.H(net898));
 TIEHIx1_ASAP7_75t_R _35373__899 (.H(net899));
 TIEHIx1_ASAP7_75t_R _35374__900 (.H(net900));
 TIEHIx1_ASAP7_75t_R _35375__901 (.H(net901));
 TIEHIx1_ASAP7_75t_R _35376__902 (.H(net902));
 TIEHIx1_ASAP7_75t_R _35377__903 (.H(net903));
 TIEHIx1_ASAP7_75t_R _35378__904 (.H(net904));
 TIEHIx1_ASAP7_75t_R _35379__905 (.H(net905));
 TIEHIx1_ASAP7_75t_R _35380__906 (.H(net906));
 TIEHIx1_ASAP7_75t_R _35381__907 (.H(net907));
 TIEHIx1_ASAP7_75t_R _35382__908 (.H(net908));
 TIEHIx1_ASAP7_75t_R _35383__909 (.H(net909));
 TIEHIx1_ASAP7_75t_R _35384__910 (.H(net910));
 TIEHIx1_ASAP7_75t_R _35385__911 (.H(net911));
 TIEHIx1_ASAP7_75t_R _35386__912 (.H(net912));
 TIEHIx1_ASAP7_75t_R _35387__913 (.H(net913));
 TIEHIx1_ASAP7_75t_R _35388__914 (.H(net914));
 TIEHIx1_ASAP7_75t_R _35389__915 (.H(net915));
 TIEHIx1_ASAP7_75t_R _35390__916 (.H(net916));
 TIEHIx1_ASAP7_75t_R _35391__917 (.H(net917));
 TIEHIx1_ASAP7_75t_R _35392__918 (.H(net918));
 TIEHIx1_ASAP7_75t_R _35393__919 (.H(net919));
 TIEHIx1_ASAP7_75t_R _35394__920 (.H(net920));
 TIEHIx1_ASAP7_75t_R _35395__921 (.H(net921));
 TIEHIx1_ASAP7_75t_R _35396__922 (.H(net922));
 TIEHIx1_ASAP7_75t_R _35397__923 (.H(net923));
 TIEHIx1_ASAP7_75t_R _35398__924 (.H(net924));
 TIEHIx1_ASAP7_75t_R _35399__925 (.H(net925));
 TIEHIx1_ASAP7_75t_R _35400__926 (.H(net926));
 TIEHIx1_ASAP7_75t_R _35401__927 (.H(net927));
 TIEHIx1_ASAP7_75t_R _35402__928 (.H(net928));
 TIEHIx1_ASAP7_75t_R _35403__929 (.H(net929));
 TIEHIx1_ASAP7_75t_R _35404__930 (.H(net930));
 TIEHIx1_ASAP7_75t_R _35405__931 (.H(net931));
 TIEHIx1_ASAP7_75t_R _35406__932 (.H(net932));
 TIEHIx1_ASAP7_75t_R _35407__933 (.H(net933));
 TIEHIx1_ASAP7_75t_R _35408__934 (.H(net934));
 TIEHIx1_ASAP7_75t_R _35409__935 (.H(net935));
 TIEHIx1_ASAP7_75t_R _35410__936 (.H(net936));
 TIEHIx1_ASAP7_75t_R _35411__937 (.H(net937));
 TIEHIx1_ASAP7_75t_R _35412__938 (.H(net938));
 TIEHIx1_ASAP7_75t_R _35413__939 (.H(net939));
 TIEHIx1_ASAP7_75t_R _35414__940 (.H(net940));
 TIEHIx1_ASAP7_75t_R _35415__941 (.H(net941));
 TIEHIx1_ASAP7_75t_R _35416__942 (.H(net942));
 TIEHIx1_ASAP7_75t_R _35417__943 (.H(net943));
 TIEHIx1_ASAP7_75t_R _35418__944 (.H(net944));
 TIEHIx1_ASAP7_75t_R _35419__945 (.H(net945));
 TIEHIx1_ASAP7_75t_R _35420__946 (.H(net946));
 TIEHIx1_ASAP7_75t_R _35421__947 (.H(net947));
 TIEHIx1_ASAP7_75t_R _35422__948 (.H(net948));
 TIEHIx1_ASAP7_75t_R _35423__949 (.H(net949));
 TIEHIx1_ASAP7_75t_R _35424__950 (.H(net950));
 TIEHIx1_ASAP7_75t_R _35425__951 (.H(net951));
 TIEHIx1_ASAP7_75t_R _35426__952 (.H(net952));
 TIEHIx1_ASAP7_75t_R _35427__953 (.H(net953));
 TIEHIx1_ASAP7_75t_R _35428__954 (.H(net954));
 TIEHIx1_ASAP7_75t_R _35429__955 (.H(net955));
 TIEHIx1_ASAP7_75t_R _35430__956 (.H(net956));
 TIEHIx1_ASAP7_75t_R _35431__957 (.H(net957));
 TIEHIx1_ASAP7_75t_R _35432__958 (.H(net958));
 TIEHIx1_ASAP7_75t_R _35433__959 (.H(net959));
 TIEHIx1_ASAP7_75t_R _35434__960 (.H(net960));
 TIEHIx1_ASAP7_75t_R _35435__961 (.H(net961));
 TIEHIx1_ASAP7_75t_R _35436__962 (.H(net962));
 TIEHIx1_ASAP7_75t_R _35437__963 (.H(net963));
 TIEHIx1_ASAP7_75t_R _35438__964 (.H(net964));
 TIEHIx1_ASAP7_75t_R _35439__965 (.H(net965));
 TIEHIx1_ASAP7_75t_R _35440__966 (.H(net966));
 TIEHIx1_ASAP7_75t_R _35441__967 (.H(net967));
 TIEHIx1_ASAP7_75t_R _35442__968 (.H(net968));
 TIEHIx1_ASAP7_75t_R _35443__969 (.H(net969));
 TIEHIx1_ASAP7_75t_R _35444__970 (.H(net970));
 TIEHIx1_ASAP7_75t_R _35445__971 (.H(net971));
 TIEHIx1_ASAP7_75t_R _35446__972 (.H(net972));
 TIEHIx1_ASAP7_75t_R _35447__973 (.H(net973));
 TIEHIx1_ASAP7_75t_R _35448__974 (.H(net974));
 TIEHIx1_ASAP7_75t_R _35449__975 (.H(net975));
 TIEHIx1_ASAP7_75t_R _35450__976 (.H(net976));
 TIEHIx1_ASAP7_75t_R _35451__977 (.H(net977));
 TIEHIx1_ASAP7_75t_R _35452__978 (.H(net978));
 TIEHIx1_ASAP7_75t_R _35453__979 (.H(net979));
 TIEHIx1_ASAP7_75t_R _35454__980 (.H(net980));
 TIEHIx1_ASAP7_75t_R _35455__981 (.H(net981));
 TIEHIx1_ASAP7_75t_R _35456__982 (.H(net982));
 TIEHIx1_ASAP7_75t_R _35457__983 (.H(net983));
 TIEHIx1_ASAP7_75t_R _35458__984 (.H(net984));
 TIEHIx1_ASAP7_75t_R _35459__985 (.H(net985));
 TIEHIx1_ASAP7_75t_R _35460__986 (.H(net986));
 TIEHIx1_ASAP7_75t_R _35461__987 (.H(net987));
 TIEHIx1_ASAP7_75t_R _35462__988 (.H(net988));
 TIEHIx1_ASAP7_75t_R _35463__989 (.H(net989));
 TIEHIx1_ASAP7_75t_R _35464__990 (.H(net990));
 TIEHIx1_ASAP7_75t_R _35465__991 (.H(net991));
 TIEHIx1_ASAP7_75t_R _35466__992 (.H(net992));
 TIEHIx1_ASAP7_75t_R _35467__993 (.H(net993));
 TIEHIx1_ASAP7_75t_R _35468__994 (.H(net994));
 TIEHIx1_ASAP7_75t_R _35469__995 (.H(net995));
 TIEHIx1_ASAP7_75t_R _35470__996 (.H(net996));
 TIEHIx1_ASAP7_75t_R _35471__997 (.H(net997));
 TIEHIx1_ASAP7_75t_R _35472__998 (.H(net998));
 TIEHIx1_ASAP7_75t_R _35473__999 (.H(net999));
 TIEHIx1_ASAP7_75t_R _35474__1000 (.H(net1000));
 TIEHIx1_ASAP7_75t_R _35475__1001 (.H(net1001));
 TIEHIx1_ASAP7_75t_R _35476__1002 (.H(net1002));
 TIEHIx1_ASAP7_75t_R _35477__1003 (.H(net1003));
 TIEHIx1_ASAP7_75t_R _35478__1004 (.H(net1004));
 TIEHIx1_ASAP7_75t_R _35479__1005 (.H(net1005));
 TIEHIx1_ASAP7_75t_R _35480__1006 (.H(net1006));
 TIEHIx1_ASAP7_75t_R _35481__1007 (.H(net1007));
 TIEHIx1_ASAP7_75t_R _35482__1008 (.H(net1008));
 TIEHIx1_ASAP7_75t_R _35483__1009 (.H(net1009));
 TIEHIx1_ASAP7_75t_R _35484__1010 (.H(net1010));
 TIEHIx1_ASAP7_75t_R _35485__1011 (.H(net1011));
 TIEHIx1_ASAP7_75t_R _35486__1012 (.H(net1012));
 TIEHIx1_ASAP7_75t_R _35487__1013 (.H(net1013));
 TIEHIx1_ASAP7_75t_R _35488__1014 (.H(net1014));
 TIEHIx1_ASAP7_75t_R _35489__1015 (.H(net1015));
 TIEHIx1_ASAP7_75t_R _35490__1016 (.H(net1016));
 TIEHIx1_ASAP7_75t_R _35491__1017 (.H(net1017));
 TIEHIx1_ASAP7_75t_R _35492__1018 (.H(net1018));
 TIEHIx1_ASAP7_75t_R _35493__1019 (.H(net1019));
 TIEHIx1_ASAP7_75t_R _35494__1020 (.H(net1020));
 TIEHIx1_ASAP7_75t_R _35495__1021 (.H(net1021));
 TIEHIx1_ASAP7_75t_R _35496__1022 (.H(net1022));
 TIEHIx1_ASAP7_75t_R _35497__1023 (.H(net1023));
 TIEHIx1_ASAP7_75t_R _35498__1024 (.H(net1024));
 TIEHIx1_ASAP7_75t_R _35499__1025 (.H(net1025));
 TIEHIx1_ASAP7_75t_R _35500__1026 (.H(net1026));
 TIEHIx1_ASAP7_75t_R _35501__1027 (.H(net1027));
 TIEHIx1_ASAP7_75t_R _35502__1028 (.H(net1028));
 TIEHIx1_ASAP7_75t_R _35503__1029 (.H(net1029));
 TIEHIx1_ASAP7_75t_R _35504__1030 (.H(net1030));
 TIEHIx1_ASAP7_75t_R _35505__1031 (.H(net1031));
 TIEHIx1_ASAP7_75t_R _35506__1032 (.H(net1032));
 TIEHIx1_ASAP7_75t_R _35507__1033 (.H(net1033));
 TIEHIx1_ASAP7_75t_R _35508__1034 (.H(net1034));
 TIEHIx1_ASAP7_75t_R _35509__1035 (.H(net1035));
 TIEHIx1_ASAP7_75t_R _35510__1036 (.H(net1036));
 TIEHIx1_ASAP7_75t_R _35511__1037 (.H(net1037));
 TIEHIx1_ASAP7_75t_R _35512__1038 (.H(net1038));
 TIEHIx1_ASAP7_75t_R _35513__1039 (.H(net1039));
 TIEHIx1_ASAP7_75t_R _35514__1040 (.H(net1040));
 TIEHIx1_ASAP7_75t_R _35515__1041 (.H(net1041));
 TIEHIx1_ASAP7_75t_R _35516__1042 (.H(net1042));
 TIEHIx1_ASAP7_75t_R _35517__1043 (.H(net1043));
 TIEHIx1_ASAP7_75t_R _35518__1044 (.H(net1044));
 TIEHIx1_ASAP7_75t_R _35519__1045 (.H(net1045));
 TIEHIx1_ASAP7_75t_R _35520__1046 (.H(net1046));
 TIEHIx1_ASAP7_75t_R _35521__1047 (.H(net1047));
 TIEHIx1_ASAP7_75t_R _35522__1048 (.H(net1048));
 TIEHIx1_ASAP7_75t_R _35523__1049 (.H(net1049));
 TIEHIx1_ASAP7_75t_R _35524__1050 (.H(net1050));
 TIEHIx1_ASAP7_75t_R _35525__1051 (.H(net1051));
 TIEHIx1_ASAP7_75t_R _35526__1052 (.H(net1052));
 TIEHIx1_ASAP7_75t_R _35527__1053 (.H(net1053));
 TIEHIx1_ASAP7_75t_R _35528__1054 (.H(net1054));
 TIEHIx1_ASAP7_75t_R _35529__1055 (.H(net1055));
 TIEHIx1_ASAP7_75t_R _35530__1056 (.H(net1056));
 TIEHIx1_ASAP7_75t_R _35531__1057 (.H(net1057));
 TIEHIx1_ASAP7_75t_R _35532__1058 (.H(net1058));
 TIEHIx1_ASAP7_75t_R _35533__1059 (.H(net1059));
 TIEHIx1_ASAP7_75t_R _35534__1060 (.H(net1060));
 TIEHIx1_ASAP7_75t_R _35535__1061 (.H(net1061));
 TIEHIx1_ASAP7_75t_R _35536__1062 (.H(net1062));
 TIEHIx1_ASAP7_75t_R _35537__1063 (.H(net1063));
 TIEHIx1_ASAP7_75t_R _35538__1064 (.H(net1064));
 TIEHIx1_ASAP7_75t_R _35539__1065 (.H(net1065));
 TIEHIx1_ASAP7_75t_R _35540__1066 (.H(net1066));
 TIEHIx1_ASAP7_75t_R _35541__1067 (.H(net1067));
 TIEHIx1_ASAP7_75t_R _35542__1068 (.H(net1068));
 TIEHIx1_ASAP7_75t_R _35543__1069 (.H(net1069));
 TIEHIx1_ASAP7_75t_R _35544__1070 (.H(net1070));
 TIEHIx1_ASAP7_75t_R _35545__1071 (.H(net1071));
 TIEHIx1_ASAP7_75t_R _35546__1072 (.H(net1072));
 TIEHIx1_ASAP7_75t_R _35547__1073 (.H(net1073));
 TIEHIx1_ASAP7_75t_R _35548__1074 (.H(net1074));
 TIEHIx1_ASAP7_75t_R _35549__1075 (.H(net1075));
 TIEHIx1_ASAP7_75t_R _35550__1076 (.H(net1076));
 TIEHIx1_ASAP7_75t_R _35551__1077 (.H(net1077));
 TIEHIx1_ASAP7_75t_R _35552__1078 (.H(net1078));
 TIEHIx1_ASAP7_75t_R _35553__1079 (.H(net1079));
 TIEHIx1_ASAP7_75t_R _35554__1080 (.H(net1080));
 TIEHIx1_ASAP7_75t_R _35555__1081 (.H(net1081));
 TIEHIx1_ASAP7_75t_R _35556__1082 (.H(net1082));
 TIEHIx1_ASAP7_75t_R _35557__1083 (.H(net1083));
 TIEHIx1_ASAP7_75t_R _35558__1084 (.H(net1084));
 TIEHIx1_ASAP7_75t_R _35559__1085 (.H(net1085));
 TIEHIx1_ASAP7_75t_R _35560__1086 (.H(net1086));
 TIEHIx1_ASAP7_75t_R _35561__1087 (.H(net1087));
 TIEHIx1_ASAP7_75t_R _35562__1088 (.H(net1088));
 TIEHIx1_ASAP7_75t_R _35563__1089 (.H(net1089));
 TIEHIx1_ASAP7_75t_R _35564__1090 (.H(net1090));
 TIEHIx1_ASAP7_75t_R _35565__1091 (.H(net1091));
 TIEHIx1_ASAP7_75t_R _35566__1092 (.H(net1092));
 TIEHIx1_ASAP7_75t_R _35567__1093 (.H(net1093));
 TIEHIx1_ASAP7_75t_R _35568__1094 (.H(net1094));
 TIEHIx1_ASAP7_75t_R _35569__1095 (.H(net1095));
 TIEHIx1_ASAP7_75t_R _35570__1096 (.H(net1096));
 TIEHIx1_ASAP7_75t_R _35571__1097 (.H(net1097));
 TIEHIx1_ASAP7_75t_R _35572__1098 (.H(net1098));
 TIEHIx1_ASAP7_75t_R _35573__1099 (.H(net1099));
 TIEHIx1_ASAP7_75t_R _35574__1100 (.H(net1100));
 TIEHIx1_ASAP7_75t_R _35575__1101 (.H(net1101));
 TIEHIx1_ASAP7_75t_R _35576__1102 (.H(net1102));
 TIEHIx1_ASAP7_75t_R _35577__1103 (.H(net1103));
 TIEHIx1_ASAP7_75t_R _35578__1104 (.H(net1104));
 TIEHIx1_ASAP7_75t_R _35579__1105 (.H(net1105));
 TIEHIx1_ASAP7_75t_R _35580__1106 (.H(net1106));
 TIEHIx1_ASAP7_75t_R _35581__1107 (.H(net1107));
 TIEHIx1_ASAP7_75t_R _35582__1108 (.H(net1108));
 TIEHIx1_ASAP7_75t_R _35583__1109 (.H(net1109));
 TIEHIx1_ASAP7_75t_R _35584__1110 (.H(net1110));
 TIEHIx1_ASAP7_75t_R _35585__1111 (.H(net1111));
 TIEHIx1_ASAP7_75t_R _35586__1112 (.H(net1112));
 TIEHIx1_ASAP7_75t_R _35587__1113 (.H(net1113));
 TIEHIx1_ASAP7_75t_R _35588__1114 (.H(net1114));
 TIEHIx1_ASAP7_75t_R _35589__1115 (.H(net1115));
 TIEHIx1_ASAP7_75t_R _35590__1116 (.H(net1116));
 TIEHIx1_ASAP7_75t_R _35591__1117 (.H(net1117));
 TIEHIx1_ASAP7_75t_R _35592__1118 (.H(net1118));
 TIEHIx1_ASAP7_75t_R _35593__1119 (.H(net1119));
 TIEHIx1_ASAP7_75t_R _35594__1120 (.H(net1120));
 TIEHIx1_ASAP7_75t_R _35595__1121 (.H(net1121));
 TIEHIx1_ASAP7_75t_R _35596__1122 (.H(net1122));
 TIEHIx1_ASAP7_75t_R _35597__1123 (.H(net1123));
 TIEHIx1_ASAP7_75t_R _35598__1124 (.H(net1124));
 TIEHIx1_ASAP7_75t_R _35599__1125 (.H(net1125));
 TIEHIx1_ASAP7_75t_R _35600__1126 (.H(net1126));
 TIEHIx1_ASAP7_75t_R _35601__1127 (.H(net1127));
 TIEHIx1_ASAP7_75t_R _35602__1128 (.H(net1128));
 TIEHIx1_ASAP7_75t_R _35603__1129 (.H(net1129));
 TIEHIx1_ASAP7_75t_R _35604__1130 (.H(net1130));
 TIEHIx1_ASAP7_75t_R _35605__1131 (.H(net1131));
 TIEHIx1_ASAP7_75t_R _35606__1132 (.H(net1132));
 TIEHIx1_ASAP7_75t_R _35607__1133 (.H(net1133));
 TIEHIx1_ASAP7_75t_R _35608__1134 (.H(net1134));
 TIEHIx1_ASAP7_75t_R _35609__1135 (.H(net1135));
 TIEHIx1_ASAP7_75t_R _35610__1136 (.H(net1136));
 TIEHIx1_ASAP7_75t_R _35611__1137 (.H(net1137));
 TIEHIx1_ASAP7_75t_R _35612__1138 (.H(net1138));
 TIEHIx1_ASAP7_75t_R _35613__1139 (.H(net1139));
 TIEHIx1_ASAP7_75t_R _35614__1140 (.H(net1140));
 TIEHIx1_ASAP7_75t_R _35615__1141 (.H(net1141));
 TIEHIx1_ASAP7_75t_R _35616__1142 (.H(net1142));
 TIEHIx1_ASAP7_75t_R _35617__1143 (.H(net1143));
 TIEHIx1_ASAP7_75t_R _35618__1144 (.H(net1144));
 TIEHIx1_ASAP7_75t_R _35619__1145 (.H(net1145));
 TIEHIx1_ASAP7_75t_R _35620__1146 (.H(net1146));
 TIEHIx1_ASAP7_75t_R _35621__1147 (.H(net1147));
 TIEHIx1_ASAP7_75t_R _35622__1148 (.H(net1148));
 TIEHIx1_ASAP7_75t_R _35623__1149 (.H(net1149));
 TIEHIx1_ASAP7_75t_R _35624__1150 (.H(net1150));
 TIEHIx1_ASAP7_75t_R _35625__1151 (.H(net1151));
 TIEHIx1_ASAP7_75t_R _35626__1152 (.H(net1152));
 TIEHIx1_ASAP7_75t_R _35627__1153 (.H(net1153));
 TIEHIx1_ASAP7_75t_R _35628__1154 (.H(net1154));
 TIEHIx1_ASAP7_75t_R _35629__1155 (.H(net1155));
 TIEHIx1_ASAP7_75t_R _35630__1156 (.H(net1156));
 TIEHIx1_ASAP7_75t_R _35631__1157 (.H(net1157));
 TIEHIx1_ASAP7_75t_R _35632__1158 (.H(net1158));
 TIEHIx1_ASAP7_75t_R _35633__1159 (.H(net1159));
 TIEHIx1_ASAP7_75t_R _35634__1160 (.H(net1160));
 TIEHIx1_ASAP7_75t_R _35635__1161 (.H(net1161));
 TIEHIx1_ASAP7_75t_R _35636__1162 (.H(net1162));
 TIEHIx1_ASAP7_75t_R _35637__1163 (.H(net1163));
 TIEHIx1_ASAP7_75t_R _35638__1164 (.H(net1164));
 TIEHIx1_ASAP7_75t_R _35639__1165 (.H(net1165));
 TIEHIx1_ASAP7_75t_R _35640__1166 (.H(net1166));
 TIEHIx1_ASAP7_75t_R _35641__1167 (.H(net1167));
 TIEHIx1_ASAP7_75t_R _35642__1168 (.H(net1168));
 TIEHIx1_ASAP7_75t_R _35643__1169 (.H(net1169));
 TIEHIx1_ASAP7_75t_R _35644__1170 (.H(net1170));
 TIEHIx1_ASAP7_75t_R _35645__1171 (.H(net1171));
 TIEHIx1_ASAP7_75t_R _35646__1172 (.H(net1172));
 TIEHIx1_ASAP7_75t_R _35647__1173 (.H(net1173));
 TIEHIx1_ASAP7_75t_R _35648__1174 (.H(net1174));
 TIEHIx1_ASAP7_75t_R _35649__1175 (.H(net1175));
 TIEHIx1_ASAP7_75t_R _35650__1176 (.H(net1176));
 TIEHIx1_ASAP7_75t_R _35651__1177 (.H(net1177));
 TIEHIx1_ASAP7_75t_R _35652__1178 (.H(net1178));
 TIEHIx1_ASAP7_75t_R _35653__1179 (.H(net1179));
 TIEHIx1_ASAP7_75t_R _35654__1180 (.H(net1180));
 TIEHIx1_ASAP7_75t_R _35655__1181 (.H(net1181));
 TIEHIx1_ASAP7_75t_R _35656__1182 (.H(net1182));
 TIEHIx1_ASAP7_75t_R _35657__1183 (.H(net1183));
 TIEHIx1_ASAP7_75t_R _35658__1184 (.H(net1184));
 TIEHIx1_ASAP7_75t_R _35659__1185 (.H(net1185));
 TIEHIx1_ASAP7_75t_R _35660__1186 (.H(net1186));
 TIEHIx1_ASAP7_75t_R _35661__1187 (.H(net1187));
 TIEHIx1_ASAP7_75t_R _35662__1188 (.H(net1188));
 TIEHIx1_ASAP7_75t_R _35663__1189 (.H(net1189));
 TIEHIx1_ASAP7_75t_R _35664__1190 (.H(net1190));
 TIEHIx1_ASAP7_75t_R _35665__1191 (.H(net1191));
 TIEHIx1_ASAP7_75t_R _35666__1192 (.H(net1192));
 TIEHIx1_ASAP7_75t_R _35667__1193 (.H(net1193));
 TIEHIx1_ASAP7_75t_R _35668__1194 (.H(net1194));
 TIEHIx1_ASAP7_75t_R _35669__1195 (.H(net1195));
 TIEHIx1_ASAP7_75t_R _35670__1196 (.H(net1196));
 TIEHIx1_ASAP7_75t_R _35671__1197 (.H(net1197));
 TIEHIx1_ASAP7_75t_R _35672__1198 (.H(net1198));
 TIEHIx1_ASAP7_75t_R _35673__1199 (.H(net1199));
 TIEHIx1_ASAP7_75t_R _35674__1200 (.H(net1200));
 TIEHIx1_ASAP7_75t_R _35675__1201 (.H(net1201));
 TIEHIx1_ASAP7_75t_R _35676__1202 (.H(net1202));
 TIEHIx1_ASAP7_75t_R _35677__1203 (.H(net1203));
 TIEHIx1_ASAP7_75t_R _35678__1204 (.H(net1204));
 TIEHIx1_ASAP7_75t_R _35679__1205 (.H(net1205));
 TIEHIx1_ASAP7_75t_R _35680__1206 (.H(net1206));
 TIEHIx1_ASAP7_75t_R _35681__1207 (.H(net1207));
 TIEHIx1_ASAP7_75t_R _35682__1208 (.H(net1208));
 TIEHIx1_ASAP7_75t_R _35683__1209 (.H(net1209));
 TIEHIx1_ASAP7_75t_R _35684__1210 (.H(net1210));
 TIEHIx1_ASAP7_75t_R _35685__1211 (.H(net1211));
 TIEHIx1_ASAP7_75t_R _35686__1212 (.H(net1212));
 TIEHIx1_ASAP7_75t_R _35687__1213 (.H(net1213));
 TIEHIx1_ASAP7_75t_R _35688__1214 (.H(net1214));
 TIEHIx1_ASAP7_75t_R _35689__1215 (.H(net1215));
 TIEHIx1_ASAP7_75t_R _35690__1216 (.H(net1216));
 TIEHIx1_ASAP7_75t_R _35691__1217 (.H(net1217));
 TIEHIx1_ASAP7_75t_R _35692__1218 (.H(net1218));
 TIEHIx1_ASAP7_75t_R _35693__1219 (.H(net1219));
 TIEHIx1_ASAP7_75t_R _35694__1220 (.H(net1220));
 TIEHIx1_ASAP7_75t_R _35695__1221 (.H(net1221));
 TIEHIx1_ASAP7_75t_R _35696__1222 (.H(net1222));
 TIEHIx1_ASAP7_75t_R _35697__1223 (.H(net1223));
 TIEHIx1_ASAP7_75t_R _35698__1224 (.H(net1224));
 TIEHIx1_ASAP7_75t_R _35699__1225 (.H(net1225));
 TIEHIx1_ASAP7_75t_R _35700__1226 (.H(net1226));
 TIEHIx1_ASAP7_75t_R _35701__1227 (.H(net1227));
 TIEHIx1_ASAP7_75t_R _35702__1228 (.H(net1228));
 TIEHIx1_ASAP7_75t_R _35703__1229 (.H(net1229));
 TIEHIx1_ASAP7_75t_R _35704__1230 (.H(net1230));
 TIEHIx1_ASAP7_75t_R _35705__1231 (.H(net1231));
 TIEHIx1_ASAP7_75t_R _35706__1232 (.H(net1232));
 TIEHIx1_ASAP7_75t_R _35707__1233 (.H(net1233));
 TIEHIx1_ASAP7_75t_R _35708__1234 (.H(net1234));
 TIEHIx1_ASAP7_75t_R _35709__1235 (.H(net1235));
 TIEHIx1_ASAP7_75t_R _35710__1236 (.H(net1236));
 TIEHIx1_ASAP7_75t_R _35711__1237 (.H(net1237));
 TIEHIx1_ASAP7_75t_R _35712__1238 (.H(net1238));
 TIEHIx1_ASAP7_75t_R _35713__1239 (.H(net1239));
 TIEHIx1_ASAP7_75t_R _35714__1240 (.H(net1240));
 TIEHIx1_ASAP7_75t_R _35715__1241 (.H(net1241));
 TIEHIx1_ASAP7_75t_R _35716__1242 (.H(net1242));
 TIEHIx1_ASAP7_75t_R _35717__1243 (.H(net1243));
 TIEHIx1_ASAP7_75t_R _35718__1244 (.H(net1244));
 TIEHIx1_ASAP7_75t_R _35719__1245 (.H(net1245));
 TIEHIx1_ASAP7_75t_R _35720__1246 (.H(net1246));
 TIEHIx1_ASAP7_75t_R _35721__1247 (.H(net1247));
 TIEHIx1_ASAP7_75t_R _35722__1248 (.H(net1248));
 TIEHIx1_ASAP7_75t_R _35723__1249 (.H(net1249));
 TIEHIx1_ASAP7_75t_R _35724__1250 (.H(net1250));
 TIEHIx1_ASAP7_75t_R _35725__1251 (.H(net1251));
 TIEHIx1_ASAP7_75t_R _35726__1252 (.H(net1252));
 TIEHIx1_ASAP7_75t_R _35727__1253 (.H(net1253));
 TIEHIx1_ASAP7_75t_R _35728__1254 (.H(net1254));
 TIEHIx1_ASAP7_75t_R _35729__1255 (.H(net1255));
 TIEHIx1_ASAP7_75t_R _35730__1256 (.H(net1256));
 TIEHIx1_ASAP7_75t_R _35731__1257 (.H(net1257));
 TIEHIx1_ASAP7_75t_R _35732__1258 (.H(net1258));
 TIEHIx1_ASAP7_75t_R _35733__1259 (.H(net1259));
 TIEHIx1_ASAP7_75t_R _35734__1260 (.H(net1260));
 TIEHIx1_ASAP7_75t_R _35735__1261 (.H(net1261));
 TIEHIx1_ASAP7_75t_R _35736__1262 (.H(net1262));
 TIEHIx1_ASAP7_75t_R _35737__1263 (.H(net1263));
 TIEHIx1_ASAP7_75t_R _35738__1264 (.H(net1264));
 TIEHIx1_ASAP7_75t_R _35739__1265 (.H(net1265));
 TIEHIx1_ASAP7_75t_R _35740__1266 (.H(net1266));
 TIEHIx1_ASAP7_75t_R _35741__1267 (.H(net1267));
 TIEHIx1_ASAP7_75t_R _35742__1268 (.H(net1268));
 TIEHIx1_ASAP7_75t_R _35743__1269 (.H(net1269));
 TIEHIx1_ASAP7_75t_R _35744__1270 (.H(net1270));
 TIEHIx1_ASAP7_75t_R _35745__1271 (.H(net1271));
 TIEHIx1_ASAP7_75t_R _35746__1272 (.H(net1272));
 TIEHIx1_ASAP7_75t_R _35747__1273 (.H(net1273));
 TIEHIx1_ASAP7_75t_R _35748__1274 (.H(net1274));
 TIEHIx1_ASAP7_75t_R _35749__1275 (.H(net1275));
 TIEHIx1_ASAP7_75t_R _35750__1276 (.H(net1276));
 TIEHIx1_ASAP7_75t_R _35751__1277 (.H(net1277));
 TIEHIx1_ASAP7_75t_R _35752__1278 (.H(net1278));
 TIEHIx1_ASAP7_75t_R _35753__1279 (.H(net1279));
 TIEHIx1_ASAP7_75t_R _35754__1280 (.H(net1280));
 TIEHIx1_ASAP7_75t_R _35755__1281 (.H(net1281));
 TIEHIx1_ASAP7_75t_R _35756__1282 (.H(net1282));
 TIEHIx1_ASAP7_75t_R _35757__1283 (.H(net1283));
 TIEHIx1_ASAP7_75t_R _35758__1284 (.H(net1284));
 TIEHIx1_ASAP7_75t_R _35759__1285 (.H(net1285));
 TIEHIx1_ASAP7_75t_R _35760__1286 (.H(net1286));
 TIEHIx1_ASAP7_75t_R _35761__1287 (.H(net1287));
 TIEHIx1_ASAP7_75t_R _35762__1288 (.H(net1288));
 TIEHIx1_ASAP7_75t_R _35763__1289 (.H(net1289));
 TIEHIx1_ASAP7_75t_R _35764__1290 (.H(net1290));
 TIEHIx1_ASAP7_75t_R _35765__1291 (.H(net1291));
 TIEHIx1_ASAP7_75t_R _35766__1292 (.H(net1292));
 TIEHIx1_ASAP7_75t_R _35767__1293 (.H(net1293));
 TIEHIx1_ASAP7_75t_R _35768__1294 (.H(net1294));
 TIEHIx1_ASAP7_75t_R _35769__1295 (.H(net1295));
 TIEHIx1_ASAP7_75t_R _35770__1296 (.H(net1296));
 TIEHIx1_ASAP7_75t_R _35771__1297 (.H(net1297));
 TIEHIx1_ASAP7_75t_R _35772__1298 (.H(net1298));
 TIEHIx1_ASAP7_75t_R _35773__1299 (.H(net1299));
 TIEHIx1_ASAP7_75t_R _35774__1300 (.H(net1300));
 TIEHIx1_ASAP7_75t_R _35775__1301 (.H(net1301));
 TIEHIx1_ASAP7_75t_R _35776__1302 (.H(net1302));
 TIEHIx1_ASAP7_75t_R _35777__1303 (.H(net1303));
 TIEHIx1_ASAP7_75t_R _35778__1304 (.H(net1304));
 TIEHIx1_ASAP7_75t_R _35779__1305 (.H(net1305));
 TIEHIx1_ASAP7_75t_R _35780__1306 (.H(net1306));
 TIEHIx1_ASAP7_75t_R _35781__1307 (.H(net1307));
 TIEHIx1_ASAP7_75t_R _35782__1308 (.H(net1308));
 TIEHIx1_ASAP7_75t_R _35783__1309 (.H(net1309));
 TIEHIx1_ASAP7_75t_R _35784__1310 (.H(net1310));
 TIEHIx1_ASAP7_75t_R _35785__1311 (.H(net1311));
 TIEHIx1_ASAP7_75t_R _35786__1312 (.H(net1312));
 TIEHIx1_ASAP7_75t_R _35787__1313 (.H(net1313));
 TIEHIx1_ASAP7_75t_R _35788__1314 (.H(net1314));
 TIEHIx1_ASAP7_75t_R _35789__1315 (.H(net1315));
 TIEHIx1_ASAP7_75t_R _35790__1316 (.H(net1316));
 TIEHIx1_ASAP7_75t_R _35791__1317 (.H(net1317));
 TIEHIx1_ASAP7_75t_R _35792__1318 (.H(net1318));
 TIEHIx1_ASAP7_75t_R _35793__1319 (.H(net1319));
 TIEHIx1_ASAP7_75t_R _35794__1320 (.H(net1320));
 TIEHIx1_ASAP7_75t_R _35795__1321 (.H(net1321));
 TIEHIx1_ASAP7_75t_R _35796__1322 (.H(net1322));
 TIEHIx1_ASAP7_75t_R _35797__1323 (.H(net1323));
 TIEHIx1_ASAP7_75t_R _35798__1324 (.H(net1324));
 TIEHIx1_ASAP7_75t_R _35799__1325 (.H(net1325));
 TIEHIx1_ASAP7_75t_R _35800__1326 (.H(net1326));
 TIEHIx1_ASAP7_75t_R _35801__1327 (.H(net1327));
 TIEHIx1_ASAP7_75t_R _35802__1328 (.H(net1328));
 TIEHIx1_ASAP7_75t_R _35803__1329 (.H(net1329));
 TIEHIx1_ASAP7_75t_R _35804__1330 (.H(net1330));
 TIEHIx1_ASAP7_75t_R _35805__1331 (.H(net1331));
 TIEHIx1_ASAP7_75t_R _35806__1332 (.H(net1332));
 TIEHIx1_ASAP7_75t_R _35807__1333 (.H(net1333));
 TIEHIx1_ASAP7_75t_R _35808__1334 (.H(net1334));
 TIEHIx1_ASAP7_75t_R _35809__1335 (.H(net1335));
 TIEHIx1_ASAP7_75t_R _35810__1336 (.H(net1336));
 TIEHIx1_ASAP7_75t_R _35811__1337 (.H(net1337));
 TIEHIx1_ASAP7_75t_R _35812__1338 (.H(net1338));
 TIEHIx1_ASAP7_75t_R _35813__1339 (.H(net1339));
 TIEHIx1_ASAP7_75t_R _35814__1340 (.H(net1340));
 TIEHIx1_ASAP7_75t_R _35815__1341 (.H(net1341));
 TIEHIx1_ASAP7_75t_R _35816__1342 (.H(net1342));
 TIEHIx1_ASAP7_75t_R _35817__1343 (.H(net1343));
 TIEHIx1_ASAP7_75t_R _35818__1344 (.H(net1344));
 TIEHIx1_ASAP7_75t_R _35819__1345 (.H(net1345));
 TIEHIx1_ASAP7_75t_R _35820__1346 (.H(net1346));
 TIEHIx1_ASAP7_75t_R _35821__1347 (.H(net1347));
 TIEHIx1_ASAP7_75t_R _35822__1348 (.H(net1348));
 TIEHIx1_ASAP7_75t_R _35823__1349 (.H(net1349));
 TIEHIx1_ASAP7_75t_R _35824__1350 (.H(net1350));
 TIEHIx1_ASAP7_75t_R _35825__1351 (.H(net1351));
 TIEHIx1_ASAP7_75t_R _35826__1352 (.H(net1352));
 TIEHIx1_ASAP7_75t_R _35827__1353 (.H(net1353));
 TIEHIx1_ASAP7_75t_R _35828__1354 (.H(net1354));
 TIEHIx1_ASAP7_75t_R _35829__1355 (.H(net1355));
 TIEHIx1_ASAP7_75t_R _35830__1356 (.H(net1356));
 TIEHIx1_ASAP7_75t_R _35831__1357 (.H(net1357));
 TIEHIx1_ASAP7_75t_R _35832__1358 (.H(net1358));
 TIEHIx1_ASAP7_75t_R _35833__1359 (.H(net1359));
 TIEHIx1_ASAP7_75t_R _35834__1360 (.H(net1360));
 TIEHIx1_ASAP7_75t_R _35835__1361 (.H(net1361));
 TIEHIx1_ASAP7_75t_R _35836__1362 (.H(net1362));
 TIEHIx1_ASAP7_75t_R _35837__1363 (.H(net1363));
 TIEHIx1_ASAP7_75t_R _35838__1364 (.H(net1364));
 TIEHIx1_ASAP7_75t_R _35839__1365 (.H(net1365));
 TIEHIx1_ASAP7_75t_R _35840__1366 (.H(net1366));
 TIEHIx1_ASAP7_75t_R _35841__1367 (.H(net1367));
 TIEHIx1_ASAP7_75t_R _35842__1368 (.H(net1368));
 TIEHIx1_ASAP7_75t_R _35843__1369 (.H(net1369));
 TIEHIx1_ASAP7_75t_R _35844__1370 (.H(net1370));
 TIEHIx1_ASAP7_75t_R _35845__1371 (.H(net1371));
 TIEHIx1_ASAP7_75t_R _35846__1372 (.H(net1372));
 TIEHIx1_ASAP7_75t_R _35847__1373 (.H(net1373));
 TIEHIx1_ASAP7_75t_R _35848__1374 (.H(net1374));
 TIEHIx1_ASAP7_75t_R _35849__1375 (.H(net1375));
 TIEHIx1_ASAP7_75t_R _35850__1376 (.H(net1376));
 TIEHIx1_ASAP7_75t_R _35851__1377 (.H(net1377));
 TIEHIx1_ASAP7_75t_R _35852__1378 (.H(net1378));
 TIEHIx1_ASAP7_75t_R _35853__1379 (.H(net1379));
 TIEHIx1_ASAP7_75t_R _35854__1380 (.H(net1380));
 TIEHIx1_ASAP7_75t_R _35855__1381 (.H(net1381));
 TIEHIx1_ASAP7_75t_R _35856__1382 (.H(net1382));
 TIEHIx1_ASAP7_75t_R _35857__1383 (.H(net1383));
 TIEHIx1_ASAP7_75t_R _35858__1384 (.H(net1384));
 TIEHIx1_ASAP7_75t_R _35859__1385 (.H(net1385));
 TIEHIx1_ASAP7_75t_R _35860__1386 (.H(net1386));
 TIEHIx1_ASAP7_75t_R _35861__1387 (.H(net1387));
 TIEHIx1_ASAP7_75t_R _35862__1388 (.H(net1388));
 TIEHIx1_ASAP7_75t_R _35863__1389 (.H(net1389));
 TIEHIx1_ASAP7_75t_R _35864__1390 (.H(net1390));
 TIEHIx1_ASAP7_75t_R _35865__1391 (.H(net1391));
 TIEHIx1_ASAP7_75t_R _35866__1392 (.H(net1392));
 TIEHIx1_ASAP7_75t_R _35867__1393 (.H(net1393));
 TIEHIx1_ASAP7_75t_R _35868__1394 (.H(net1394));
 TIEHIx1_ASAP7_75t_R _35869__1395 (.H(net1395));
 TIEHIx1_ASAP7_75t_R _35870__1396 (.H(net1396));
 TIEHIx1_ASAP7_75t_R _35871__1397 (.H(net1397));
 TIEHIx1_ASAP7_75t_R _35872__1398 (.H(net1398));
 TIEHIx1_ASAP7_75t_R _35873__1399 (.H(net1399));
 TIEHIx1_ASAP7_75t_R _35874__1400 (.H(net1400));
 TIEHIx1_ASAP7_75t_R _35875__1401 (.H(net1401));
 TIEHIx1_ASAP7_75t_R _35876__1402 (.H(net1402));
 TIEHIx1_ASAP7_75t_R _35877__1403 (.H(net1403));
 TIEHIx1_ASAP7_75t_R _35878__1404 (.H(net1404));
 TIEHIx1_ASAP7_75t_R _35879__1405 (.H(net1405));
 TIEHIx1_ASAP7_75t_R _35880__1406 (.H(net1406));
 TIEHIx1_ASAP7_75t_R _35881__1407 (.H(net1407));
 TIEHIx1_ASAP7_75t_R _35882__1408 (.H(net1408));
 TIEHIx1_ASAP7_75t_R _35883__1409 (.H(net1409));
 TIEHIx1_ASAP7_75t_R _35884__1410 (.H(net1410));
 TIEHIx1_ASAP7_75t_R _35885__1411 (.H(net1411));
 TIEHIx1_ASAP7_75t_R _35886__1412 (.H(net1412));
 TIEHIx1_ASAP7_75t_R _35887__1413 (.H(net1413));
 TIEHIx1_ASAP7_75t_R _35888__1414 (.H(net1414));
 TIEHIx1_ASAP7_75t_R _35889__1415 (.H(net1415));
 TIEHIx1_ASAP7_75t_R _35890__1416 (.H(net1416));
 TIEHIx1_ASAP7_75t_R _35891__1417 (.H(net1417));
 TIEHIx1_ASAP7_75t_R _35892__1418 (.H(net1418));
 TIEHIx1_ASAP7_75t_R _35893__1419 (.H(net1419));
 TIEHIx1_ASAP7_75t_R _35894__1420 (.H(net1420));
 TIEHIx1_ASAP7_75t_R _35895__1421 (.H(net1421));
 TIEHIx1_ASAP7_75t_R _35896__1422 (.H(net1422));
 TIEHIx1_ASAP7_75t_R _35897__1423 (.H(net1423));
 TIEHIx1_ASAP7_75t_R _35898__1424 (.H(net1424));
 TIEHIx1_ASAP7_75t_R _35899__1425 (.H(net1425));
 TIEHIx1_ASAP7_75t_R _35900__1426 (.H(net1426));
 TIEHIx1_ASAP7_75t_R _35901__1427 (.H(net1427));
 TIEHIx1_ASAP7_75t_R _35902__1428 (.H(net1428));
 TIEHIx1_ASAP7_75t_R _35903__1429 (.H(net1429));
 TIEHIx1_ASAP7_75t_R _35904__1430 (.H(net1430));
 TIEHIx1_ASAP7_75t_R _35905__1431 (.H(net1431));
 TIEHIx1_ASAP7_75t_R _35906__1432 (.H(net1432));
 TIEHIx1_ASAP7_75t_R _35907__1433 (.H(net1433));
 TIEHIx1_ASAP7_75t_R _35908__1434 (.H(net1434));
 TIEHIx1_ASAP7_75t_R _35909__1435 (.H(net1435));
 TIEHIx1_ASAP7_75t_R _35910__1436 (.H(net1436));
 TIEHIx1_ASAP7_75t_R _35911__1437 (.H(net1437));
 TIEHIx1_ASAP7_75t_R _35912__1438 (.H(net1438));
 TIEHIx1_ASAP7_75t_R _35913__1439 (.H(net1439));
 TIEHIx1_ASAP7_75t_R _35914__1440 (.H(net1440));
 TIEHIx1_ASAP7_75t_R _35915__1441 (.H(net1441));
 TIEHIx1_ASAP7_75t_R _35916__1442 (.H(net1442));
 TIEHIx1_ASAP7_75t_R _35917__1443 (.H(net1443));
 TIEHIx1_ASAP7_75t_R _35918__1444 (.H(net1444));
 TIEHIx1_ASAP7_75t_R _35919__1445 (.H(net1445));
 TIEHIx1_ASAP7_75t_R _35920__1446 (.H(net1446));
 TIEHIx1_ASAP7_75t_R _35921__1447 (.H(net1447));
 TIEHIx1_ASAP7_75t_R _35922__1448 (.H(net1448));
 TIEHIx1_ASAP7_75t_R _35923__1449 (.H(net1449));
 TIEHIx1_ASAP7_75t_R _35924__1450 (.H(net1450));
 TIEHIx1_ASAP7_75t_R _35925__1451 (.H(net1451));
 TIEHIx1_ASAP7_75t_R _35926__1452 (.H(net1452));
 TIEHIx1_ASAP7_75t_R _35927__1453 (.H(net1453));
 TIEHIx1_ASAP7_75t_R _35928__1454 (.H(net1454));
 TIEHIx1_ASAP7_75t_R _35929__1455 (.H(net1455));
 TIEHIx1_ASAP7_75t_R _35930__1456 (.H(net1456));
 TIEHIx1_ASAP7_75t_R _35931__1457 (.H(net1457));
 TIEHIx1_ASAP7_75t_R _35932__1458 (.H(net1458));
 TIEHIx1_ASAP7_75t_R _35933__1459 (.H(net1459));
 TIEHIx1_ASAP7_75t_R _35934__1460 (.H(net1460));
 TIEHIx1_ASAP7_75t_R _35935__1461 (.H(net1461));
 TIEHIx1_ASAP7_75t_R _35936__1462 (.H(net1462));
 TIEHIx1_ASAP7_75t_R _35937__1463 (.H(net1463));
 TIEHIx1_ASAP7_75t_R _35938__1464 (.H(net1464));
 TIEHIx1_ASAP7_75t_R _35939__1465 (.H(net1465));
 TIEHIx1_ASAP7_75t_R _35940__1466 (.H(net1466));
 TIEHIx1_ASAP7_75t_R _35941__1467 (.H(net1467));
 TIEHIx1_ASAP7_75t_R _35942__1468 (.H(net1468));
 TIEHIx1_ASAP7_75t_R _35943__1469 (.H(net1469));
 TIEHIx1_ASAP7_75t_R _35944__1470 (.H(net1470));
 TIEHIx1_ASAP7_75t_R _35945__1471 (.H(net1471));
 TIEHIx1_ASAP7_75t_R _35946__1472 (.H(net1472));
 TIEHIx1_ASAP7_75t_R _35947__1473 (.H(net1473));
 TIEHIx1_ASAP7_75t_R _35948__1474 (.H(net1474));
 TIEHIx1_ASAP7_75t_R _35949__1475 (.H(net1475));
 TIEHIx1_ASAP7_75t_R _35950__1476 (.H(net1476));
 TIEHIx1_ASAP7_75t_R _35951__1477 (.H(net1477));
 TIEHIx1_ASAP7_75t_R _35952__1478 (.H(net1478));
 TIEHIx1_ASAP7_75t_R _35953__1479 (.H(net1479));
 TIEHIx1_ASAP7_75t_R _35954__1480 (.H(net1480));
 TIEHIx1_ASAP7_75t_R _35955__1481 (.H(net1481));
 TIEHIx1_ASAP7_75t_R _35956__1482 (.H(net1482));
 TIEHIx1_ASAP7_75t_R _35957__1483 (.H(net1483));
 TIEHIx1_ASAP7_75t_R _35958__1484 (.H(net1484));
 TIEHIx1_ASAP7_75t_R _35959__1485 (.H(net1485));
 TIEHIx1_ASAP7_75t_R _35960__1486 (.H(net1486));
 TIEHIx1_ASAP7_75t_R _35961__1487 (.H(net1487));
 TIEHIx1_ASAP7_75t_R _35962__1488 (.H(net1488));
 TIEHIx1_ASAP7_75t_R _35963__1489 (.H(net1489));
 TIEHIx1_ASAP7_75t_R _35964__1490 (.H(net1490));
 TIEHIx1_ASAP7_75t_R _35965__1491 (.H(net1491));
 TIEHIx1_ASAP7_75t_R _35966__1492 (.H(net1492));
 TIEHIx1_ASAP7_75t_R _35967__1493 (.H(net1493));
 TIEHIx1_ASAP7_75t_R _35968__1494 (.H(net1494));
 TIEHIx1_ASAP7_75t_R _35969__1495 (.H(net1495));
 TIEHIx1_ASAP7_75t_R _35970__1496 (.H(net1496));
 TIEHIx1_ASAP7_75t_R _35971__1497 (.H(net1497));
 TIEHIx1_ASAP7_75t_R _35972__1498 (.H(net1498));
 TIEHIx1_ASAP7_75t_R _35973__1499 (.H(net1499));
 TIEHIx1_ASAP7_75t_R _35974__1500 (.H(net1500));
 TIEHIx1_ASAP7_75t_R _35975__1501 (.H(net1501));
 TIEHIx1_ASAP7_75t_R _35976__1502 (.H(net1502));
 TIEHIx1_ASAP7_75t_R _35977__1503 (.H(net1503));
 TIEHIx1_ASAP7_75t_R _35978__1504 (.H(net1504));
 TIEHIx1_ASAP7_75t_R _35979__1505 (.H(net1505));
 TIEHIx1_ASAP7_75t_R _35980__1506 (.H(net1506));
 TIEHIx1_ASAP7_75t_R _35981__1507 (.H(net1507));
 TIEHIx1_ASAP7_75t_R _35982__1508 (.H(net1508));
 TIEHIx1_ASAP7_75t_R _35983__1509 (.H(net1509));
 TIEHIx1_ASAP7_75t_R _35984__1510 (.H(net1510));
 TIEHIx1_ASAP7_75t_R _35985__1511 (.H(net1511));
 TIEHIx1_ASAP7_75t_R _35986__1512 (.H(net1512));
 TIEHIx1_ASAP7_75t_R _35987__1513 (.H(net1513));
 TIEHIx1_ASAP7_75t_R _35988__1514 (.H(net1514));
 TIEHIx1_ASAP7_75t_R _35989__1515 (.H(net1515));
 TIEHIx1_ASAP7_75t_R _35990__1516 (.H(net1516));
 TIEHIx1_ASAP7_75t_R _35991__1517 (.H(net1517));
 TIEHIx1_ASAP7_75t_R _35992__1518 (.H(net1518));
 TIEHIx1_ASAP7_75t_R _35993__1519 (.H(net1519));
 TIEHIx1_ASAP7_75t_R _35994__1520 (.H(net1520));
 TIEHIx1_ASAP7_75t_R _35995__1521 (.H(net1521));
 TIEHIx1_ASAP7_75t_R _35996__1522 (.H(net1522));
 TIEHIx1_ASAP7_75t_R _35997__1523 (.H(net1523));
 TIEHIx1_ASAP7_75t_R _35998__1524 (.H(net1524));
 TIEHIx1_ASAP7_75t_R _35999__1525 (.H(net1525));
 TIEHIx1_ASAP7_75t_R _36000__1526 (.H(net1526));
 TIEHIx1_ASAP7_75t_R _36001__1527 (.H(net1527));
 TIEHIx1_ASAP7_75t_R _36002__1528 (.H(net1528));
 TIEHIx1_ASAP7_75t_R _36003__1529 (.H(net1529));
 TIEHIx1_ASAP7_75t_R _36004__1530 (.H(net1530));
 TIEHIx1_ASAP7_75t_R _36005__1531 (.H(net1531));
 TIEHIx1_ASAP7_75t_R _36006__1532 (.H(net1532));
 TIEHIx1_ASAP7_75t_R _36007__1533 (.H(net1533));
 TIEHIx1_ASAP7_75t_R _36008__1534 (.H(net1534));
 TIEHIx1_ASAP7_75t_R _36009__1535 (.H(net1535));
 TIEHIx1_ASAP7_75t_R _36010__1536 (.H(net1536));
 TIEHIx1_ASAP7_75t_R _36011__1537 (.H(net1537));
 TIEHIx1_ASAP7_75t_R _36012__1538 (.H(net1538));
 TIEHIx1_ASAP7_75t_R _36013__1539 (.H(net1539));
 TIEHIx1_ASAP7_75t_R _36014__1540 (.H(net1540));
 TIEHIx1_ASAP7_75t_R _36015__1541 (.H(net1541));
 TIEHIx1_ASAP7_75t_R _36016__1542 (.H(net1542));
 TIEHIx1_ASAP7_75t_R _36017__1543 (.H(net1543));
 TIEHIx1_ASAP7_75t_R _36018__1544 (.H(net1544));
 TIEHIx1_ASAP7_75t_R _36019__1545 (.H(net1545));
 TIEHIx1_ASAP7_75t_R _36020__1546 (.H(net1546));
 TIEHIx1_ASAP7_75t_R _36021__1547 (.H(net1547));
 TIEHIx1_ASAP7_75t_R _36022__1548 (.H(net1548));
 TIEHIx1_ASAP7_75t_R _36023__1549 (.H(net1549));
 TIEHIx1_ASAP7_75t_R _36024__1550 (.H(net1550));
 TIEHIx1_ASAP7_75t_R _36025__1551 (.H(net1551));
 TIEHIx1_ASAP7_75t_R _36026__1552 (.H(net1552));
 TIEHIx1_ASAP7_75t_R _36027__1553 (.H(net1553));
 TIEHIx1_ASAP7_75t_R _36028__1554 (.H(net1554));
 TIEHIx1_ASAP7_75t_R _36029__1555 (.H(net1555));
 TIEHIx1_ASAP7_75t_R _36030__1556 (.H(net1556));
 TIEHIx1_ASAP7_75t_R _36031__1557 (.H(net1557));
 TIEHIx1_ASAP7_75t_R _36032__1558 (.H(net1558));
 TIEHIx1_ASAP7_75t_R _36033__1559 (.H(net1559));
 TIEHIx1_ASAP7_75t_R _36034__1560 (.H(net1560));
 TIEHIx1_ASAP7_75t_R _36035__1561 (.H(net1561));
 TIEHIx1_ASAP7_75t_R _36036__1562 (.H(net1562));
 TIEHIx1_ASAP7_75t_R _36037__1563 (.H(net1563));
 TIEHIx1_ASAP7_75t_R _36038__1564 (.H(net1564));
 TIEHIx1_ASAP7_75t_R _36039__1565 (.H(net1565));
 TIEHIx1_ASAP7_75t_R _36040__1566 (.H(net1566));
 TIEHIx1_ASAP7_75t_R _36041__1567 (.H(net1567));
 TIEHIx1_ASAP7_75t_R _36042__1568 (.H(net1568));
 TIEHIx1_ASAP7_75t_R _36043__1569 (.H(net1569));
 TIEHIx1_ASAP7_75t_R _36044__1570 (.H(net1570));
 TIEHIx1_ASAP7_75t_R _36045__1571 (.H(net1571));
 TIEHIx1_ASAP7_75t_R _36046__1572 (.H(net1572));
 TIEHIx1_ASAP7_75t_R _36047__1573 (.H(net1573));
 TIEHIx1_ASAP7_75t_R _36048__1574 (.H(net1574));
 TIEHIx1_ASAP7_75t_R _36049__1575 (.H(net1575));
 TIEHIx1_ASAP7_75t_R _36050__1576 (.H(net1576));
 TIEHIx1_ASAP7_75t_R _36051__1577 (.H(net1577));
 TIEHIx1_ASAP7_75t_R _36052__1578 (.H(net1578));
 TIEHIx1_ASAP7_75t_R _36053__1579 (.H(net1579));
 TIEHIx1_ASAP7_75t_R _36054__1580 (.H(net1580));
 TIEHIx1_ASAP7_75t_R _36055__1581 (.H(net1581));
 TIEHIx1_ASAP7_75t_R _36056__1582 (.H(net1582));
 TIEHIx1_ASAP7_75t_R _36057__1583 (.H(net1583));
 TIEHIx1_ASAP7_75t_R _36058__1584 (.H(net1584));
 TIEHIx1_ASAP7_75t_R _36059__1585 (.H(net1585));
 TIEHIx1_ASAP7_75t_R _36060__1586 (.H(net1586));
 TIEHIx1_ASAP7_75t_R _36061__1587 (.H(net1587));
 TIEHIx1_ASAP7_75t_R _36062__1588 (.H(net1588));
 TIEHIx1_ASAP7_75t_R _36063__1589 (.H(net1589));
 TIEHIx1_ASAP7_75t_R _36064__1590 (.H(net1590));
 TIEHIx1_ASAP7_75t_R _36065__1591 (.H(net1591));
 TIEHIx1_ASAP7_75t_R _36066__1592 (.H(net1592));
 TIEHIx1_ASAP7_75t_R _36067__1593 (.H(net1593));
 TIEHIx1_ASAP7_75t_R _36068__1594 (.H(net1594));
 TIEHIx1_ASAP7_75t_R _36069__1595 (.H(net1595));
 TIEHIx1_ASAP7_75t_R _36070__1596 (.H(net1596));
 TIEHIx1_ASAP7_75t_R _36071__1597 (.H(net1597));
 TIEHIx1_ASAP7_75t_R _36072__1598 (.H(net1598));
 TIEHIx1_ASAP7_75t_R _36073__1599 (.H(net1599));
 TIEHIx1_ASAP7_75t_R _36074__1600 (.H(net1600));
 TIEHIx1_ASAP7_75t_R _36075__1601 (.H(net1601));
 TIEHIx1_ASAP7_75t_R _36076__1602 (.H(net1602));
 TIEHIx1_ASAP7_75t_R _36077__1603 (.H(net1603));
 TIEHIx1_ASAP7_75t_R _36078__1604 (.H(net1604));
 TIEHIx1_ASAP7_75t_R _36079__1605 (.H(net1605));
 TIEHIx1_ASAP7_75t_R _36080__1606 (.H(net1606));
 TIEHIx1_ASAP7_75t_R _36081__1607 (.H(net1607));
 TIEHIx1_ASAP7_75t_R _36082__1608 (.H(net1608));
 TIEHIx1_ASAP7_75t_R _36083__1609 (.H(net1609));
 TIEHIx1_ASAP7_75t_R _36084__1610 (.H(net1610));
 TIEHIx1_ASAP7_75t_R _36085__1611 (.H(net1611));
 TIEHIx1_ASAP7_75t_R _36086__1612 (.H(net1612));
 TIEHIx1_ASAP7_75t_R _36087__1613 (.H(net1613));
 TIEHIx1_ASAP7_75t_R _36088__1614 (.H(net1614));
 TIEHIx1_ASAP7_75t_R _36089__1615 (.H(net1615));
 TIEHIx1_ASAP7_75t_R _36090__1616 (.H(net1616));
 TIEHIx1_ASAP7_75t_R _36091__1617 (.H(net1617));
 TIEHIx1_ASAP7_75t_R _36092__1618 (.H(net1618));
 TIEHIx1_ASAP7_75t_R _36093__1619 (.H(net1619));
 TIEHIx1_ASAP7_75t_R _36094__1620 (.H(net1620));
 TIEHIx1_ASAP7_75t_R _36095__1621 (.H(net1621));
 TIEHIx1_ASAP7_75t_R _36096__1622 (.H(net1622));
 TIEHIx1_ASAP7_75t_R _36097__1623 (.H(net1623));
 TIEHIx1_ASAP7_75t_R _36098__1624 (.H(net1624));
 TIEHIx1_ASAP7_75t_R _36099__1625 (.H(net1625));
 TIEHIx1_ASAP7_75t_R _36100__1626 (.H(net1626));
 TIEHIx1_ASAP7_75t_R _36101__1627 (.H(net1627));
 TIEHIx1_ASAP7_75t_R _36102__1628 (.H(net1628));
 TIEHIx1_ASAP7_75t_R _36103__1629 (.H(net1629));
 TIEHIx1_ASAP7_75t_R _36104__1630 (.H(net1630));
 TIEHIx1_ASAP7_75t_R _36105__1631 (.H(net1631));
 TIEHIx1_ASAP7_75t_R _36106__1632 (.H(net1632));
 TIEHIx1_ASAP7_75t_R _36107__1633 (.H(net1633));
 TIEHIx1_ASAP7_75t_R _36108__1634 (.H(net1634));
 TIEHIx1_ASAP7_75t_R _36109__1635 (.H(net1635));
 TIEHIx1_ASAP7_75t_R _36110__1636 (.H(net1636));
 TIEHIx1_ASAP7_75t_R _36111__1637 (.H(net1637));
 TIEHIx1_ASAP7_75t_R _36112__1638 (.H(net1638));
 TIEHIx1_ASAP7_75t_R _36113__1639 (.H(net1639));
 TIEHIx1_ASAP7_75t_R _36114__1640 (.H(net1640));
 TIEHIx1_ASAP7_75t_R _36115__1641 (.H(net1641));
 TIEHIx1_ASAP7_75t_R _36116__1642 (.H(net1642));
 TIEHIx1_ASAP7_75t_R _36117__1643 (.H(net1643));
 TIEHIx1_ASAP7_75t_R _36118__1644 (.H(net1644));
 TIEHIx1_ASAP7_75t_R _36119__1645 (.H(net1645));
 TIEHIx1_ASAP7_75t_R _36120__1646 (.H(net1646));
 TIEHIx1_ASAP7_75t_R _36121__1647 (.H(net1647));
 TIEHIx1_ASAP7_75t_R _36122__1648 (.H(net1648));
 TIEHIx1_ASAP7_75t_R _36123__1649 (.H(net1649));
 TIEHIx1_ASAP7_75t_R _36124__1650 (.H(net1650));
 TIEHIx1_ASAP7_75t_R _36125__1651 (.H(net1651));
 TIEHIx1_ASAP7_75t_R _36126__1652 (.H(net1652));
 TIEHIx1_ASAP7_75t_R _36127__1653 (.H(net1653));
 TIEHIx1_ASAP7_75t_R _36128__1654 (.H(net1654));
 TIEHIx1_ASAP7_75t_R _36129__1655 (.H(net1655));
 TIEHIx1_ASAP7_75t_R _36130__1656 (.H(net1656));
 TIEHIx1_ASAP7_75t_R _36131__1657 (.H(net1657));
 TIEHIx1_ASAP7_75t_R _36132__1658 (.H(net1658));
 TIEHIx1_ASAP7_75t_R _36133__1659 (.H(net1659));
 TIEHIx1_ASAP7_75t_R _36134__1660 (.H(net1660));
 TIEHIx1_ASAP7_75t_R _36135__1661 (.H(net1661));
 TIEHIx1_ASAP7_75t_R _36136__1662 (.H(net1662));
 TIEHIx1_ASAP7_75t_R _36137__1663 (.H(net1663));
 TIEHIx1_ASAP7_75t_R _36138__1664 (.H(net1664));
 TIEHIx1_ASAP7_75t_R _36139__1665 (.H(net1665));
 TIEHIx1_ASAP7_75t_R _36140__1666 (.H(net1666));
 TIEHIx1_ASAP7_75t_R _36141__1667 (.H(net1667));
 TIEHIx1_ASAP7_75t_R _36142__1668 (.H(net1668));
 TIEHIx1_ASAP7_75t_R _36143__1669 (.H(net1669));
 TIEHIx1_ASAP7_75t_R _36144__1670 (.H(net1670));
 TIEHIx1_ASAP7_75t_R _36145__1671 (.H(net1671));
 TIEHIx1_ASAP7_75t_R _36146__1672 (.H(net1672));
 TIEHIx1_ASAP7_75t_R _36147__1673 (.H(net1673));
 TIEHIx1_ASAP7_75t_R _36148__1674 (.H(net1674));
 TIEHIx1_ASAP7_75t_R _36149__1675 (.H(net1675));
 TIEHIx1_ASAP7_75t_R _36150__1676 (.H(net1676));
 TIEHIx1_ASAP7_75t_R _36151__1677 (.H(net1677));
 TIEHIx1_ASAP7_75t_R _36152__1678 (.H(net1678));
 TIEHIx1_ASAP7_75t_R _36153__1679 (.H(net1679));
 TIEHIx1_ASAP7_75t_R _36154__1680 (.H(net1680));
 TIEHIx1_ASAP7_75t_R _36155__1681 (.H(net1681));
 TIEHIx1_ASAP7_75t_R _36156__1682 (.H(net1682));
 TIEHIx1_ASAP7_75t_R _36157__1683 (.H(net1683));
 TIEHIx1_ASAP7_75t_R _36158__1684 (.H(net1684));
 TIEHIx1_ASAP7_75t_R _36159__1685 (.H(net1685));
 TIEHIx1_ASAP7_75t_R _36160__1686 (.H(net1686));
 TIEHIx1_ASAP7_75t_R _36161__1687 (.H(net1687));
 TIEHIx1_ASAP7_75t_R _36162__1688 (.H(net1688));
 TIEHIx1_ASAP7_75t_R _36163__1689 (.H(net1689));
 TIEHIx1_ASAP7_75t_R _36164__1690 (.H(net1690));
 TIEHIx1_ASAP7_75t_R _36165__1691 (.H(net1691));
 TIEHIx1_ASAP7_75t_R _36166__1692 (.H(net1692));
 TIEHIx1_ASAP7_75t_R _36167__1693 (.H(net1693));
 TIEHIx1_ASAP7_75t_R _36168__1694 (.H(net1694));
 TIEHIx1_ASAP7_75t_R _36169__1695 (.H(net1695));
 TIEHIx1_ASAP7_75t_R _36170__1696 (.H(net1696));
 TIEHIx1_ASAP7_75t_R _36171__1697 (.H(net1697));
 TIEHIx1_ASAP7_75t_R _36172__1698 (.H(net1698));
 TIEHIx1_ASAP7_75t_R _36173__1699 (.H(net1699));
 TIEHIx1_ASAP7_75t_R _36174__1700 (.H(net1700));
 TIEHIx1_ASAP7_75t_R _36175__1701 (.H(net1701));
 TIEHIx1_ASAP7_75t_R _36176__1702 (.H(net1702));
 TIEHIx1_ASAP7_75t_R _36177__1703 (.H(net1703));
 TIEHIx1_ASAP7_75t_R _36178__1704 (.H(net1704));
 TIEHIx1_ASAP7_75t_R _36179__1705 (.H(net1705));
 TIEHIx1_ASAP7_75t_R _36180__1706 (.H(net1706));
 TIEHIx1_ASAP7_75t_R _36181__1707 (.H(net1707));
 TIEHIx1_ASAP7_75t_R _36182__1708 (.H(net1708));
 TIEHIx1_ASAP7_75t_R _36183__1709 (.H(net1709));
 TIEHIx1_ASAP7_75t_R _36184__1710 (.H(net1710));
 TIEHIx1_ASAP7_75t_R _36185__1711 (.H(net1711));
 TIEHIx1_ASAP7_75t_R _36186__1712 (.H(net1712));
 TIEHIx1_ASAP7_75t_R _36187__1713 (.H(net1713));
 TIEHIx1_ASAP7_75t_R _36188__1714 (.H(net1714));
 TIEHIx1_ASAP7_75t_R _36189__1715 (.H(net1715));
 TIEHIx1_ASAP7_75t_R _36190__1716 (.H(net1716));
 TIEHIx1_ASAP7_75t_R _36191__1717 (.H(net1717));
 TIEHIx1_ASAP7_75t_R _36192__1718 (.H(net1718));
 TIEHIx1_ASAP7_75t_R _36193__1719 (.H(net1719));
 TIEHIx1_ASAP7_75t_R _36194__1720 (.H(net1720));
 TIEHIx1_ASAP7_75t_R _36195__1721 (.H(net1721));
 TIEHIx1_ASAP7_75t_R _36196__1722 (.H(net1722));
 TIEHIx1_ASAP7_75t_R _36197__1723 (.H(net1723));
 TIEHIx1_ASAP7_75t_R _36198__1724 (.H(net1724));
 TIEHIx1_ASAP7_75t_R _36199__1725 (.H(net1725));
 TIEHIx1_ASAP7_75t_R _36200__1726 (.H(net1726));
 TIEHIx1_ASAP7_75t_R _36201__1727 (.H(net1727));
 TIEHIx1_ASAP7_75t_R _36202__1728 (.H(net1728));
 TIEHIx1_ASAP7_75t_R _36203__1729 (.H(net1729));
 TIEHIx1_ASAP7_75t_R _36204__1730 (.H(net1730));
 TIEHIx1_ASAP7_75t_R _36205__1731 (.H(net1731));
 TIEHIx1_ASAP7_75t_R _36206__1732 (.H(net1732));
 TIEHIx1_ASAP7_75t_R _36207__1733 (.H(net1733));
 TIEHIx1_ASAP7_75t_R _36208__1734 (.H(net1734));
 TIEHIx1_ASAP7_75t_R _36209__1735 (.H(net1735));
 TIEHIx1_ASAP7_75t_R _36210__1736 (.H(net1736));
 TIEHIx1_ASAP7_75t_R _36211__1737 (.H(net1737));
 TIEHIx1_ASAP7_75t_R _36212__1738 (.H(net1738));
 TIEHIx1_ASAP7_75t_R _36213__1739 (.H(net1739));
 TIEHIx1_ASAP7_75t_R _36214__1740 (.H(net1740));
 TIEHIx1_ASAP7_75t_R _36215__1741 (.H(net1741));
 TIEHIx1_ASAP7_75t_R _36216__1742 (.H(net1742));
 TIEHIx1_ASAP7_75t_R _36217__1743 (.H(net1743));
 TIEHIx1_ASAP7_75t_R _36218__1744 (.H(net1744));
 TIEHIx1_ASAP7_75t_R _36219__1745 (.H(net1745));
 TIEHIx1_ASAP7_75t_R _36220__1746 (.H(net1746));
 TIEHIx1_ASAP7_75t_R _36221__1747 (.H(net1747));
 TIEHIx1_ASAP7_75t_R _36222__1748 (.H(net1748));
 TIEHIx1_ASAP7_75t_R _36223__1749 (.H(net1749));
 TIEHIx1_ASAP7_75t_R _36224__1750 (.H(net1750));
 TIEHIx1_ASAP7_75t_R _36225__1751 (.H(net1751));
 TIEHIx1_ASAP7_75t_R _36226__1752 (.H(net1752));
 TIEHIx1_ASAP7_75t_R _36227__1753 (.H(net1753));
 TIEHIx1_ASAP7_75t_R _36228__1754 (.H(net1754));
 TIEHIx1_ASAP7_75t_R _36229__1755 (.H(net1755));
 TIEHIx1_ASAP7_75t_R _36260__1756 (.H(net1756));
 TIEHIx1_ASAP7_75t_R _36261__1757 (.H(net1757));
 TIEHIx1_ASAP7_75t_R _36262__1758 (.H(net1758));
 TIEHIx1_ASAP7_75t_R _36263__1759 (.H(net1759));
 TIEHIx1_ASAP7_75t_R _36264__1760 (.H(net1760));
 TIEHIx1_ASAP7_75t_R _36265__1761 (.H(net1761));
 TIEHIx1_ASAP7_75t_R _36266__1762 (.H(net1762));
 TIEHIx1_ASAP7_75t_R _36267__1763 (.H(net1763));
 TIEHIx1_ASAP7_75t_R _36268__1764 (.H(net1764));
 TIEHIx1_ASAP7_75t_R _36269__1765 (.H(net1765));
 TIEHIx1_ASAP7_75t_R _36270__1766 (.H(net1766));
 TIEHIx1_ASAP7_75t_R _36271__1767 (.H(net1767));
 TIEHIx1_ASAP7_75t_R _36272__1768 (.H(net1768));
 TIEHIx1_ASAP7_75t_R _36273__1769 (.H(net1769));
 TIEHIx1_ASAP7_75t_R _36274__1770 (.H(net1770));
 TIEHIx1_ASAP7_75t_R _36275__1771 (.H(net1771));
 TIEHIx1_ASAP7_75t_R _36276__1772 (.H(net1772));
 TIEHIx1_ASAP7_75t_R _36277__1773 (.H(net1773));
 TIEHIx1_ASAP7_75t_R _36278__1774 (.H(net1774));
 TIEHIx1_ASAP7_75t_R _36279__1775 (.H(net1775));
 TIEHIx1_ASAP7_75t_R _36280__1776 (.H(net1776));
 TIEHIx1_ASAP7_75t_R _36281__1777 (.H(net1777));
 TIEHIx1_ASAP7_75t_R _36282__1778 (.H(net1778));
 TIEHIx1_ASAP7_75t_R _36283__1779 (.H(net1779));
 TIEHIx1_ASAP7_75t_R _36284__1780 (.H(net1780));
 TIEHIx1_ASAP7_75t_R _36285__1781 (.H(net1781));
 TIEHIx1_ASAP7_75t_R _36286__1782 (.H(net1782));
 TIEHIx1_ASAP7_75t_R _36287__1783 (.H(net1783));
 TIEHIx1_ASAP7_75t_R _36288__1784 (.H(net1784));
 TIEHIx1_ASAP7_75t_R _36289__1785 (.H(net1785));
 TIEHIx1_ASAP7_75t_R _36290__1786 (.H(net1786));
 TIEHIx1_ASAP7_75t_R _36291__1787 (.H(net1787));
 TIEHIx1_ASAP7_75t_R _36292__1788 (.H(net1788));
 TIEHIx1_ASAP7_75t_R _36293__1789 (.H(net1789));
 TIEHIx1_ASAP7_75t_R _36294__1790 (.H(net1790));
 TIEHIx1_ASAP7_75t_R _36295__1791 (.H(net1791));
 TIEHIx1_ASAP7_75t_R _36296__1792 (.H(net1792));
 TIEHIx1_ASAP7_75t_R _36297__1793 (.H(net1793));
 TIEHIx1_ASAP7_75t_R _36298__1794 (.H(net1794));
 TIEHIx1_ASAP7_75t_R _36299__1795 (.H(net1795));
 TIEHIx1_ASAP7_75t_R _36300__1796 (.H(net1796));
 TIEHIx1_ASAP7_75t_R _36301__1797 (.H(net1797));
 TIEHIx1_ASAP7_75t_R _36302__1798 (.H(net1798));
 TIEHIx1_ASAP7_75t_R _36303__1799 (.H(net1799));
 TIEHIx1_ASAP7_75t_R _36304__1800 (.H(net1800));
 TIEHIx1_ASAP7_75t_R _36305__1801 (.H(net1801));
 TIEHIx1_ASAP7_75t_R _36306__1802 (.H(net1802));
 TIEHIx1_ASAP7_75t_R _36307__1803 (.H(net1803));
 TIEHIx1_ASAP7_75t_R _36308__1804 (.H(net1804));
 TIEHIx1_ASAP7_75t_R _36309__1805 (.H(net1805));
 TIEHIx1_ASAP7_75t_R _36310__1806 (.H(net1806));
 TIEHIx1_ASAP7_75t_R _36311__1807 (.H(net1807));
 TIEHIx1_ASAP7_75t_R _36312__1808 (.H(net1808));
 TIEHIx1_ASAP7_75t_R _36313__1809 (.H(net1809));
 TIEHIx1_ASAP7_75t_R _36314__1810 (.H(net1810));
 TIEHIx1_ASAP7_75t_R _36315__1811 (.H(net1811));
 TIEHIx1_ASAP7_75t_R _36316__1812 (.H(net1812));
 TIEHIx1_ASAP7_75t_R _36317__1813 (.H(net1813));
 TIEHIx1_ASAP7_75t_R _36318__1814 (.H(net1814));
 TIEHIx1_ASAP7_75t_R _36319__1815 (.H(net1815));
 TIEHIx1_ASAP7_75t_R _36320__1816 (.H(net1816));
 TIEHIx1_ASAP7_75t_R _36321__1817 (.H(net1817));
 TIEHIx1_ASAP7_75t_R _36322__1818 (.H(net1818));
 TIEHIx1_ASAP7_75t_R _36323__1819 (.H(net1819));
 TIEHIx1_ASAP7_75t_R _36324__1820 (.H(net1820));
 TIEHIx1_ASAP7_75t_R _36325__1821 (.H(net1821));
 TIEHIx1_ASAP7_75t_R _36326__1822 (.H(net1822));
 TIEHIx1_ASAP7_75t_R _36327__1823 (.H(net1823));
 TIEHIx1_ASAP7_75t_R _36328__1824 (.H(net1824));
 TIEHIx1_ASAP7_75t_R _36329__1825 (.H(net1825));
 TIEHIx1_ASAP7_75t_R _36330__1826 (.H(net1826));
 TIEHIx1_ASAP7_75t_R _36331__1827 (.H(net1827));
 TIEHIx1_ASAP7_75t_R _36332__1828 (.H(net1828));
 TIEHIx1_ASAP7_75t_R _36333__1829 (.H(net1829));
 TIEHIx1_ASAP7_75t_R _36334__1830 (.H(net1830));
 TIEHIx1_ASAP7_75t_R _36335__1831 (.H(net1831));
 TIEHIx1_ASAP7_75t_R _36336__1832 (.H(net1832));
 TIEHIx1_ASAP7_75t_R _36337__1833 (.H(net1833));
 TIEHIx1_ASAP7_75t_R _36338__1834 (.H(net1834));
 TIEHIx1_ASAP7_75t_R _36339__1835 (.H(net1835));
 TIEHIx1_ASAP7_75t_R _36340__1836 (.H(net1836));
 TIEHIx1_ASAP7_75t_R _36341__1837 (.H(net1837));
 TIEHIx1_ASAP7_75t_R _36342__1838 (.H(net1838));
 TIEHIx1_ASAP7_75t_R _36343__1839 (.H(net1839));
 TIEHIx1_ASAP7_75t_R _36344__1840 (.H(net1840));
 TIEHIx1_ASAP7_75t_R _36345__1841 (.H(net1841));
 TIEHIx1_ASAP7_75t_R _36346__1842 (.H(net1842));
 TIEHIx1_ASAP7_75t_R _36347__1843 (.H(net1843));
 TIEHIx1_ASAP7_75t_R _36348__1844 (.H(net1844));
 TIEHIx1_ASAP7_75t_R _36349__1845 (.H(net1845));
 TIEHIx1_ASAP7_75t_R _36350__1846 (.H(net1846));
 TIEHIx1_ASAP7_75t_R _36351__1847 (.H(net1847));
 TIEHIx1_ASAP7_75t_R _36352__1848 (.H(net1848));
 TIEHIx1_ASAP7_75t_R _36353__1849 (.H(net1849));
 TIEHIx1_ASAP7_75t_R _36354__1850 (.H(net1850));
 TIEHIx1_ASAP7_75t_R _36355__1851 (.H(net1851));
 TIEHIx1_ASAP7_75t_R _36356__1852 (.H(net1852));
 TIEHIx1_ASAP7_75t_R _36357__1853 (.H(net1853));
 TIEHIx1_ASAP7_75t_R _36358__1854 (.H(net1854));
 TIEHIx1_ASAP7_75t_R _36359__1855 (.H(net1855));
 TIEHIx1_ASAP7_75t_R _36360__1856 (.H(net1856));
 TIEHIx1_ASAP7_75t_R _36361__1857 (.H(net1857));
 TIEHIx1_ASAP7_75t_R _36362__1858 (.H(net1858));
 TIEHIx1_ASAP7_75t_R _36363__1859 (.H(net1859));
 TIEHIx1_ASAP7_75t_R _36364__1860 (.H(net1860));
 TIEHIx1_ASAP7_75t_R _36365__1861 (.H(net1861));
 TIEHIx1_ASAP7_75t_R _36366__1862 (.H(net1862));
 TIEHIx1_ASAP7_75t_R _36367__1863 (.H(net1863));
 TIEHIx1_ASAP7_75t_R _36368__1864 (.H(net1864));
 TIEHIx1_ASAP7_75t_R _36369__1865 (.H(net1865));
 TIEHIx1_ASAP7_75t_R _36370__1866 (.H(net1866));
 TIEHIx1_ASAP7_75t_R _36371__1867 (.H(net1867));
 TIEHIx1_ASAP7_75t_R _36372__1868 (.H(net1868));
 TIEHIx1_ASAP7_75t_R _36373__1869 (.H(net1869));
 TIEHIx1_ASAP7_75t_R _36374__1870 (.H(net1870));
 TIEHIx1_ASAP7_75t_R _36375__1871 (.H(net1871));
 TIEHIx1_ASAP7_75t_R _36376__1872 (.H(net1872));
 TIEHIx1_ASAP7_75t_R _36377__1873 (.H(net1873));
 TIEHIx1_ASAP7_75t_R _36378__1874 (.H(net1874));
 TIEHIx1_ASAP7_75t_R _36379__1875 (.H(net1875));
 TIEHIx1_ASAP7_75t_R _36380__1876 (.H(net1876));
 TIEHIx1_ASAP7_75t_R _36381__1877 (.H(net1877));
 TIEHIx1_ASAP7_75t_R _36382__1878 (.H(net1878));
 TIEHIx1_ASAP7_75t_R _36383__1879 (.H(net1879));
 TIEHIx1_ASAP7_75t_R _36384__1880 (.H(net1880));
 TIEHIx1_ASAP7_75t_R _36385__1881 (.H(net1881));
 TIEHIx1_ASAP7_75t_R _36386__1882 (.H(net1882));
 TIEHIx1_ASAP7_75t_R _36387__1883 (.H(net1883));
 TIEHIx1_ASAP7_75t_R _36388__1884 (.H(net1884));
 TIEHIx1_ASAP7_75t_R _36389__1885 (.H(net1885));
 TIEHIx1_ASAP7_75t_R _36390__1886 (.H(net1886));
 TIEHIx1_ASAP7_75t_R _36391__1887 (.H(net1887));
 TIEHIx1_ASAP7_75t_R _36392__1888 (.H(net1888));
 TIEHIx1_ASAP7_75t_R _36393__1889 (.H(net1889));
 TIEHIx1_ASAP7_75t_R _36394__1890 (.H(net1890));
 TIEHIx1_ASAP7_75t_R _36395__1891 (.H(net1891));
 TIEHIx1_ASAP7_75t_R _36396__1892 (.H(net1892));
 TIEHIx1_ASAP7_75t_R _36397__1893 (.H(net1893));
 TIEHIx1_ASAP7_75t_R _36398__1894 (.H(net1894));
 TIEHIx1_ASAP7_75t_R _36399__1895 (.H(net1895));
 TIEHIx1_ASAP7_75t_R _36400__1896 (.H(net1896));
 TIEHIx1_ASAP7_75t_R _36401__1897 (.H(net1897));
 TIEHIx1_ASAP7_75t_R _36402__1898 (.H(net1898));
 TIEHIx1_ASAP7_75t_R _36403__1899 (.H(net1899));
 TIEHIx1_ASAP7_75t_R _36404__1900 (.H(net1900));
 TIEHIx1_ASAP7_75t_R _36405__1901 (.H(net1901));
 TIEHIx1_ASAP7_75t_R _36406__1902 (.H(net1902));
 TIEHIx1_ASAP7_75t_R _36407__1903 (.H(net1903));
 TIEHIx1_ASAP7_75t_R _36408__1904 (.H(net1904));
 TIEHIx1_ASAP7_75t_R _36409__1905 (.H(net1905));
 TIEHIx1_ASAP7_75t_R _36410__1906 (.H(net1906));
 TIEHIx1_ASAP7_75t_R _36411__1907 (.H(net1907));
 TIEHIx1_ASAP7_75t_R _36412__1908 (.H(net1908));
 TIEHIx1_ASAP7_75t_R _36413__1909 (.H(net1909));
 TIEHIx1_ASAP7_75t_R _36414__1910 (.H(net1910));
 TIEHIx1_ASAP7_75t_R _36415__1911 (.H(net1911));
 TIEHIx1_ASAP7_75t_R _36416__1912 (.H(net1912));
 TIEHIx1_ASAP7_75t_R _36417__1913 (.H(net1913));
 TIEHIx1_ASAP7_75t_R _36418__1914 (.H(net1914));
 TIEHIx1_ASAP7_75t_R _36419__1915 (.H(net1915));
 TIEHIx1_ASAP7_75t_R _36420__1916 (.H(net1916));
 TIEHIx1_ASAP7_75t_R _36421__1917 (.H(net1917));
 TIEHIx1_ASAP7_75t_R _36422__1918 (.H(net1918));
 TIEHIx1_ASAP7_75t_R _36423__1919 (.H(net1919));
 TIEHIx1_ASAP7_75t_R _36424__1920 (.H(net1920));
 TIEHIx1_ASAP7_75t_R _36425__1921 (.H(net1921));
 TIEHIx1_ASAP7_75t_R _36426__1922 (.H(net1922));
 TIEHIx1_ASAP7_75t_R _36427__1923 (.H(net1923));
 TIEHIx1_ASAP7_75t_R _36428__1924 (.H(net1924));
 TIEHIx1_ASAP7_75t_R _36429__1925 (.H(net1925));
 TIEHIx1_ASAP7_75t_R _36430__1926 (.H(net1926));
 TIEHIx1_ASAP7_75t_R _36431__1927 (.H(net1927));
 TIEHIx1_ASAP7_75t_R _36432__1928 (.H(net1928));
 TIEHIx1_ASAP7_75t_R _36433__1929 (.H(net1929));
 TIEHIx1_ASAP7_75t_R _36434__1930 (.H(net1930));
 TIEHIx1_ASAP7_75t_R _36435__1931 (.H(net1931));
 TIEHIx1_ASAP7_75t_R _36436__1932 (.H(net1932));
 TIEHIx1_ASAP7_75t_R _36437__1933 (.H(net1933));
 TIEHIx1_ASAP7_75t_R _36438__1934 (.H(net1934));
 TIEHIx1_ASAP7_75t_R _36439__1935 (.H(net1935));
 TIEHIx1_ASAP7_75t_R _36440__1936 (.H(net1936));
 TIEHIx1_ASAP7_75t_R _36441__1937 (.H(net1937));
 TIEHIx1_ASAP7_75t_R _36442__1938 (.H(net1938));
 TIEHIx1_ASAP7_75t_R _36443__1939 (.H(net1939));
 TIEHIx1_ASAP7_75t_R _36444__1940 (.H(net1940));
 TIEHIx1_ASAP7_75t_R _36445__1941 (.H(net1941));
 TIEHIx1_ASAP7_75t_R _36446__1942 (.H(net1942));
 TIEHIx1_ASAP7_75t_R _36447__1943 (.H(net1943));
 TIEHIx1_ASAP7_75t_R _36448__1944 (.H(net1944));
 TIEHIx1_ASAP7_75t_R _36449__1945 (.H(net1945));
 TIEHIx1_ASAP7_75t_R _36450__1946 (.H(net1946));
 TIEHIx1_ASAP7_75t_R _36451__1947 (.H(net1947));
 TIEHIx1_ASAP7_75t_R _36452__1948 (.H(net1948));
 TIEHIx1_ASAP7_75t_R _36453__1949 (.H(net1949));
 TIEHIx1_ASAP7_75t_R _36454__1950 (.H(net1950));
 TIEHIx1_ASAP7_75t_R _36455__1951 (.H(net1951));
 TIEHIx1_ASAP7_75t_R _36456__1952 (.H(net1952));
 TIEHIx1_ASAP7_75t_R _36457__1953 (.H(net1953));
 TIEHIx1_ASAP7_75t_R _36458__1954 (.H(net1954));
 TIEHIx1_ASAP7_75t_R _36459__1955 (.H(net1955));
 TIEHIx1_ASAP7_75t_R _36460__1956 (.H(net1956));
 TIEHIx1_ASAP7_75t_R _36461__1957 (.H(net1957));
 TIEHIx1_ASAP7_75t_R _36462__1958 (.H(net1958));
 TIEHIx1_ASAP7_75t_R _36463__1959 (.H(net1959));
 TIEHIx1_ASAP7_75t_R _36464__1960 (.H(net1960));
 TIEHIx1_ASAP7_75t_R _36465__1961 (.H(net1961));
 TIEHIx1_ASAP7_75t_R _36466__1962 (.H(net1962));
 TIEHIx1_ASAP7_75t_R _36467__1963 (.H(net1963));
 TIEHIx1_ASAP7_75t_R _36468__1964 (.H(net1964));
 TIEHIx1_ASAP7_75t_R _36469__1965 (.H(net1965));
 TIEHIx1_ASAP7_75t_R _36470__1966 (.H(net1966));
 TIEHIx1_ASAP7_75t_R _36471__1967 (.H(net1967));
 TIEHIx1_ASAP7_75t_R _36472__1968 (.H(net1968));
 TIEHIx1_ASAP7_75t_R _36473__1969 (.H(net1969));
 TIEHIx1_ASAP7_75t_R _36474__1970 (.H(net1970));
 TIEHIx1_ASAP7_75t_R _36475__1971 (.H(net1971));
 TIEHIx1_ASAP7_75t_R _36476__1972 (.H(net1972));
 TIEHIx1_ASAP7_75t_R _36477__1973 (.H(net1973));
 TIEHIx1_ASAP7_75t_R _36478__1974 (.H(net1974));
 TIEHIx1_ASAP7_75t_R _36479__1975 (.H(net1975));
 TIEHIx1_ASAP7_75t_R _36480__1976 (.H(net1976));
 TIEHIx1_ASAP7_75t_R _36481__1977 (.H(net1977));
 TIEHIx1_ASAP7_75t_R _36482__1978 (.H(net1978));
 TIEHIx1_ASAP7_75t_R _36483__1979 (.H(net1979));
 TIEHIx1_ASAP7_75t_R _36484__1980 (.H(net1980));
 TIEHIx1_ASAP7_75t_R _36485__1981 (.H(net1981));
 TIEHIx1_ASAP7_75t_R _36486__1982 (.H(net1982));
 TIEHIx1_ASAP7_75t_R _36487__1983 (.H(net1983));
 TIEHIx1_ASAP7_75t_R _36488__1984 (.H(net1984));
 TIEHIx1_ASAP7_75t_R _36489__1985 (.H(net1985));
 TIEHIx1_ASAP7_75t_R _36490__1986 (.H(net1986));
 TIEHIx1_ASAP7_75t_R _36491__1987 (.H(net1987));
 TIEHIx1_ASAP7_75t_R _36492__1988 (.H(net1988));
 TIEHIx1_ASAP7_75t_R _36493__1989 (.H(net1989));
 TIEHIx1_ASAP7_75t_R _36494__1990 (.H(net1990));
 TIEHIx1_ASAP7_75t_R _36495__1991 (.H(net1991));
 TIEHIx1_ASAP7_75t_R _36496__1992 (.H(net1992));
 TIEHIx1_ASAP7_75t_R _36497__1993 (.H(net1993));
 TIEHIx1_ASAP7_75t_R _36498__1994 (.H(net1994));
 TIEHIx1_ASAP7_75t_R _36499__1995 (.H(net1995));
 TIEHIx1_ASAP7_75t_R _36500__1996 (.H(net1996));
 TIEHIx1_ASAP7_75t_R _36501__1997 (.H(net1997));
 TIEHIx1_ASAP7_75t_R _36502__1998 (.H(net1998));
 TIEHIx1_ASAP7_75t_R _36503__1999 (.H(net1999));
 TIEHIx1_ASAP7_75t_R _36504__2000 (.H(net2000));
 TIEHIx1_ASAP7_75t_R _36505__2001 (.H(net2001));
 TIEHIx1_ASAP7_75t_R _36506__2002 (.H(net2002));
 TIEHIx1_ASAP7_75t_R _36507__2003 (.H(net2003));
 TIEHIx1_ASAP7_75t_R _36508__2004 (.H(net2004));
 TIEHIx1_ASAP7_75t_R _36509__2005 (.H(net2005));
 TIEHIx1_ASAP7_75t_R _36510__2006 (.H(net2006));
 TIEHIx1_ASAP7_75t_R _36511__2007 (.H(net2007));
 TIEHIx1_ASAP7_75t_R _36512__2008 (.H(net2008));
 TIEHIx1_ASAP7_75t_R _36513__2009 (.H(net2009));
 TIEHIx1_ASAP7_75t_R _36514__2010 (.H(net2010));
 TIEHIx1_ASAP7_75t_R _36515__2011 (.H(net2011));
 TIEHIx1_ASAP7_75t_R _36516__2012 (.H(net2012));
 TIEHIx1_ASAP7_75t_R _36517__2013 (.H(net2013));
 TIEHIx1_ASAP7_75t_R _36518__2014 (.H(net2014));
 TIEHIx1_ASAP7_75t_R _36519__2015 (.H(net2015));
 TIEHIx1_ASAP7_75t_R _36520__2016 (.H(net2016));
 TIEHIx1_ASAP7_75t_R _36521__2017 (.H(net2017));
 TIEHIx1_ASAP7_75t_R _36522__2018 (.H(net2018));
 TIEHIx1_ASAP7_75t_R _36523__2019 (.H(net2019));
 TIEHIx1_ASAP7_75t_R _36524__2020 (.H(net2020));
 TIEHIx1_ASAP7_75t_R _36525__2021 (.H(net2021));
 TIEHIx1_ASAP7_75t_R _36526__2022 (.H(net2022));
 TIEHIx1_ASAP7_75t_R _36527__2023 (.H(net2023));
 TIEHIx1_ASAP7_75t_R _36528__2024 (.H(net2024));
 TIEHIx1_ASAP7_75t_R _36529__2025 (.H(net2025));
 TIEHIx1_ASAP7_75t_R _36530__2026 (.H(net2026));
 TIEHIx1_ASAP7_75t_R _36531__2027 (.H(net2027));
 TIEHIx1_ASAP7_75t_R _36532__2028 (.H(net2028));
 TIEHIx1_ASAP7_75t_R _36533__2029 (.H(net2029));
 TIEHIx1_ASAP7_75t_R _36534__2030 (.H(net2030));
 TIEHIx1_ASAP7_75t_R _36535__2031 (.H(net2031));
 TIEHIx1_ASAP7_75t_R _36536__2032 (.H(net2032));
 TIEHIx1_ASAP7_75t_R _36537__2033 (.H(net2033));
 TIEHIx1_ASAP7_75t_R _36538__2034 (.H(net2034));
 TIEHIx1_ASAP7_75t_R _36539__2035 (.H(net2035));
 TIEHIx1_ASAP7_75t_R _36540__2036 (.H(net2036));
 TIEHIx1_ASAP7_75t_R _36541__2037 (.H(net2037));
 TIEHIx1_ASAP7_75t_R _36542__2038 (.H(net2038));
 TIEHIx1_ASAP7_75t_R _36543__2039 (.H(net2039));
 TIEHIx1_ASAP7_75t_R _36544__2040 (.H(net2040));
 TIEHIx1_ASAP7_75t_R _36545__2041 (.H(net2041));
 TIEHIx1_ASAP7_75t_R _36546__2042 (.H(net2042));
 TIEHIx1_ASAP7_75t_R _36547__2043 (.H(net2043));
 TIEHIx1_ASAP7_75t_R _36548__2044 (.H(net2044));
 TIEHIx1_ASAP7_75t_R _36549__2045 (.H(net2045));
 TIEHIx1_ASAP7_75t_R _36550__2046 (.H(net2046));
 TIEHIx1_ASAP7_75t_R _36551__2047 (.H(net2047));
 TIEHIx1_ASAP7_75t_R _36552__2048 (.H(net2048));
 TIEHIx1_ASAP7_75t_R _36553__2049 (.H(net2049));
 TIEHIx1_ASAP7_75t_R _36554__2050 (.H(net2050));
 TIEHIx1_ASAP7_75t_R _36555__2051 (.H(net2051));
 TIEHIx1_ASAP7_75t_R _36556__2052 (.H(net2052));
 TIEHIx1_ASAP7_75t_R _36557__2053 (.H(net2053));
 TIEHIx1_ASAP7_75t_R _36558__2054 (.H(net2054));
 TIEHIx1_ASAP7_75t_R _36559__2055 (.H(net2055));
 TIEHIx1_ASAP7_75t_R _36560__2056 (.H(net2056));
 TIEHIx1_ASAP7_75t_R _36561__2057 (.H(net2057));
 TIEHIx1_ASAP7_75t_R _36562__2058 (.H(net2058));
 TIEHIx1_ASAP7_75t_R _36563__2059 (.H(net2059));
 TIEHIx1_ASAP7_75t_R _36564__2060 (.H(net2060));
 TIEHIx1_ASAP7_75t_R _36565__2061 (.H(net2061));
 TIEHIx1_ASAP7_75t_R _36566__2062 (.H(net2062));
 TIEHIx1_ASAP7_75t_R _36567__2063 (.H(net2063));
 TIEHIx1_ASAP7_75t_R _36568__2064 (.H(net2064));
 TIEHIx1_ASAP7_75t_R _36569__2065 (.H(net2065));
 TIEHIx1_ASAP7_75t_R _36570__2066 (.H(net2066));
 TIEHIx1_ASAP7_75t_R _36571__2067 (.H(net2067));
 TIEHIx1_ASAP7_75t_R _36572__2068 (.H(net2068));
 TIEHIx1_ASAP7_75t_R _36573__2069 (.H(net2069));
 TIEHIx1_ASAP7_75t_R _36574__2070 (.H(net2070));
 TIEHIx1_ASAP7_75t_R _36575__2071 (.H(net2071));
 TIEHIx1_ASAP7_75t_R _36576__2072 (.H(net2072));
 TIEHIx1_ASAP7_75t_R _36577__2073 (.H(net2073));
 TIEHIx1_ASAP7_75t_R _36578__2074 (.H(net2074));
 TIEHIx1_ASAP7_75t_R _36579__2075 (.H(net2075));
 TIEHIx1_ASAP7_75t_R _36580__2076 (.H(net2076));
 TIEHIx1_ASAP7_75t_R _36581__2077 (.H(net2077));
 TIEHIx1_ASAP7_75t_R _36582__2078 (.H(net2078));
 TIEHIx1_ASAP7_75t_R _36583__2079 (.H(net2079));
 TIEHIx1_ASAP7_75t_R _36584__2080 (.H(net2080));
 TIEHIx1_ASAP7_75t_R _36585__2081 (.H(net2081));
 TIEHIx1_ASAP7_75t_R _36586__2082 (.H(net2082));
 TIEHIx1_ASAP7_75t_R _36587__2083 (.H(net2083));
 TIEHIx1_ASAP7_75t_R _36588__2084 (.H(net2084));
 TIEHIx1_ASAP7_75t_R _36589__2085 (.H(net2085));
 TIEHIx1_ASAP7_75t_R _36590__2086 (.H(net2086));
 TIEHIx1_ASAP7_75t_R _36591__2087 (.H(net2087));
 TIEHIx1_ASAP7_75t_R _36592__2088 (.H(net2088));
 TIEHIx1_ASAP7_75t_R _36593__2089 (.H(net2089));
 TIEHIx1_ASAP7_75t_R _36594__2090 (.H(net2090));
 TIEHIx1_ASAP7_75t_R _36595__2091 (.H(net2091));
 TIEHIx1_ASAP7_75t_R _36596__2092 (.H(net2092));
 TIEHIx1_ASAP7_75t_R _36597__2093 (.H(net2093));
 TIEHIx1_ASAP7_75t_R _36598__2094 (.H(net2094));
 TIEHIx1_ASAP7_75t_R _36599__2095 (.H(net2095));
 TIEHIx1_ASAP7_75t_R _36600__2096 (.H(net2096));
 TIEHIx1_ASAP7_75t_R _36601__2097 (.H(net2097));
 TIEHIx1_ASAP7_75t_R _36602__2098 (.H(net2098));
 TIEHIx1_ASAP7_75t_R _36603__2099 (.H(net2099));
 TIEHIx1_ASAP7_75t_R _36604__2100 (.H(net2100));
 TIEHIx1_ASAP7_75t_R _36605__2101 (.H(net2101));
 TIEHIx1_ASAP7_75t_R _36606__2102 (.H(net2102));
 TIEHIx1_ASAP7_75t_R _36607__2103 (.H(net2103));
 TIEHIx1_ASAP7_75t_R _36608__2104 (.H(net2104));
 TIEHIx1_ASAP7_75t_R _36609__2105 (.H(net2105));
 TIEHIx1_ASAP7_75t_R _36610__2106 (.H(net2106));
 TIEHIx1_ASAP7_75t_R _36611__2107 (.H(net2107));
 TIEHIx1_ASAP7_75t_R _36612__2108 (.H(net2108));
 TIEHIx1_ASAP7_75t_R _36613__2109 (.H(net2109));
 TIEHIx1_ASAP7_75t_R _36614__2110 (.H(net2110));
 TIEHIx1_ASAP7_75t_R _36615__2111 (.H(net2111));
 TIEHIx1_ASAP7_75t_R _36616__2112 (.H(net2112));
 TIEHIx1_ASAP7_75t_R _36617__2113 (.H(net2113));
 TIEHIx1_ASAP7_75t_R _36619__2114 (.H(net2114));
 TIEHIx1_ASAP7_75t_R _36620__2115 (.H(net2115));
 TIEHIx1_ASAP7_75t_R _36621__2116 (.H(net2116));
 TIEHIx1_ASAP7_75t_R _36622__2117 (.H(net2117));
 TIEHIx1_ASAP7_75t_R _36623__2118 (.H(net2118));
 TIEHIx1_ASAP7_75t_R _36624__2119 (.H(net2119));
 TIEHIx1_ASAP7_75t_R _36658__2120 (.H(net2120));
 TIEHIx1_ASAP7_75t_R _36659__2121 (.H(net2121));
 TIEHIx1_ASAP7_75t_R _36660__2122 (.H(net2122));
 TIEHIx1_ASAP7_75t_R _36728__2123 (.H(net2123));
 TIEHIx1_ASAP7_75t_R _36761__2124 (.H(net2124));
 BUFx4_ASAP7_75t_R clkbuf_leaf_1_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_1_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_2_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_2_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_3_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_3_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_4_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_4_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_5_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_5_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_6_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_6_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_7_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_7_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_8_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_8_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_9_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_9_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_10_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_10_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_11_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_11_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_12_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_12_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_13_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_13_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_14_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_14_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_15_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_15_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_16_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_16_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_17_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_17_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_18_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_18_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_19_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_19_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_20_clk_i (.A(clknet_2_2__leaf_clk_i),
    .Y(clknet_leaf_20_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_21_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_21_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_22_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_22_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_23_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_23_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_24_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_24_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_25_clk_i (.A(clknet_2_3__leaf_clk_i),
    .Y(clknet_leaf_25_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_26_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_26_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_27_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_27_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_28_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_28_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_29_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_29_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_30_clk_i (.A(clknet_2_1__leaf_clk_i),
    .Y(clknet_leaf_30_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_31_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_31_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_32_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_32_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_leaf_33_clk_i (.A(clknet_2_0__leaf_clk_i),
    .Y(clknet_leaf_33_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_0_clk_i (.A(clk_i),
    .Y(clknet_0_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_0__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_0__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_1__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_1__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_2__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_2__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_2_3__f_clk_i (.A(clknet_0_clk_i),
    .Y(clknet_2_3__leaf_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_10_clk_i (.A(clknet_leaf_0_clk_i),
    .Y(clknet_level_0_1_10_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_11_clk_i (.A(clknet_level_0_1_10_clk_i),
    .Y(clknet_level_1_1_11_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_12_clk_i (.A(clknet_level_1_1_11_clk_i),
    .Y(clknet_level_2_1_12_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_13_clk_i (.A(clknet_level_2_1_12_clk_i),
    .Y(clknet_level_3_1_13_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_24_clk_i (.A(clknet_leaf_1_clk_i),
    .Y(clknet_level_0_1_24_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_25_clk_i (.A(clknet_level_0_1_24_clk_i),
    .Y(clknet_level_1_1_25_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_26_clk_i (.A(clknet_level_1_1_25_clk_i),
    .Y(clknet_level_2_1_26_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_27_clk_i (.A(clknet_level_2_1_26_clk_i),
    .Y(clknet_level_3_1_27_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_38_clk_i (.A(clknet_leaf_2_clk_i),
    .Y(clknet_level_0_1_38_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_39_clk_i (.A(clknet_level_0_1_38_clk_i),
    .Y(clknet_level_1_1_39_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_310_clk_i (.A(clknet_level_1_1_39_clk_i),
    .Y(clknet_level_2_1_310_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_311_clk_i (.A(clknet_level_2_1_310_clk_i),
    .Y(clknet_level_3_1_311_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_412_clk_i (.A(clknet_leaf_3_clk_i),
    .Y(clknet_level_0_1_412_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_413_clk_i (.A(clknet_level_0_1_412_clk_i),
    .Y(clknet_level_1_1_413_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_414_clk_i (.A(clknet_level_1_1_413_clk_i),
    .Y(clknet_level_2_1_414_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_415_clk_i (.A(clknet_level_2_1_414_clk_i),
    .Y(clknet_level_3_1_415_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_516_clk_i (.A(clknet_leaf_4_clk_i),
    .Y(clknet_level_0_1_516_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_517_clk_i (.A(clknet_level_0_1_516_clk_i),
    .Y(clknet_level_1_1_517_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_518_clk_i (.A(clknet_level_1_1_517_clk_i),
    .Y(clknet_level_2_1_518_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_519_clk_i (.A(clknet_level_2_1_518_clk_i),
    .Y(clknet_level_3_1_519_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_620_clk_i (.A(clknet_leaf_5_clk_i),
    .Y(clknet_level_0_1_620_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_621_clk_i (.A(clknet_level_0_1_620_clk_i),
    .Y(clknet_level_1_1_621_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_622_clk_i (.A(clknet_level_1_1_621_clk_i),
    .Y(clknet_level_2_1_622_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_623_clk_i (.A(clknet_level_2_1_622_clk_i),
    .Y(clknet_level_3_1_623_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_724_clk_i (.A(clknet_leaf_6_clk_i),
    .Y(clknet_level_0_1_724_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_725_clk_i (.A(clknet_level_0_1_724_clk_i),
    .Y(clknet_level_1_1_725_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_726_clk_i (.A(clknet_level_1_1_725_clk_i),
    .Y(clknet_level_2_1_726_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_727_clk_i (.A(clknet_level_2_1_726_clk_i),
    .Y(clknet_level_3_1_727_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_828_clk_i (.A(clknet_leaf_7_clk_i),
    .Y(clknet_level_0_1_828_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_829_clk_i (.A(clknet_level_0_1_828_clk_i),
    .Y(clknet_level_1_1_829_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_830_clk_i (.A(clknet_level_1_1_829_clk_i),
    .Y(clknet_level_2_1_830_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_831_clk_i (.A(clknet_level_2_1_830_clk_i),
    .Y(clknet_level_3_1_831_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_932_clk_i (.A(clknet_leaf_8_clk_i),
    .Y(clknet_level_0_1_932_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_933_clk_i (.A(clknet_level_0_1_932_clk_i),
    .Y(clknet_level_1_1_933_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_934_clk_i (.A(clknet_level_1_1_933_clk_i),
    .Y(clknet_level_2_1_934_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_935_clk_i (.A(clknet_level_2_1_934_clk_i),
    .Y(clknet_level_3_1_935_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1036_clk_i (.A(clknet_leaf_9_clk_i),
    .Y(clknet_level_0_1_1036_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1037_clk_i (.A(clknet_level_0_1_1036_clk_i),
    .Y(clknet_level_1_1_1037_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1038_clk_i (.A(clknet_level_1_1_1037_clk_i),
    .Y(clknet_level_2_1_1038_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1039_clk_i (.A(clknet_level_2_1_1038_clk_i),
    .Y(clknet_level_3_1_1039_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1140_clk_i (.A(clknet_leaf_10_clk_i),
    .Y(clknet_level_0_1_1140_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1141_clk_i (.A(clknet_level_0_1_1140_clk_i),
    .Y(clknet_level_1_1_1141_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1142_clk_i (.A(clknet_level_1_1_1141_clk_i),
    .Y(clknet_level_2_1_1142_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1143_clk_i (.A(clknet_level_2_1_1142_clk_i),
    .Y(clknet_level_3_1_1143_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1244_clk_i (.A(clknet_leaf_11_clk_i),
    .Y(clknet_level_0_1_1244_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1245_clk_i (.A(clknet_level_0_1_1244_clk_i),
    .Y(clknet_level_1_1_1245_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1246_clk_i (.A(clknet_level_1_1_1245_clk_i),
    .Y(clknet_level_2_1_1246_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1247_clk_i (.A(clknet_level_2_1_1246_clk_i),
    .Y(clknet_level_3_1_1247_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1348_clk_i (.A(clknet_leaf_12_clk_i),
    .Y(clknet_level_0_1_1348_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1349_clk_i (.A(clknet_level_0_1_1348_clk_i),
    .Y(clknet_level_1_1_1349_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1350_clk_i (.A(clknet_level_1_1_1349_clk_i),
    .Y(clknet_level_2_1_1350_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1351_clk_i (.A(clknet_level_2_1_1350_clk_i),
    .Y(clknet_level_3_1_1351_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1452_clk_i (.A(clknet_leaf_13_clk_i),
    .Y(clknet_level_0_1_1452_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1453_clk_i (.A(clknet_level_0_1_1452_clk_i),
    .Y(clknet_level_1_1_1453_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1454_clk_i (.A(clknet_level_1_1_1453_clk_i),
    .Y(clknet_level_2_1_1454_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1455_clk_i (.A(clknet_level_2_1_1454_clk_i),
    .Y(clknet_level_3_1_1455_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1556_clk_i (.A(clknet_leaf_14_clk_i),
    .Y(clknet_level_0_1_1556_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1557_clk_i (.A(clknet_level_0_1_1556_clk_i),
    .Y(clknet_level_1_1_1557_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1558_clk_i (.A(clknet_level_1_1_1557_clk_i),
    .Y(clknet_level_2_1_1558_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1559_clk_i (.A(clknet_level_2_1_1558_clk_i),
    .Y(clknet_level_3_1_1559_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1660_clk_i (.A(clknet_leaf_15_clk_i),
    .Y(clknet_level_0_1_1660_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1661_clk_i (.A(clknet_level_0_1_1660_clk_i),
    .Y(clknet_level_1_1_1661_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1662_clk_i (.A(clknet_level_1_1_1661_clk_i),
    .Y(clknet_level_2_1_1662_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1663_clk_i (.A(clknet_level_2_1_1662_clk_i),
    .Y(clknet_level_3_1_1663_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1764_clk_i (.A(clknet_leaf_16_clk_i),
    .Y(clknet_level_0_1_1764_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1765_clk_i (.A(clknet_level_0_1_1764_clk_i),
    .Y(clknet_level_1_1_1765_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1766_clk_i (.A(clknet_level_1_1_1765_clk_i),
    .Y(clknet_level_2_1_1766_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1767_clk_i (.A(clknet_level_2_1_1766_clk_i),
    .Y(clknet_level_3_1_1767_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1868_clk_i (.A(clknet_leaf_17_clk_i),
    .Y(clknet_level_0_1_1868_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1869_clk_i (.A(clknet_level_0_1_1868_clk_i),
    .Y(clknet_level_1_1_1869_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1870_clk_i (.A(clknet_level_1_1_1869_clk_i),
    .Y(clknet_level_2_1_1870_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1871_clk_i (.A(clknet_level_2_1_1870_clk_i),
    .Y(clknet_level_3_1_1871_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_1972_clk_i (.A(clknet_leaf_18_clk_i),
    .Y(clknet_level_0_1_1972_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_1973_clk_i (.A(clknet_level_0_1_1972_clk_i),
    .Y(clknet_level_1_1_1973_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_1974_clk_i (.A(clknet_level_1_1_1973_clk_i),
    .Y(clknet_level_2_1_1974_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_1975_clk_i (.A(clknet_level_2_1_1974_clk_i),
    .Y(clknet_level_3_1_1975_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2076_clk_i (.A(clknet_leaf_19_clk_i),
    .Y(clknet_level_0_1_2076_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2077_clk_i (.A(clknet_level_0_1_2076_clk_i),
    .Y(clknet_level_1_1_2077_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2078_clk_i (.A(clknet_level_1_1_2077_clk_i),
    .Y(clknet_level_2_1_2078_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2079_clk_i (.A(clknet_level_2_1_2078_clk_i),
    .Y(clknet_level_3_1_2079_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2180_clk_i (.A(clknet_leaf_20_clk_i),
    .Y(clknet_level_0_1_2180_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2181_clk_i (.A(clknet_level_0_1_2180_clk_i),
    .Y(clknet_level_1_1_2181_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2182_clk_i (.A(clknet_level_1_1_2181_clk_i),
    .Y(clknet_level_2_1_2182_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2183_clk_i (.A(clknet_level_2_1_2182_clk_i),
    .Y(clknet_level_3_1_2183_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2284_clk_i (.A(clknet_leaf_21_clk_i),
    .Y(clknet_level_0_1_2284_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2285_clk_i (.A(clknet_level_0_1_2284_clk_i),
    .Y(clknet_level_1_1_2285_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2286_clk_i (.A(clknet_level_1_1_2285_clk_i),
    .Y(clknet_level_2_1_2286_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2287_clk_i (.A(clknet_level_2_1_2286_clk_i),
    .Y(clknet_level_3_1_2287_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2388_clk_i (.A(clknet_leaf_22_clk_i),
    .Y(clknet_level_0_1_2388_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2389_clk_i (.A(clknet_level_0_1_2388_clk_i),
    .Y(clknet_level_1_1_2389_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2390_clk_i (.A(clknet_level_1_1_2389_clk_i),
    .Y(clknet_level_2_1_2390_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2391_clk_i (.A(clknet_level_2_1_2390_clk_i),
    .Y(clknet_level_3_1_2391_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2492_clk_i (.A(clknet_leaf_23_clk_i),
    .Y(clknet_level_0_1_2492_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2493_clk_i (.A(clknet_level_0_1_2492_clk_i),
    .Y(clknet_level_1_1_2493_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2494_clk_i (.A(clknet_level_1_1_2493_clk_i),
    .Y(clknet_level_2_1_2494_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2495_clk_i (.A(clknet_level_2_1_2494_clk_i),
    .Y(clknet_level_3_1_2495_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_2596_clk_i (.A(clknet_leaf_24_clk_i),
    .Y(clknet_level_0_1_2596_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_2597_clk_i (.A(clknet_level_0_1_2596_clk_i),
    .Y(clknet_level_1_1_2597_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_2598_clk_i (.A(clknet_level_1_1_2597_clk_i),
    .Y(clknet_level_2_1_2598_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_2599_clk_i (.A(clknet_level_2_1_2598_clk_i),
    .Y(clknet_level_3_1_2599_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_26100_clk_i (.A(clknet_leaf_25_clk_i),
    .Y(clknet_level_0_1_26100_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_26101_clk_i (.A(clknet_level_0_1_26100_clk_i),
    .Y(clknet_level_1_1_26101_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_26102_clk_i (.A(clknet_level_1_1_26101_clk_i),
    .Y(clknet_level_2_1_26102_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_26103_clk_i (.A(clknet_level_2_1_26102_clk_i),
    .Y(clknet_level_3_1_26103_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_27104_clk_i (.A(clknet_leaf_26_clk_i),
    .Y(clknet_level_0_1_27104_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_27105_clk_i (.A(clknet_level_0_1_27104_clk_i),
    .Y(clknet_level_1_1_27105_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_27106_clk_i (.A(clknet_level_1_1_27105_clk_i),
    .Y(clknet_level_2_1_27106_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_27107_clk_i (.A(clknet_level_2_1_27106_clk_i),
    .Y(clknet_level_3_1_27107_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_28108_clk_i (.A(clknet_leaf_27_clk_i),
    .Y(clknet_level_0_1_28108_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_28109_clk_i (.A(clknet_level_0_1_28108_clk_i),
    .Y(clknet_level_1_1_28109_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_28110_clk_i (.A(clknet_level_1_1_28109_clk_i),
    .Y(clknet_level_2_1_28110_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_28111_clk_i (.A(clknet_level_2_1_28110_clk_i),
    .Y(clknet_level_3_1_28111_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_29112_clk_i (.A(clknet_leaf_28_clk_i),
    .Y(clknet_level_0_1_29112_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_29113_clk_i (.A(clknet_level_0_1_29112_clk_i),
    .Y(clknet_level_1_1_29113_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_29114_clk_i (.A(clknet_level_1_1_29113_clk_i),
    .Y(clknet_level_2_1_29114_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_29115_clk_i (.A(clknet_level_2_1_29114_clk_i),
    .Y(clknet_level_3_1_29115_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_30116_clk_i (.A(clknet_leaf_29_clk_i),
    .Y(clknet_level_0_1_30116_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_30117_clk_i (.A(clknet_level_0_1_30116_clk_i),
    .Y(clknet_level_1_1_30117_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_30118_clk_i (.A(clknet_level_1_1_30117_clk_i),
    .Y(clknet_level_2_1_30118_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_30119_clk_i (.A(clknet_level_2_1_30118_clk_i),
    .Y(clknet_level_3_1_30119_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_31120_clk_i (.A(clknet_leaf_30_clk_i),
    .Y(clknet_level_0_1_31120_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_31121_clk_i (.A(clknet_level_0_1_31120_clk_i),
    .Y(clknet_level_1_1_31121_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_31122_clk_i (.A(clknet_level_1_1_31121_clk_i),
    .Y(clknet_level_2_1_31122_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_31123_clk_i (.A(clknet_level_2_1_31122_clk_i),
    .Y(clknet_level_3_1_31123_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_32124_clk_i (.A(clknet_leaf_31_clk_i),
    .Y(clknet_level_0_1_32124_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_32125_clk_i (.A(clknet_level_0_1_32124_clk_i),
    .Y(clknet_level_1_1_32125_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_32126_clk_i (.A(clknet_level_1_1_32125_clk_i),
    .Y(clknet_level_2_1_32126_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_32127_clk_i (.A(clknet_level_2_1_32126_clk_i),
    .Y(clknet_level_3_1_32127_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_33128_clk_i (.A(clknet_leaf_32_clk_i),
    .Y(clknet_level_0_1_33128_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_33129_clk_i (.A(clknet_level_0_1_33128_clk_i),
    .Y(clknet_level_1_1_33129_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_33130_clk_i (.A(clknet_level_1_1_33129_clk_i),
    .Y(clknet_level_2_1_33130_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_33131_clk_i (.A(clknet_level_2_1_33130_clk_i),
    .Y(clknet_level_3_1_33131_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_0_1_34132_clk_i (.A(clknet_leaf_33_clk_i),
    .Y(clknet_level_0_1_34132_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_1_1_34133_clk_i (.A(clknet_level_0_1_34132_clk_i),
    .Y(clknet_level_1_1_34133_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_2_1_34134_clk_i (.A(clknet_level_1_1_34133_clk_i),
    .Y(clknet_level_2_1_34134_clk_i));
 BUFx4_ASAP7_75t_R clkbuf_level_3_1_34135_clk_i (.A(clknet_level_2_1_34134_clk_i),
    .Y(clknet_level_3_1_34135_clk_i));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_0_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_0_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_1_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_1_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_2_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_2_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_3_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_3_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_4_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_4_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_5_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_5_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_6_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_6_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_7_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_7_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_8_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_8_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_9_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_9_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_10_core_clock_gate_i.clk_o  (.A(\clknet_2_2__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_10_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_11_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_11_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_12_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_12_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_13_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_13_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_14_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_14_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_15_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_15_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_16_core_clock_gate_i.clk_o  (.A(\clknet_2_3__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_16_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_17_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_17_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_18_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_18_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_19_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_19_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_20_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_20_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_21_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_21_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_22_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_22_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_23_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_23_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_24_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_24_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_25_core_clock_gate_i.clk_o  (.A(\clknet_2_1__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_25_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_26_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_26_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_27_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_27_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_28_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_28_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_29_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_29_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_30_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_30_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_leaf_31_core_clock_gate_i.clk_o  (.A(\clknet_2_0__leaf_core_clock_gate_i.clk_o ),
    .Y(\clknet_leaf_31_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_0_core_clock_gate_i.clk_o  (.A(\core_clock_gate_i.clk_o ),
    .Y(\clknet_0_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_0__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_0__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_1__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_1__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_2__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_2__leaf_core_clock_gate_i.clk_o ));
 BUFx4_ASAP7_75t_R \clkbuf_2_3__f_core_clock_gate_i.clk_o  (.A(\clknet_0_core_clock_gate_i.clk_o ),
    .Y(\clknet_2_3__leaf_core_clock_gate_i.clk_o ));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_00051_),
    .Y(net2125));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(net2125),
    .Y(net2126));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(_17267_),
    .Y(net2127));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net2127),
    .Y(net2128));
 BUFx2_ASAP7_75t_R rebuffer5 (.A(_17267_),
    .Y(net2129));
 BUFx2_ASAP7_75t_R rebuffer6 (.A(net2129),
    .Y(net2130));
 BUFx3_ASAP7_75t_R rebuffer7 (.A(_17397_),
    .Y(net2131));
 BUFx2_ASAP7_75t_R rebuffer8 (.A(net2131),
    .Y(net2132));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net2131),
    .Y(net2133));
 BUFx3_ASAP7_75t_R rebuffer10 (.A(_00052_),
    .Y(net2134));
 BUFx2_ASAP7_75t_R rebuffer11 (.A(net2134),
    .Y(net2135));
 BUFx2_ASAP7_75t_R rebuffer12 (.A(net170),
    .Y(net2136));
 BUFx2_ASAP7_75t_R rebuffer13 (.A(net2136),
    .Y(net2137));
 BUFx3_ASAP7_75t_R rebuffer14 (.A(net170),
    .Y(net2138));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(net2138),
    .Y(net2139));
 BUFx2_ASAP7_75t_R rebuffer16 (.A(net2138),
    .Y(net2140));
 BUFx2_ASAP7_75t_R rebuffer17 (.A(net170),
    .Y(net2141));
 BUFx2_ASAP7_75t_R rebuffer18 (.A(net2141),
    .Y(net2142));
 BUFx2_ASAP7_75t_R rebuffer19 (.A(net2297),
    .Y(net2143));
 BUFx2_ASAP7_75t_R rebuffer20 (.A(net2143),
    .Y(net2144));
 BUFx2_ASAP7_75t_R rebuffer21 (.A(_00015_),
    .Y(net2145));
 BUFx2_ASAP7_75t_R rebuffer22 (.A(net2145),
    .Y(net2146));
 BUFx2_ASAP7_75t_R rebuffer23 (.A(_17588_),
    .Y(net2147));
 BUFx2_ASAP7_75t_R rebuffer24 (.A(net2147),
    .Y(net2148));
 BUFx2_ASAP7_75t_R rebuffer25 (.A(net2148),
    .Y(net2149));
 BUFx2_ASAP7_75t_R rebuffer26 (.A(net2149),
    .Y(net2150));
 BUFx2_ASAP7_75t_R rebuffer27 (.A(_17531_),
    .Y(net2151));
 BUFx3_ASAP7_75t_R rebuffer28 (.A(net168),
    .Y(net2152));
 BUFx2_ASAP7_75t_R rebuffer29 (.A(net2152),
    .Y(net2153));
 BUFx2_ASAP7_75t_R rebuffer30 (.A(net2153),
    .Y(net2154));
 BUFx3_ASAP7_75t_R rebuffer31 (.A(net2153),
    .Y(net2155));
 BUFx2_ASAP7_75t_R rebuffer32 (.A(net2155),
    .Y(net2156));
 BUFx2_ASAP7_75t_R rebuffer33 (.A(net168),
    .Y(net2157));
 BUFx2_ASAP7_75t_R rebuffer34 (.A(net2157),
    .Y(net2158));
 BUFx2_ASAP7_75t_R rebuffer35 (.A(_02352_),
    .Y(net2159));
 BUFx6f_ASAP7_75t_R rebuffer36 (.A(_02352_),
    .Y(net2160));
 BUFx2_ASAP7_75t_R rebuffer37 (.A(_17274_),
    .Y(net2161));
 BUFx2_ASAP7_75t_R rebuffer38 (.A(net2161),
    .Y(net2162));
 BUFx3_ASAP7_75t_R rebuffer39 (.A(_00038_),
    .Y(net2163));
 BUFx2_ASAP7_75t_R rebuffer40 (.A(net2163),
    .Y(net2164));
 BUFx2_ASAP7_75t_R rebuffer41 (.A(net2164),
    .Y(net2165));
 BUFx2_ASAP7_75t_R rebuffer42 (.A(_17076_),
    .Y(net2166));
 BUFx2_ASAP7_75t_R rebuffer43 (.A(_17077_),
    .Y(net2167));
 BUFx2_ASAP7_75t_R rebuffer44 (.A(_16991_),
    .Y(net2168));
 BUFx2_ASAP7_75t_R rebuffer45 (.A(_16923_),
    .Y(net2169));
 BUFx2_ASAP7_75t_R rebuffer46 (.A(net2251),
    .Y(net2170));
 BUFx3_ASAP7_75t_R rebuffer47 (.A(net166),
    .Y(net2171));
 BUFx2_ASAP7_75t_R rebuffer48 (.A(net2171),
    .Y(net2172));
 BUFx2_ASAP7_75t_R rebuffer49 (.A(net2171),
    .Y(net2173));
 BUFx2_ASAP7_75t_R rebuffer50 (.A(net2173),
    .Y(net2174));
 BUFx3_ASAP7_75t_R rebuffer51 (.A(net2173),
    .Y(net2175));
 BUFx2_ASAP7_75t_R rebuffer52 (.A(net2175),
    .Y(net2176));
 BUFx2_ASAP7_75t_R rebuffer53 (.A(net164),
    .Y(net2177));
 BUFx2_ASAP7_75t_R rebuffer54 (.A(net2177),
    .Y(net2178));
 BUFx3_ASAP7_75t_R rebuffer55 (.A(net164),
    .Y(net2179));
 BUFx2_ASAP7_75t_R rebuffer56 (.A(net2179),
    .Y(net2180));
 BUFx2_ASAP7_75t_R rebuffer57 (.A(_16568_),
    .Y(net2181));
 BUFx2_ASAP7_75t_R rebuffer58 (.A(net2181),
    .Y(net2182));
 BUFx2_ASAP7_75t_R rebuffer59 (.A(net2182),
    .Y(net2183));
 BUFx2_ASAP7_75t_R rebuffer60 (.A(net2182),
    .Y(net2184));
 BUFx6f_ASAP7_75t_R rebuffer61 (.A(_05964_),
    .Y(net2185));
 BUFx3_ASAP7_75t_R rebuffer62 (.A(net2185),
    .Y(net2186));
 BUFx2_ASAP7_75t_R rebuffer63 (.A(net2185),
    .Y(net2187));
 BUFx2_ASAP7_75t_R rebuffer64 (.A(net2185),
    .Y(net2188));
 BUFx2_ASAP7_75t_R rebuffer65 (.A(net2185),
    .Y(net2189));
 BUFx12f_ASAP7_75t_R rebuffer66 (.A(_05883_),
    .Y(net2190));
 BUFx2_ASAP7_75t_R rebuffer67 (.A(net2190),
    .Y(net2191));
 BUFx2_ASAP7_75t_R rebuffer68 (.A(net2190),
    .Y(net2192));
 BUFx2_ASAP7_75t_R rebuffer69 (.A(_17558_),
    .Y(net2193));
 BUFx2_ASAP7_75t_R rebuffer70 (.A(_17558_),
    .Y(net2194));
 BUFx2_ASAP7_75t_R rebuffer71 (.A(net2194),
    .Y(net2195));
 BUFx2_ASAP7_75t_R rebuffer72 (.A(_00031_),
    .Y(net2196));
 BUFx12_ASAP7_75t_R split73 (.A(_08621_),
    .Y(net2197));
 BUFx6f_ASAP7_75t_R rebuffer74 (.A(_08621_),
    .Y(net2198));
 BUFx2_ASAP7_75t_R rebuffer75 (.A(net180),
    .Y(net2199));
 BUFx2_ASAP7_75t_R rebuffer76 (.A(net2199),
    .Y(net2200));
 BUFx2_ASAP7_75t_R rebuffer77 (.A(net2199),
    .Y(net2201));
 BUFx3_ASAP7_75t_R rebuffer78 (.A(net2201),
    .Y(net2202));
 BUFx2_ASAP7_75t_R rebuffer79 (.A(net2201),
    .Y(net2203));
 BUFx2_ASAP7_75t_R rebuffer80 (.A(net180),
    .Y(net2204));
 BUFx2_ASAP7_75t_R rebuffer81 (.A(net2204),
    .Y(net2205));
 BUFx2_ASAP7_75t_R rebuffer82 (.A(_05849_),
    .Y(net2206));
 BUFx3_ASAP7_75t_R rebuffer83 (.A(net2206),
    .Y(net2207));
 BUFx2_ASAP7_75t_R rebuffer84 (.A(net2207),
    .Y(net2208));
 BUFx2_ASAP7_75t_R rebuffer85 (.A(_00289_),
    .Y(net2209));
 BUFx6f_ASAP7_75t_R rebuffer86 (.A(_00289_),
    .Y(net2210));
 BUFx2_ASAP7_75t_R rebuffer87 (.A(net2210),
    .Y(net2211));
 BUFx2_ASAP7_75t_R rebuffer88 (.A(net2378),
    .Y(net2212));
 BUFx2_ASAP7_75t_R rebuffer89 (.A(net2212),
    .Y(net2213));
 BUFx2_ASAP7_75t_R rebuffer90 (.A(net2378),
    .Y(net2214));
 BUFx2_ASAP7_75t_R rebuffer91 (.A(net2244),
    .Y(net2215));
 BUFx2_ASAP7_75t_R rebuffer92 (.A(net2244),
    .Y(net2216));
 BUFx2_ASAP7_75t_R rebuffer93 (.A(net2227),
    .Y(net2217));
 BUFx2_ASAP7_75t_R rebuffer94 (.A(_14290_),
    .Y(net2218));
 BUFx2_ASAP7_75t_R rebuffer95 (.A(net2218),
    .Y(net2219));
 BUFx2_ASAP7_75t_R rebuffer96 (.A(net2218),
    .Y(net2220));
 BUFx2_ASAP7_75t_R rebuffer97 (.A(net2218),
    .Y(net2221));
 BUFx2_ASAP7_75t_R rebuffer98 (.A(_14126_),
    .Y(net2222));
 BUFx3_ASAP7_75t_R rebuffer99 (.A(_05833_),
    .Y(net2223));
 BUFx2_ASAP7_75t_R rebuffer100 (.A(net2223),
    .Y(net2224));
 BUFx2_ASAP7_75t_R rebuffer101 (.A(net2223),
    .Y(net2225));
 BUFx2_ASAP7_75t_R rebuffer102 (.A(net2223),
    .Y(net2226));
 BUFx12f_ASAP7_75t_R rebuffer103 (.A(_13391_),
    .Y(net2227));
 BUFx2_ASAP7_75t_R rebuffer104 (.A(net2227),
    .Y(net2228));
 BUFx2_ASAP7_75t_R rebuffer105 (.A(net2227),
    .Y(net2229));
 BUFx2_ASAP7_75t_R rebuffer106 (.A(_14233_),
    .Y(net2230));
 BUFx2_ASAP7_75t_R rebuffer107 (.A(_14233_),
    .Y(net2231));
 BUFx2_ASAP7_75t_R rebuffer108 (.A(_18031_),
    .Y(net2232));
 BUFx2_ASAP7_75t_R rebuffer109 (.A(net2232),
    .Y(net2233));
 BUFx2_ASAP7_75t_R rebuffer110 (.A(_05852_),
    .Y(net2234));
 BUFx2_ASAP7_75t_R rebuffer111 (.A(net2234),
    .Y(net2235));
 BUFx2_ASAP7_75t_R rebuffer112 (.A(_00024_),
    .Y(net2236));
 BUFx2_ASAP7_75t_R rebuffer113 (.A(net2236),
    .Y(net2237));
 BUFx2_ASAP7_75t_R rebuffer114 (.A(_17617_),
    .Y(net2238));
 BUFx2_ASAP7_75t_R rebuffer115 (.A(net2238),
    .Y(net2239));
 BUFx2_ASAP7_75t_R rebuffer116 (.A(net2238),
    .Y(net2240));
 BUFx2_ASAP7_75t_R rebuffer117 (.A(_17617_),
    .Y(net2241));
 BUFx4f_ASAP7_75t_R split118 (.A(_13391_),
    .Y(net2242));
 BUFx3_ASAP7_75t_R split119 (.A(_05964_),
    .Y(net2243));
 BUFx12f_ASAP7_75t_R rebuffer120 (.A(_13391_),
    .Y(net2244));
 BUFx4f_ASAP7_75t_R rebuffer121 (.A(_05821_),
    .Y(net2245));
 BUFx2_ASAP7_75t_R rebuffer122 (.A(net2245),
    .Y(net2246));
 BUFx2_ASAP7_75t_R rebuffer123 (.A(net2245),
    .Y(net2247));
 BUFx10_ASAP7_75t_R split124 (.A(net367),
    .Y(net2248));
 BUFx4f_ASAP7_75t_R split125 (.A(net367),
    .Y(net2249));
 BUFx3_ASAP7_75t_R rebuffer126 (.A(_17313_),
    .Y(net2250));
 BUFx2_ASAP7_75t_R split127 (.A(_16924_),
    .Y(net2251));
 BUFx2_ASAP7_75t_R rebuffer128 (.A(_05962_),
    .Y(net2252));
 BUFx2_ASAP7_75t_R split129 (.A(_05849_),
    .Y(net2253));
 BUFx2_ASAP7_75t_R rebuffer130 (.A(net158),
    .Y(net2254));
 BUFx2_ASAP7_75t_R rebuffer131 (.A(net2254),
    .Y(net2255));
 BUFx2_ASAP7_75t_R rebuffer132 (.A(net2255),
    .Y(net2256));
 BUFx12_ASAP7_75t_R split133 (.A(net2265),
    .Y(net2257));
 BUFx10_ASAP7_75t_R split134 (.A(net360),
    .Y(net2258));
 BUFx4f_ASAP7_75t_R split135 (.A(net364),
    .Y(net2259));
 BUFx12f_ASAP7_75t_R split136 (.A(_13359_),
    .Y(net2260));
 BUFx2_ASAP7_75t_R rebuffer137 (.A(_00290_),
    .Y(net2261));
 BUFx2_ASAP7_75t_R rebuffer138 (.A(net2261),
    .Y(net2262));
 BUFx2_ASAP7_75t_R rebuffer139 (.A(net2262),
    .Y(net2263));
 BUFx2_ASAP7_75t_R rebuffer140 (.A(_00290_),
    .Y(net2264));
 BUFx3_ASAP7_75t_R split141 (.A(net364),
    .Y(net2265));
 BUFx2_ASAP7_75t_R rebuffer142 (.A(net360),
    .Y(net2266));
 BUFx3_ASAP7_75t_R rebuffer143 (.A(net2266),
    .Y(net2267));
 BUFx2_ASAP7_75t_R rebuffer144 (.A(net2267),
    .Y(net2268));
 BUFx6f_ASAP7_75t_R split145 (.A(net2276),
    .Y(net2269));
 BUFx2_ASAP7_75t_R rebuffer146 (.A(_05912_),
    .Y(net2270));
 BUFx3_ASAP7_75t_R rebuffer147 (.A(net2270),
    .Y(net2271));
 BUFx2_ASAP7_75t_R rebuffer148 (.A(net2271),
    .Y(net2272));
 BUFx3_ASAP7_75t_R rebuffer149 (.A(net2272),
    .Y(net2273));
 BUFx2_ASAP7_75t_R rebuffer150 (.A(net2273),
    .Y(net2274));
 BUFx2_ASAP7_75t_R rebuffer151 (.A(_05912_),
    .Y(net2275));
 BUFx4f_ASAP7_75t_R split152 (.A(net365),
    .Y(net2276));
 BUFx6f_ASAP7_75t_R split153 (.A(net2336),
    .Y(net2277));
 BUFx16f_ASAP7_75t_R split154 (.A(net326),
    .Y(net2278));
 BUFx12f_ASAP7_75t_R split155 (.A(net353),
    .Y(net2279));
 BUFx6f_ASAP7_75t_R split156 (.A(net358),
    .Y(net2280));
 BUFx2_ASAP7_75t_R rebuffer157 (.A(net2375),
    .Y(net2281));
 BUFx2_ASAP7_75t_R rebuffer158 (.A(net2375),
    .Y(net2282));
 BUFx2_ASAP7_75t_R rebuffer159 (.A(net2375),
    .Y(net2283));
 BUFx12f_ASAP7_75t_R split160 (.A(net2294),
    .Y(net2284));
 BUFx4f_ASAP7_75t_R rebuffer161 (.A(_05863_),
    .Y(net2285));
 BUFx2_ASAP7_75t_R rebuffer162 (.A(net2285),
    .Y(net2286));
 BUFx2_ASAP7_75t_R rebuffer163 (.A(net2286),
    .Y(net2287));
 BUFx2_ASAP7_75t_R rebuffer164 (.A(net358),
    .Y(net2288));
 BUFx2_ASAP7_75t_R rebuffer165 (.A(_14008_),
    .Y(net2289));
 BUFx12f_ASAP7_75t_R rebuffer166 (.A(_14008_),
    .Y(net2290));
 BUFx2_ASAP7_75t_R rebuffer167 (.A(net2290),
    .Y(net2291));
 BUFx2_ASAP7_75t_R rebuffer168 (.A(_14008_),
    .Y(net2292));
 BUFx2_ASAP7_75t_R rebuffer169 (.A(net2292),
    .Y(net2293));
 BUFx12f_ASAP7_75t_R split170 (.A(net354),
    .Y(net2294));
 BUFx2_ASAP7_75t_R rebuffer171 (.A(_05837_),
    .Y(net2295));
 BUFx2_ASAP7_75t_R rebuffer172 (.A(net2295),
    .Y(net2296));
 BUFx6f_ASAP7_75t_R rebuffer173 (.A(_01745_),
    .Y(net2297));
 BUFx2_ASAP7_75t_R rebuffer174 (.A(net2297),
    .Y(net2298));
 BUFx2_ASAP7_75t_R rebuffer175 (.A(net2297),
    .Y(net2299));
 BUFx2_ASAP7_75t_R rebuffer176 (.A(_00288_),
    .Y(net2300));
 BUFx6f_ASAP7_75t_R rebuffer177 (.A(net2300),
    .Y(net2301));
 BUFx2_ASAP7_75t_R rebuffer178 (.A(net2301),
    .Y(net2302));
 BUFx2_ASAP7_75t_R rebuffer179 (.A(net2302),
    .Y(net2303));
 BUFx2_ASAP7_75t_R rebuffer180 (.A(net2301),
    .Y(net2304));
 BUFx2_ASAP7_75t_R rebuffer181 (.A(_05938_),
    .Y(net2305));
 BUFx2_ASAP7_75t_R rebuffer182 (.A(net2305),
    .Y(net2306));
 BUFx2_ASAP7_75t_R rebuffer183 (.A(_05938_),
    .Y(net2307));
 BUFx2_ASAP7_75t_R rebuffer184 (.A(_05938_),
    .Y(net2308));
 BUFx2_ASAP7_75t_R rebuffer185 (.A(net2308),
    .Y(net2309));
 BUFx2_ASAP7_75t_R rebuffer186 (.A(_15396_),
    .Y(net2310));
 BUFx2_ASAP7_75t_R rebuffer187 (.A(net2310),
    .Y(net2311));
 BUFx2_ASAP7_75t_R rebuffer188 (.A(net2310),
    .Y(net2312));
 BUFx2_ASAP7_75t_R rebuffer189 (.A(_00246_),
    .Y(net2313));
 BUFx3_ASAP7_75t_R rebuffer190 (.A(net2313),
    .Y(net2314));
 BUFx3_ASAP7_75t_R rebuffer191 (.A(net2313),
    .Y(net2315));
 BUFx2_ASAP7_75t_R rebuffer192 (.A(_05887_),
    .Y(net2316));
 BUFx4f_ASAP7_75t_R rebuffer193 (.A(net2316),
    .Y(net2317));
 BUFx3_ASAP7_75t_R rebuffer194 (.A(net2316),
    .Y(net2318));
 BUFx2_ASAP7_75t_R rebuffer195 (.A(net2318),
    .Y(net2319));
 BUFx2_ASAP7_75t_R rebuffer196 (.A(net2318),
    .Y(net2320));
 BUFx2_ASAP7_75t_R rebuffer197 (.A(net354),
    .Y(net2321));
 BUFx2_ASAP7_75t_R rebuffer198 (.A(_15050_),
    .Y(net2322));
 BUFx2_ASAP7_75t_R rebuffer199 (.A(net2322),
    .Y(net2323));
 BUFx2_ASAP7_75t_R rebuffer200 (.A(_05904_),
    .Y(net2324));
 BUFx2_ASAP7_75t_R rebuffer201 (.A(net2324),
    .Y(net2325));
 BUFx2_ASAP7_75t_R rebuffer202 (.A(net2324),
    .Y(net2326));
 BUFx2_ASAP7_75t_R rebuffer203 (.A(net2326),
    .Y(net2327));
 BUFx2_ASAP7_75t_R rebuffer204 (.A(_05904_),
    .Y(net2328));
 BUFx12f_ASAP7_75t_R split205 (.A(net2198),
    .Y(net2329));
 BUFx6f_ASAP7_75t_R split206 (.A(net2198),
    .Y(net2330));
 BUFx4f_ASAP7_75t_R split207 (.A(net355),
    .Y(net2331));
 BUFx3_ASAP7_75t_R split208 (.A(net359),
    .Y(net2332));
 BUFx6f_ASAP7_75t_R split209 (.A(net363),
    .Y(net2333));
 BUFx3_ASAP7_75t_R rebuffer210 (.A(_01410_),
    .Y(net2334));
 BUFx2_ASAP7_75t_R rebuffer211 (.A(net2334),
    .Y(net2335));
 BUFx2_ASAP7_75t_R split212 (.A(net366),
    .Y(net2336));
 BUFx6f_ASAP7_75t_R rebuffer213 (.A(_05845_),
    .Y(net2337));
 BUFx6f_ASAP7_75t_R rebuffer214 (.A(net2337),
    .Y(net2338));
 BUFx2_ASAP7_75t_R rebuffer215 (.A(net2338),
    .Y(net2339));
 BUFx2_ASAP7_75t_R rebuffer216 (.A(net2339),
    .Y(net2340));
 BUFx2_ASAP7_75t_R rebuffer217 (.A(net2337),
    .Y(net2341));
 BUFx2_ASAP7_75t_R rebuffer218 (.A(net355),
    .Y(net2342));
 BUFx6f_ASAP7_75t_R rebuffer219 (.A(net2342),
    .Y(net2343));
 BUFx2_ASAP7_75t_R rebuffer220 (.A(net2342),
    .Y(net2344));
 BUFx4f_ASAP7_75t_R rebuffer221 (.A(_05855_),
    .Y(net2345));
 BUFx2_ASAP7_75t_R rebuffer222 (.A(net2345),
    .Y(net2346));
 BUFx2_ASAP7_75t_R rebuffer223 (.A(net2345),
    .Y(net2347));
 BUFx2_ASAP7_75t_R rebuffer224 (.A(net2345),
    .Y(net2348));
 BUFx2_ASAP7_75t_R rebuffer225 (.A(_05870_),
    .Y(net2349));
 BUFx2_ASAP7_75t_R rebuffer226 (.A(net2349),
    .Y(net2350));
 BUFx2_ASAP7_75t_R rebuffer227 (.A(net2350),
    .Y(net2351));
 BUFx6f_ASAP7_75t_R split228 (.A(net406),
    .Y(net2352));
 BUFx3_ASAP7_75t_R rebuffer229 (.A(_05879_),
    .Y(net2353));
 BUFx2_ASAP7_75t_R rebuffer230 (.A(net2353),
    .Y(net2354));
 BUFx2_ASAP7_75t_R rebuffer231 (.A(net2353),
    .Y(net2355));
 BUFx2_ASAP7_75t_R rebuffer232 (.A(net2355),
    .Y(net2356));
 BUFx3_ASAP7_75t_R split233 (.A(net365),
    .Y(net2357));
 BUFx2_ASAP7_75t_R rebuffer234 (.A(_01744_),
    .Y(net2358));
 BUFx2_ASAP7_75t_R rebuffer235 (.A(net2358),
    .Y(net2359));
 BUFx2_ASAP7_75t_R rebuffer236 (.A(net2358),
    .Y(net2360));
 BUFx2_ASAP7_75t_R rebuffer237 (.A(net2358),
    .Y(net2361));
 BUFx2_ASAP7_75t_R rebuffer238 (.A(net2361),
    .Y(net2362));
 BUFx2_ASAP7_75t_R rebuffer239 (.A(net2361),
    .Y(net2363));
 BUFx2_ASAP7_75t_R rebuffer240 (.A(_05894_),
    .Y(net2364));
 BUFx6f_ASAP7_75t_R rebuffer241 (.A(net2364),
    .Y(net2365));
 BUFx2_ASAP7_75t_R rebuffer242 (.A(net2365),
    .Y(net2366));
 BUFx2_ASAP7_75t_R rebuffer243 (.A(net2366),
    .Y(net2367));
 BUFx2_ASAP7_75t_R rebuffer244 (.A(net2365),
    .Y(net2368));
 BUFx4f_ASAP7_75t_R rebuffer245 (.A(net406),
    .Y(net2369));
 BUFx3_ASAP7_75t_R split246 (.A(_05837_),
    .Y(net2370));
 BUFx4f_ASAP7_75t_R split247 (.A(net2284),
    .Y(net2371));
 BUFx2_ASAP7_75t_R rebuffer248 (.A(net2279),
    .Y(net2372));
 BUFx12f_ASAP7_75t_R split249 (.A(net353),
    .Y(net2373));
 BUFx2_ASAP7_75t_R rebuffer250 (.A(net363),
    .Y(net2374));
 BUFx12f_ASAP7_75t_R rebuffer251 (.A(net353),
    .Y(net2375));
 BUFx6f_ASAP7_75t_R split252 (.A(net402),
    .Y(net2376));
 BUFx4f_ASAP7_75t_R split253 (.A(net406),
    .Y(net2377));
 BUFx3_ASAP7_75t_R split254 (.A(net2210),
    .Y(net2378));
 BUFx10_ASAP7_75t_R split255 (.A(net411),
    .Y(net2379));
 BUFx2_ASAP7_75t_R hold256 (.A(net2387),
    .Y(net2380));
 BUFx2_ASAP7_75t_R hold257 (.A(net2384),
    .Y(net2381));
 BUFx2_ASAP7_75t_R hold258 (.A(net2386),
    .Y(net2382));
 BUFx2_ASAP7_75t_R hold259 (.A(net2388),
    .Y(net2383));
 BUFx2_ASAP7_75t_R hold260 (.A(net2390),
    .Y(net2384));
 BUFx2_ASAP7_75t_R hold261 (.A(net2381),
    .Y(net2385));
 BUFx2_ASAP7_75t_R hold262 (.A(rst_ni),
    .Y(net2386));
 BUFx2_ASAP7_75t_R hold263 (.A(net2382),
    .Y(net2387));
 BUFx2_ASAP7_75t_R hold264 (.A(net2380),
    .Y(net2388));
 BUFx2_ASAP7_75t_R hold265 (.A(net2383),
    .Y(net2389));
 BUFx2_ASAP7_75t_R hold266 (.A(net148),
    .Y(net2390));
 BUFx2_ASAP7_75t_R hold267 (.A(net3938),
    .Y(net2391));
 BUFx2_ASAP7_75t_R hold268 (.A(net3942),
    .Y(net2392));
 BUFx2_ASAP7_75t_R hold269 (.A(_04362_),
    .Y(net2393));
 BUFx2_ASAP7_75t_R hold270 (.A(net3968),
    .Y(net2394));
 BUFx2_ASAP7_75t_R hold271 (.A(net3972),
    .Y(net2395));
 BUFx2_ASAP7_75t_R hold272 (.A(net3800),
    .Y(net2396));
 BUFx2_ASAP7_75t_R hold273 (.A(net3905),
    .Y(net2397));
 BUFx2_ASAP7_75t_R hold274 (.A(net3909),
    .Y(net2398));
 BUFx2_ASAP7_75t_R hold275 (.A(net3911),
    .Y(net2399));
 BUFx2_ASAP7_75t_R hold276 (.A(net2762),
    .Y(net2400));
 BUFx2_ASAP7_75t_R hold277 (.A(net2766),
    .Y(net2401));
 BUFx2_ASAP7_75t_R hold278 (.A(_04452_),
    .Y(net2402));
 BUFx2_ASAP7_75t_R hold279 (.A(net2775),
    .Y(net2403));
 BUFx2_ASAP7_75t_R hold280 (.A(net2779),
    .Y(net2404));
 BUFx2_ASAP7_75t_R hold281 (.A(_04465_),
    .Y(net2405));
 BUFx2_ASAP7_75t_R hold282 (.A(net2783),
    .Y(net2406));
 BUFx2_ASAP7_75t_R hold283 (.A(net2787),
    .Y(net2407));
 BUFx2_ASAP7_75t_R hold284 (.A(_04449_),
    .Y(net2408));
 BUFx2_ASAP7_75t_R hold285 (.A(net2808),
    .Y(net2409));
 BUFx2_ASAP7_75t_R hold286 (.A(net2812),
    .Y(net2410));
 BUFx2_ASAP7_75t_R hold287 (.A(_04467_),
    .Y(net2411));
 BUFx2_ASAP7_75t_R hold288 (.A(net3974),
    .Y(net2412));
 BUFx2_ASAP7_75t_R hold289 (.A(net3978),
    .Y(net2413));
 BUFx2_ASAP7_75t_R hold290 (.A(net3806),
    .Y(net2414));
 BUFx2_ASAP7_75t_R hold291 (.A(net3980),
    .Y(net2415));
 BUFx2_ASAP7_75t_R hold292 (.A(net3984),
    .Y(net2416));
 BUFx2_ASAP7_75t_R hold293 (.A(net3818),
    .Y(net2417));
 BUFx2_ASAP7_75t_R hold294 (.A(net3986),
    .Y(net2418));
 BUFx2_ASAP7_75t_R hold295 (.A(net3810),
    .Y(net2419));
 BUFx2_ASAP7_75t_R hold296 (.A(net3812),
    .Y(net2420));
 BUFx2_ASAP7_75t_R hold297 (.A(net3991),
    .Y(net2421));
 BUFx2_ASAP7_75t_R hold298 (.A(net3822),
    .Y(net2422));
 BUFx2_ASAP7_75t_R hold299 (.A(net3824),
    .Y(net2423));
 BUFx2_ASAP7_75t_R hold300 (.A(net2840),
    .Y(net2424));
 BUFx2_ASAP7_75t_R hold301 (.A(net2844),
    .Y(net2425));
 BUFx2_ASAP7_75t_R hold302 (.A(_04439_),
    .Y(net2426));
 BUFx2_ASAP7_75t_R hold303 (.A(net2824),
    .Y(net2427));
 BUFx2_ASAP7_75t_R hold304 (.A(net2828),
    .Y(net2428));
 BUFx2_ASAP7_75t_R hold305 (.A(_04451_),
    .Y(net2429));
 BUFx2_ASAP7_75t_R hold306 (.A(net2832),
    .Y(net2430));
 BUFx2_ASAP7_75t_R hold307 (.A(net2836),
    .Y(net2431));
 BUFx2_ASAP7_75t_R hold308 (.A(_04448_),
    .Y(net2432));
 BUFx2_ASAP7_75t_R hold309 (.A(net3914),
    .Y(net2433));
 BUFx2_ASAP7_75t_R hold310 (.A(net3918),
    .Y(net2434));
 BUFx2_ASAP7_75t_R hold311 (.A(net3920),
    .Y(net2435));
 BUFx2_ASAP7_75t_R hold312 (.A(net3996),
    .Y(net2436));
 BUFx2_ASAP7_75t_R hold313 (.A(net3834),
    .Y(net2437));
 BUFx2_ASAP7_75t_R hold314 (.A(net3836),
    .Y(net2438));
 BUFx2_ASAP7_75t_R hold315 (.A(net4006),
    .Y(net2439));
 BUFx2_ASAP7_75t_R hold316 (.A(net3828),
    .Y(net2440));
 BUFx2_ASAP7_75t_R hold317 (.A(net3830),
    .Y(net2441));
 BUFx2_ASAP7_75t_R hold318 (.A(net2856),
    .Y(net2442));
 BUFx2_ASAP7_75t_R hold319 (.A(net2860),
    .Y(net2443));
 BUFx2_ASAP7_75t_R hold320 (.A(_04468_),
    .Y(net2444));
 BUFx2_ASAP7_75t_R hold321 (.A(net2872),
    .Y(net2445));
 BUFx2_ASAP7_75t_R hold322 (.A(net2876),
    .Y(net2446));
 BUFx2_ASAP7_75t_R hold323 (.A(_04458_),
    .Y(net2447));
 BUFx2_ASAP7_75t_R hold324 (.A(net2791),
    .Y(net2448));
 BUFx2_ASAP7_75t_R hold325 (.A(net2795),
    .Y(net2449));
 BUFx2_ASAP7_75t_R hold326 (.A(_04446_),
    .Y(net2450));
 BUFx2_ASAP7_75t_R hold327 (.A(net2880),
    .Y(net2451));
 BUFx2_ASAP7_75t_R hold328 (.A(net2884),
    .Y(net2452));
 BUFx2_ASAP7_75t_R hold329 (.A(_04442_),
    .Y(net2453));
 BUFx2_ASAP7_75t_R hold330 (.A(net2848),
    .Y(net2454));
 BUFx2_ASAP7_75t_R hold331 (.A(net2852),
    .Y(net2455));
 BUFx2_ASAP7_75t_R hold332 (.A(_04464_),
    .Y(net2456));
 BUFx2_ASAP7_75t_R hold333 (.A(net4001),
    .Y(net2457));
 BUFx2_ASAP7_75t_R hold334 (.A(net3840),
    .Y(net2458));
 BUFx2_ASAP7_75t_R hold335 (.A(net3842),
    .Y(net2459));
 BUFx2_ASAP7_75t_R hold336 (.A(net3292),
    .Y(net2460));
 BUFx2_ASAP7_75t_R hold337 (.A(net3296),
    .Y(net2461));
 BUFx2_ASAP7_75t_R hold338 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .Y(net2462));
 BUFx2_ASAP7_75t_R hold339 (.A(net2888),
    .Y(net2463));
 BUFx2_ASAP7_75t_R hold340 (.A(net2892),
    .Y(net2464));
 BUFx2_ASAP7_75t_R hold341 (.A(_04455_),
    .Y(net2465));
 BUFx2_ASAP7_75t_R hold342 (.A(net3071),
    .Y(net2466));
 BUFx2_ASAP7_75t_R hold343 (.A(net3075),
    .Y(net2467));
 BUFx2_ASAP7_75t_R hold344 (.A(_04443_),
    .Y(net2468));
 BUFx2_ASAP7_75t_R hold345 (.A(net2864),
    .Y(net2469));
 BUFx2_ASAP7_75t_R hold346 (.A(net2868),
    .Y(net2470));
 BUFx2_ASAP7_75t_R hold347 (.A(_04444_),
    .Y(net2471));
 BUFx2_ASAP7_75t_R hold348 (.A(net2896),
    .Y(net2472));
 BUFx2_ASAP7_75t_R hold349 (.A(net2900),
    .Y(net2473));
 BUFx2_ASAP7_75t_R hold350 (.A(_04454_),
    .Y(net2474));
 BUFx2_ASAP7_75t_R hold351 (.A(net3954),
    .Y(net2475));
 BUFx2_ASAP7_75t_R hold352 (.A(net3958),
    .Y(net2476));
 BUFx2_ASAP7_75t_R hold353 (.A(_04367_),
    .Y(net2477));
 BUFx2_ASAP7_75t_R hold354 (.A(net3079),
    .Y(net2478));
 BUFx2_ASAP7_75t_R hold355 (.A(net3083),
    .Y(net2479));
 BUFx2_ASAP7_75t_R hold356 (.A(_04459_),
    .Y(net2480));
 BUFx2_ASAP7_75t_R hold357 (.A(net4016),
    .Y(net2481));
 BUFx2_ASAP7_75t_R hold358 (.A(net3852),
    .Y(net2482));
 BUFx2_ASAP7_75t_R hold359 (.A(net3854),
    .Y(net2483));
 BUFx2_ASAP7_75t_R hold360 (.A(net2912),
    .Y(net2484));
 BUFx2_ASAP7_75t_R hold361 (.A(net2916),
    .Y(net2485));
 BUFx2_ASAP7_75t_R hold362 (.A(_04462_),
    .Y(net2486));
 BUFx2_ASAP7_75t_R hold363 (.A(net3922),
    .Y(net2487));
 BUFx2_ASAP7_75t_R hold364 (.A(net3926),
    .Y(net2488));
 BUFx2_ASAP7_75t_R hold365 (.A(net3928),
    .Y(net2489));
 BUFx2_ASAP7_75t_R hold366 (.A(net2904),
    .Y(net2490));
 BUFx2_ASAP7_75t_R hold367 (.A(net2908),
    .Y(net2491));
 BUFx2_ASAP7_75t_R hold368 (.A(_04466_),
    .Y(net2492));
 BUFx2_ASAP7_75t_R hold369 (.A(net4021),
    .Y(net2493));
 BUFx2_ASAP7_75t_R hold370 (.A(net3858),
    .Y(net2494));
 BUFx2_ASAP7_75t_R hold371 (.A(net3860),
    .Y(net2495));
 BUFx2_ASAP7_75t_R hold372 (.A(net4011),
    .Y(net2496));
 BUFx2_ASAP7_75t_R hold373 (.A(net3846),
    .Y(net2497));
 BUFx2_ASAP7_75t_R hold374 (.A(net3848),
    .Y(net2498));
 BUFx2_ASAP7_75t_R hold375 (.A(net2816),
    .Y(net2499));
 BUFx2_ASAP7_75t_R hold376 (.A(net2820),
    .Y(net2500));
 BUFx2_ASAP7_75t_R hold377 (.A(_04450_),
    .Y(net2501));
 BUFx2_ASAP7_75t_R hold378 (.A(net2761),
    .Y(net2502));
 BUFx2_ASAP7_75t_R hold379 (.A(net2763),
    .Y(net2503));
 BUFx2_ASAP7_75t_R hold380 (.A(net2765),
    .Y(net2504));
 BUFx2_ASAP7_75t_R hold381 (.A(net2767),
    .Y(net2505));
 BUFx2_ASAP7_75t_R hold382 (.A(net2925),
    .Y(net2506));
 BUFx2_ASAP7_75t_R hold383 (.A(net2929),
    .Y(net2507));
 BUFx2_ASAP7_75t_R hold384 (.A(_04460_),
    .Y(net2508));
 BUFx2_ASAP7_75t_R hold385 (.A(net4036),
    .Y(net2509));
 BUFx2_ASAP7_75t_R hold386 (.A(net3864),
    .Y(net2510));
 BUFx2_ASAP7_75t_R hold387 (.A(net3866),
    .Y(net2511));
 BUFx2_ASAP7_75t_R hold388 (.A(net2939),
    .Y(net2512));
 BUFx2_ASAP7_75t_R hold389 (.A(net2943),
    .Y(net2513));
 BUFx2_ASAP7_75t_R hold390 (.A(_04463_),
    .Y(net2514));
 BUFx2_ASAP7_75t_R hold391 (.A(net2947),
    .Y(net2515));
 BUFx2_ASAP7_75t_R hold392 (.A(net2951),
    .Y(net2516));
 BUFx2_ASAP7_75t_R hold393 (.A(_04447_),
    .Y(net2517));
 BUFx2_ASAP7_75t_R hold394 (.A(net3108),
    .Y(net2518));
 BUFx2_ASAP7_75t_R hold395 (.A(net3112),
    .Y(net2519));
 BUFx2_ASAP7_75t_R hold396 (.A(_04461_),
    .Y(net2520));
 BUFx2_ASAP7_75t_R hold397 (.A(net2774),
    .Y(net2521));
 BUFx2_ASAP7_75t_R hold398 (.A(net2776),
    .Y(net2522));
 BUFx2_ASAP7_75t_R hold399 (.A(net2778),
    .Y(net2523));
 BUFx2_ASAP7_75t_R hold400 (.A(net2780),
    .Y(net2524));
 BUFx2_ASAP7_75t_R hold401 (.A(net4031),
    .Y(net2525));
 BUFx2_ASAP7_75t_R hold402 (.A(net3870),
    .Y(net2526));
 BUFx2_ASAP7_75t_R hold403 (.A(net3872),
    .Y(net2527));
 BUFx2_ASAP7_75t_R hold404 (.A(net2963),
    .Y(net2528));
 BUFx2_ASAP7_75t_R hold405 (.A(net2967),
    .Y(net2529));
 BUFx2_ASAP7_75t_R hold406 (.A(_04469_),
    .Y(net2530));
 BUFx2_ASAP7_75t_R hold407 (.A(net3180),
    .Y(net2531));
 BUFx2_ASAP7_75t_R hold408 (.A(net3184),
    .Y(net2532));
 BUFx2_ASAP7_75t_R hold409 (.A(_02654_),
    .Y(net2533));
 BUFx2_ASAP7_75t_R hold410 (.A(net2855),
    .Y(net2534));
 BUFx2_ASAP7_75t_R hold411 (.A(net2857),
    .Y(net2535));
 BUFx2_ASAP7_75t_R hold412 (.A(net2859),
    .Y(net2536));
 BUFx2_ASAP7_75t_R hold413 (.A(net2861),
    .Y(net2537));
 BUFx2_ASAP7_75t_R hold414 (.A(net2782),
    .Y(net2538));
 BUFx2_ASAP7_75t_R hold415 (.A(net2784),
    .Y(net2539));
 BUFx2_ASAP7_75t_R hold416 (.A(net2786),
    .Y(net2540));
 BUFx2_ASAP7_75t_R hold417 (.A(net2788),
    .Y(net2541));
 BUFx2_ASAP7_75t_R hold418 (.A(net2955),
    .Y(net2542));
 BUFx2_ASAP7_75t_R hold419 (.A(net2959),
    .Y(net2543));
 BUFx2_ASAP7_75t_R hold420 (.A(_04440_),
    .Y(net2544));
 BUFx2_ASAP7_75t_R hold421 (.A(net2807),
    .Y(net2545));
 BUFx2_ASAP7_75t_R hold422 (.A(net2809),
    .Y(net2546));
 BUFx2_ASAP7_75t_R hold423 (.A(net2811),
    .Y(net2547));
 BUFx2_ASAP7_75t_R hold424 (.A(net2813),
    .Y(net2548));
 BUFx2_ASAP7_75t_R hold425 (.A(net4026),
    .Y(net2549));
 BUFx2_ASAP7_75t_R hold426 (.A(net3876),
    .Y(net2550));
 BUFx2_ASAP7_75t_R hold427 (.A(net3878),
    .Y(net2551));
 BUFx2_ASAP7_75t_R hold428 (.A(net3016),
    .Y(net2552));
 BUFx2_ASAP7_75t_R hold429 (.A(net3020),
    .Y(net2553));
 BUFx2_ASAP7_75t_R hold430 (.A(_04438_),
    .Y(net2554));
 BUFx2_ASAP7_75t_R hold431 (.A(net2823),
    .Y(net2555));
 BUFx2_ASAP7_75t_R hold432 (.A(net2825),
    .Y(net2556));
 BUFx2_ASAP7_75t_R hold433 (.A(net2827),
    .Y(net2557));
 BUFx2_ASAP7_75t_R hold434 (.A(net2829),
    .Y(net2558));
 BUFx2_ASAP7_75t_R hold435 (.A(net2980),
    .Y(net2559));
 BUFx2_ASAP7_75t_R hold436 (.A(net2984),
    .Y(net2560));
 BUFx2_ASAP7_75t_R hold437 (.A(_04445_),
    .Y(net2561));
 BUFx2_ASAP7_75t_R hold438 (.A(net4041),
    .Y(net2562));
 BUFx2_ASAP7_75t_R hold439 (.A(net3882),
    .Y(net2563));
 BUFx2_ASAP7_75t_R hold440 (.A(net3884),
    .Y(net2564));
 BUFx2_ASAP7_75t_R hold441 (.A(net3930),
    .Y(net2565));
 BUFx2_ASAP7_75t_R hold442 (.A(net3934),
    .Y(net2566));
 BUFx2_ASAP7_75t_R hold443 (.A(net3936),
    .Y(net2567));
 BUFx2_ASAP7_75t_R hold444 (.A(net4051),
    .Y(net2568));
 BUFx2_ASAP7_75t_R hold445 (.A(net3888),
    .Y(net2569));
 BUFx2_ASAP7_75t_R hold446 (.A(net3890),
    .Y(net2570));
 BUFx2_ASAP7_75t_R hold447 (.A(net4046),
    .Y(net2571));
 BUFx2_ASAP7_75t_R hold448 (.A(net3894),
    .Y(net2572));
 BUFx2_ASAP7_75t_R hold449 (.A(net3896),
    .Y(net2573));
 BUFx2_ASAP7_75t_R hold450 (.A(net2996),
    .Y(net2574));
 BUFx2_ASAP7_75t_R hold451 (.A(net3000),
    .Y(net2575));
 BUFx2_ASAP7_75t_R hold452 (.A(_04437_),
    .Y(net2576));
 BUFx2_ASAP7_75t_R hold453 (.A(net2839),
    .Y(net2577));
 BUFx2_ASAP7_75t_R hold454 (.A(net2841),
    .Y(net2578));
 BUFx2_ASAP7_75t_R hold455 (.A(net2843),
    .Y(net2579));
 BUFx2_ASAP7_75t_R hold456 (.A(net2845),
    .Y(net2580));
 BUFx2_ASAP7_75t_R hold457 (.A(net2831),
    .Y(net2581));
 BUFx2_ASAP7_75t_R hold458 (.A(net2833),
    .Y(net2582));
 BUFx2_ASAP7_75t_R hold459 (.A(net2835),
    .Y(net2583));
 BUFx2_ASAP7_75t_R hold460 (.A(net2837),
    .Y(net2584));
 BUFx2_ASAP7_75t_R hold461 (.A(net3004),
    .Y(net2585));
 BUFx2_ASAP7_75t_R hold462 (.A(net3008),
    .Y(net2586));
 BUFx2_ASAP7_75t_R hold463 (.A(_04456_),
    .Y(net2587));
 BUFx2_ASAP7_75t_R hold464 (.A(net2790),
    .Y(net2588));
 BUFx2_ASAP7_75t_R hold465 (.A(net2792),
    .Y(net2589));
 BUFx2_ASAP7_75t_R hold466 (.A(net2794),
    .Y(net2590));
 BUFx2_ASAP7_75t_R hold467 (.A(net2796),
    .Y(net2591));
 BUFx2_ASAP7_75t_R hold468 (.A(net2847),
    .Y(net2592));
 BUFx2_ASAP7_75t_R hold469 (.A(net2849),
    .Y(net2593));
 BUFx2_ASAP7_75t_R hold470 (.A(net2851),
    .Y(net2594));
 BUFx2_ASAP7_75t_R hold471 (.A(net2853),
    .Y(net2595));
 BUFx2_ASAP7_75t_R hold472 (.A(net2871),
    .Y(net2596));
 BUFx2_ASAP7_75t_R hold473 (.A(net2873),
    .Y(net2597));
 BUFx2_ASAP7_75t_R hold474 (.A(net2875),
    .Y(net2598));
 BUFx2_ASAP7_75t_R hold475 (.A(net2877),
    .Y(net2599));
 BUFx2_ASAP7_75t_R hold476 (.A(net2879),
    .Y(net2600));
 BUFx2_ASAP7_75t_R hold477 (.A(net2881),
    .Y(net2601));
 BUFx2_ASAP7_75t_R hold478 (.A(net2883),
    .Y(net2602));
 BUFx2_ASAP7_75t_R hold479 (.A(net2885),
    .Y(net2603));
 BUFx2_ASAP7_75t_R hold480 (.A(net2863),
    .Y(net2604));
 BUFx2_ASAP7_75t_R hold481 (.A(net2865),
    .Y(net2605));
 BUFx2_ASAP7_75t_R hold482 (.A(net2867),
    .Y(net2606));
 BUFx2_ASAP7_75t_R hold483 (.A(net2869),
    .Y(net2607));
 BUFx2_ASAP7_75t_R hold484 (.A(net2988),
    .Y(net2608));
 BUFx2_ASAP7_75t_R hold485 (.A(net2992),
    .Y(net2609));
 BUFx2_ASAP7_75t_R hold486 (.A(_04453_),
    .Y(net2610));
 BUFx2_ASAP7_75t_R hold487 (.A(net3070),
    .Y(net2611));
 BUFx2_ASAP7_75t_R hold488 (.A(net3072),
    .Y(net2612));
 BUFx2_ASAP7_75t_R hold489 (.A(net3074),
    .Y(net2613));
 BUFx2_ASAP7_75t_R hold490 (.A(net3076),
    .Y(net2614));
 BUFx2_ASAP7_75t_R hold491 (.A(net2887),
    .Y(net2615));
 BUFx2_ASAP7_75t_R hold492 (.A(net2889),
    .Y(net2616));
 BUFx2_ASAP7_75t_R hold493 (.A(net2891),
    .Y(net2617));
 BUFx2_ASAP7_75t_R hold494 (.A(net2893),
    .Y(net2618));
 BUFx2_ASAP7_75t_R hold495 (.A(net4056),
    .Y(net2619));
 BUFx2_ASAP7_75t_R hold496 (.A(net3900),
    .Y(net2620));
 BUFx2_ASAP7_75t_R hold497 (.A(net3902),
    .Y(net2621));
 BUFx2_ASAP7_75t_R hold498 (.A(net2895),
    .Y(net2622));
 BUFx2_ASAP7_75t_R hold499 (.A(net2897),
    .Y(net2623));
 BUFx2_ASAP7_75t_R hold500 (.A(net2899),
    .Y(net2624));
 BUFx2_ASAP7_75t_R hold501 (.A(net2901),
    .Y(net2625));
 BUFx2_ASAP7_75t_R hold502 (.A(net3078),
    .Y(net2626));
 BUFx2_ASAP7_75t_R hold503 (.A(net3080),
    .Y(net2627));
 BUFx2_ASAP7_75t_R hold504 (.A(net3082),
    .Y(net2628));
 BUFx2_ASAP7_75t_R hold505 (.A(net3084),
    .Y(net2629));
 BUFx2_ASAP7_75t_R hold506 (.A(net2815),
    .Y(net2630));
 BUFx2_ASAP7_75t_R hold507 (.A(net2817),
    .Y(net2631));
 BUFx2_ASAP7_75t_R hold508 (.A(net2819),
    .Y(net2632));
 BUFx2_ASAP7_75t_R hold509 (.A(net2821),
    .Y(net2633));
 BUFx2_ASAP7_75t_R hold510 (.A(net2903),
    .Y(net2634));
 BUFx2_ASAP7_75t_R hold511 (.A(net2905),
    .Y(net2635));
 BUFx2_ASAP7_75t_R hold512 (.A(net2907),
    .Y(net2636));
 BUFx2_ASAP7_75t_R hold513 (.A(net2909),
    .Y(net2637));
 BUFx2_ASAP7_75t_R hold514 (.A(net2924),
    .Y(net2638));
 BUFx2_ASAP7_75t_R hold515 (.A(net2926),
    .Y(net2639));
 BUFx2_ASAP7_75t_R hold516 (.A(net2928),
    .Y(net2640));
 BUFx2_ASAP7_75t_R hold517 (.A(net2930),
    .Y(net2641));
 BUFx2_ASAP7_75t_R hold518 (.A(net3754),
    .Y(net2642));
 BUFx2_ASAP7_75t_R hold519 (.A(net3758),
    .Y(net2643));
 BUFx2_ASAP7_75t_R hold520 (.A(_02647_),
    .Y(net2644));
 BUFx2_ASAP7_75t_R hold521 (.A(net2911),
    .Y(net2645));
 BUFx2_ASAP7_75t_R hold522 (.A(net2913),
    .Y(net2646));
 BUFx2_ASAP7_75t_R hold523 (.A(net2915),
    .Y(net2647));
 BUFx2_ASAP7_75t_R hold524 (.A(net2917),
    .Y(net2648));
 BUFx2_ASAP7_75t_R hold525 (.A(net3003),
    .Y(net2649));
 BUFx2_ASAP7_75t_R hold526 (.A(net3005),
    .Y(net2650));
 BUFx2_ASAP7_75t_R hold527 (.A(net3007),
    .Y(net2651));
 BUFx2_ASAP7_75t_R hold528 (.A(net3009),
    .Y(net2652));
 BUFx2_ASAP7_75t_R hold529 (.A(net3092),
    .Y(net2653));
 BUFx2_ASAP7_75t_R hold530 (.A(net3096),
    .Y(net2654));
 BUFx2_ASAP7_75t_R hold531 (.A(net2946),
    .Y(net2655));
 BUFx2_ASAP7_75t_R hold532 (.A(net2948),
    .Y(net2656));
 BUFx2_ASAP7_75t_R hold533 (.A(net2950),
    .Y(net2657));
 BUFx2_ASAP7_75t_R hold534 (.A(net2952),
    .Y(net2658));
 BUFx2_ASAP7_75t_R hold535 (.A(net2938),
    .Y(net2659));
 BUFx2_ASAP7_75t_R hold536 (.A(net2940),
    .Y(net2660));
 BUFx2_ASAP7_75t_R hold537 (.A(net2942),
    .Y(net2661));
 BUFx2_ASAP7_75t_R hold538 (.A(net2944),
    .Y(net2662));
 BUFx2_ASAP7_75t_R hold539 (.A(net3107),
    .Y(net2663));
 BUFx2_ASAP7_75t_R hold540 (.A(net3109),
    .Y(net2664));
 BUFx2_ASAP7_75t_R hold541 (.A(net3111),
    .Y(net2665));
 BUFx2_ASAP7_75t_R hold542 (.A(net3113),
    .Y(net2666));
 BUFx2_ASAP7_75t_R hold543 (.A(net2954),
    .Y(net2667));
 BUFx2_ASAP7_75t_R hold544 (.A(net2956),
    .Y(net2668));
 BUFx2_ASAP7_75t_R hold545 (.A(net2958),
    .Y(net2669));
 BUFx2_ASAP7_75t_R hold546 (.A(net2960),
    .Y(net2670));
 BUFx2_ASAP7_75t_R hold547 (.A(net3239),
    .Y(net2671));
 BUFx2_ASAP7_75t_R hold548 (.A(net3243),
    .Y(net2672));
 BUFx2_ASAP7_75t_R hold549 (.A(net3424),
    .Y(net2673));
 BUFx2_ASAP7_75t_R hold550 (.A(net3428),
    .Y(net2674));
 BUFx2_ASAP7_75t_R hold551 (.A(net3116),
    .Y(net2675));
 BUFx2_ASAP7_75t_R hold552 (.A(net3120),
    .Y(net2676));
 BUFx2_ASAP7_75t_R hold553 (.A(net3322),
    .Y(net2677));
 BUFx2_ASAP7_75t_R hold554 (.A(net3326),
    .Y(net2678));
 BUFx2_ASAP7_75t_R hold555 (.A(net2979),
    .Y(net2679));
 BUFx2_ASAP7_75t_R hold556 (.A(net2981),
    .Y(net2680));
 BUFx2_ASAP7_75t_R hold557 (.A(net2983),
    .Y(net2681));
 BUFx2_ASAP7_75t_R hold558 (.A(net2985),
    .Y(net2682));
 BUFx2_ASAP7_75t_R hold559 (.A(net3469),
    .Y(net2683));
 BUFx2_ASAP7_75t_R hold560 (.A(net3473),
    .Y(net2684));
 BUFx2_ASAP7_75t_R hold561 (.A(net2995),
    .Y(net2685));
 BUFx2_ASAP7_75t_R hold562 (.A(net2997),
    .Y(net2686));
 BUFx2_ASAP7_75t_R hold563 (.A(net2999),
    .Y(net2687));
 BUFx2_ASAP7_75t_R hold564 (.A(net3001),
    .Y(net2688));
 BUFx2_ASAP7_75t_R hold565 (.A(net2987),
    .Y(net2689));
 BUFx2_ASAP7_75t_R hold566 (.A(net2989),
    .Y(net2690));
 BUFx2_ASAP7_75t_R hold567 (.A(net2991),
    .Y(net2691));
 BUFx2_ASAP7_75t_R hold568 (.A(net2993),
    .Y(net2692));
 BUFx2_ASAP7_75t_R hold569 (.A(net3015),
    .Y(net2693));
 BUFx2_ASAP7_75t_R hold570 (.A(net3017),
    .Y(net2694));
 BUFx2_ASAP7_75t_R hold571 (.A(net3019),
    .Y(net2695));
 BUFx2_ASAP7_75t_R hold572 (.A(net3021),
    .Y(net2696));
 BUFx2_ASAP7_75t_R hold573 (.A(net3346),
    .Y(net2697));
 BUFx2_ASAP7_75t_R hold574 (.A(net3350),
    .Y(net2698));
 BUFx2_ASAP7_75t_R hold575 (.A(net3454),
    .Y(net2699));
 BUFx2_ASAP7_75t_R hold576 (.A(net3458),
    .Y(net2700));
 BUFx2_ASAP7_75t_R hold577 (.A(net3330),
    .Y(net2701));
 BUFx2_ASAP7_75t_R hold578 (.A(net3334),
    .Y(net2702));
 BUFx2_ASAP7_75t_R hold579 (.A(net3338),
    .Y(net2703));
 BUFx2_ASAP7_75t_R hold580 (.A(net3342),
    .Y(net2704));
 BUFx2_ASAP7_75t_R hold581 (.A(net3270),
    .Y(net2705));
 BUFx2_ASAP7_75t_R hold582 (.A(net3274),
    .Y(net2706));
 BUFx2_ASAP7_75t_R hold583 (.A(net3262),
    .Y(net2707));
 BUFx2_ASAP7_75t_R hold584 (.A(net3266),
    .Y(net2708));
 BUFx2_ASAP7_75t_R hold585 (.A(net3416),
    .Y(net2709));
 BUFx2_ASAP7_75t_R hold586 (.A(net3420),
    .Y(net2710));
 BUFx2_ASAP7_75t_R hold587 (.A(net3446),
    .Y(net2711));
 BUFx2_ASAP7_75t_R hold588 (.A(net3450),
    .Y(net2712));
 BUFx2_ASAP7_75t_R hold589 (.A(net2970),
    .Y(net2713));
 BUFx2_ASAP7_75t_R hold590 (.A(net2974),
    .Y(net2714));
 BUFx2_ASAP7_75t_R hold591 (.A(net2740),
    .Y(net2715));
 BUFx2_ASAP7_75t_R hold592 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .Y(net2716));
 BUFx2_ASAP7_75t_R hold593 (.A(net3247),
    .Y(net2717));
 BUFx2_ASAP7_75t_R hold594 (.A(net3251),
    .Y(net2718));
 BUFx2_ASAP7_75t_R hold595 (.A(net3360),
    .Y(net2719));
 BUFx2_ASAP7_75t_R hold596 (.A(net3364),
    .Y(net2720));
 BUFx2_ASAP7_75t_R hold597 (.A(net3314),
    .Y(net2721));
 BUFx2_ASAP7_75t_R hold598 (.A(net3318),
    .Y(net2722));
 BUFx2_ASAP7_75t_R hold599 (.A(net3278),
    .Y(net2723));
 BUFx2_ASAP7_75t_R hold600 (.A(net3282),
    .Y(net2724));
 BUFx2_ASAP7_75t_R hold601 (.A(net3462),
    .Y(net2725));
 BUFx2_ASAP7_75t_R hold602 (.A(net3466),
    .Y(net2726));
 BUFx2_ASAP7_75t_R hold603 (.A(net3046),
    .Y(net2727));
 BUFx2_ASAP7_75t_R hold604 (.A(net3050),
    .Y(net2728));
 BUFx2_ASAP7_75t_R hold605 (.A(net3307),
    .Y(net2729));
 BUFx2_ASAP7_75t_R hold606 (.A(net3311),
    .Y(net2730));
 BUFx2_ASAP7_75t_R hold607 (.A(net3727),
    .Y(net2731));
 BUFx2_ASAP7_75t_R hold608 (.A(net3035),
    .Y(net2732));
 BUFx2_ASAP7_75t_R hold609 (.A(_09314_),
    .Y(net2733));
 BUFx2_ASAP7_75t_R hold610 (.A(_09315_),
    .Y(net2734));
 BUFx2_ASAP7_75t_R hold611 (.A(_02830_),
    .Y(net2735));
 BUFx2_ASAP7_75t_R hold612 (.A(net2969),
    .Y(net2736));
 BUFx2_ASAP7_75t_R hold613 (.A(net2971),
    .Y(net2737));
 BUFx2_ASAP7_75t_R hold614 (.A(net2973),
    .Y(net2738));
 BUFx2_ASAP7_75t_R hold615 (.A(net2975),
    .Y(net2739));
 BUFx2_ASAP7_75t_R hold616 (.A(_06571_),
    .Y(net2740));
 BUFx2_ASAP7_75t_R hold617 (.A(net2715),
    .Y(net2741));
 BUFx2_ASAP7_75t_R hold618 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .Y(net2742));
 BUFx2_ASAP7_75t_R hold619 (.A(net3255),
    .Y(net2743));
 BUFx2_ASAP7_75t_R hold620 (.A(net3259),
    .Y(net2744));
 BUFx2_ASAP7_75t_R hold621 (.A(net3400),
    .Y(net2745));
 BUFx2_ASAP7_75t_R hold622 (.A(net3404),
    .Y(net2746));
 BUFx2_ASAP7_75t_R hold623 (.A(net3439),
    .Y(net2747));
 BUFx2_ASAP7_75t_R hold624 (.A(net3443),
    .Y(net2748));
 BUFx2_ASAP7_75t_R hold625 (.A(net3393),
    .Y(net2749));
 BUFx2_ASAP7_75t_R hold626 (.A(net3397),
    .Y(net2750));
 BUFx2_ASAP7_75t_R hold627 (.A(net3432),
    .Y(net2751));
 BUFx2_ASAP7_75t_R hold628 (.A(net3436),
    .Y(net2752));
 BUFx2_ASAP7_75t_R hold629 (.A(net3285),
    .Y(net2753));
 BUFx2_ASAP7_75t_R hold630 (.A(net3289),
    .Y(net2754));
 BUFx2_ASAP7_75t_R hold631 (.A(net3291),
    .Y(net2755));
 BUFx2_ASAP7_75t_R hold632 (.A(net3293),
    .Y(net2756));
 BUFx2_ASAP7_75t_R hold633 (.A(net3295),
    .Y(net2757));
 BUFx2_ASAP7_75t_R hold634 (.A(net3297),
    .Y(net2758));
 BUFx2_ASAP7_75t_R hold635 (.A(_06567_),
    .Y(net2759));
 BUFx2_ASAP7_75t_R hold636 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .Y(net2760));
 BUFx2_ASAP7_75t_R hold637 (.A(instr_rdata_i[15]),
    .Y(net2761));
 BUFx2_ASAP7_75t_R hold638 (.A(net2502),
    .Y(net2762));
 BUFx2_ASAP7_75t_R hold639 (.A(net2400),
    .Y(net2763));
 BUFx2_ASAP7_75t_R hold640 (.A(net2503),
    .Y(net2764));
 BUFx2_ASAP7_75t_R hold641 (.A(net102),
    .Y(net2765));
 BUFx2_ASAP7_75t_R hold642 (.A(net2504),
    .Y(net2766));
 BUFx2_ASAP7_75t_R hold643 (.A(net2401),
    .Y(net2767));
 BUFx2_ASAP7_75t_R hold644 (.A(net2505),
    .Y(net2768));
 BUFx2_ASAP7_75t_R hold645 (.A(net3091),
    .Y(net2769));
 BUFx2_ASAP7_75t_R hold646 (.A(net3093),
    .Y(net2770));
 BUFx2_ASAP7_75t_R hold647 (.A(net3095),
    .Y(net2771));
 BUFx2_ASAP7_75t_R hold648 (.A(net3097),
    .Y(net2772));
 BUFx2_ASAP7_75t_R hold649 (.A(_04457_),
    .Y(net2773));
 BUFx2_ASAP7_75t_R hold650 (.A(instr_rdata_i[28]),
    .Y(net2774));
 BUFx2_ASAP7_75t_R hold651 (.A(net2521),
    .Y(net2775));
 BUFx2_ASAP7_75t_R hold652 (.A(net2403),
    .Y(net2776));
 BUFx2_ASAP7_75t_R hold653 (.A(net2522),
    .Y(net2777));
 BUFx2_ASAP7_75t_R hold654 (.A(net116),
    .Y(net2778));
 BUFx2_ASAP7_75t_R hold655 (.A(net2523),
    .Y(net2779));
 BUFx2_ASAP7_75t_R hold656 (.A(net2404),
    .Y(net2780));
 BUFx2_ASAP7_75t_R hold657 (.A(net2524),
    .Y(net2781));
 BUFx2_ASAP7_75t_R hold658 (.A(instr_rdata_i[12]),
    .Y(net2782));
 BUFx2_ASAP7_75t_R hold659 (.A(net2538),
    .Y(net2783));
 BUFx2_ASAP7_75t_R hold660 (.A(net2406),
    .Y(net2784));
 BUFx2_ASAP7_75t_R hold661 (.A(net2539),
    .Y(net2785));
 BUFx2_ASAP7_75t_R hold662 (.A(net99),
    .Y(net2786));
 BUFx2_ASAP7_75t_R hold663 (.A(net2540),
    .Y(net2787));
 BUFx2_ASAP7_75t_R hold664 (.A(net2407),
    .Y(net2788));
 BUFx2_ASAP7_75t_R hold665 (.A(net2541),
    .Y(net2789));
 BUFx2_ASAP7_75t_R hold666 (.A(instr_rdata_i[9]),
    .Y(net2790));
 BUFx2_ASAP7_75t_R hold667 (.A(net2588),
    .Y(net2791));
 BUFx2_ASAP7_75t_R hold668 (.A(net2448),
    .Y(net2792));
 BUFx2_ASAP7_75t_R hold669 (.A(net2589),
    .Y(net2793));
 BUFx2_ASAP7_75t_R hold670 (.A(net127),
    .Y(net2794));
 BUFx2_ASAP7_75t_R hold671 (.A(net2590),
    .Y(net2795));
 BUFx2_ASAP7_75t_R hold672 (.A(net2449),
    .Y(net2796));
 BUFx2_ASAP7_75t_R hold673 (.A(net2591),
    .Y(net2797));
 BUFx2_ASAP7_75t_R hold674 (.A(net3115),
    .Y(net2798));
 BUFx2_ASAP7_75t_R hold675 (.A(net3117),
    .Y(net2799));
 BUFx2_ASAP7_75t_R hold676 (.A(net3119),
    .Y(net2800));
 BUFx2_ASAP7_75t_R hold677 (.A(net3121),
    .Y(net2801));
 BUFx2_ASAP7_75t_R hold678 (.A(_04441_),
    .Y(net2802));
 BUFx2_ASAP7_75t_R hold679 (.A(net3136),
    .Y(net2803));
 BUFx2_ASAP7_75t_R hold680 (.A(net3054),
    .Y(net2804));
 BUFx2_ASAP7_75t_R hold681 (.A(_09309_),
    .Y(net2805));
 BUFx2_ASAP7_75t_R hold682 (.A(_02829_),
    .Y(net2806));
 BUFx2_ASAP7_75t_R hold683 (.A(instr_rdata_i[30]),
    .Y(net2807));
 BUFx2_ASAP7_75t_R hold684 (.A(net2545),
    .Y(net2808));
 BUFx2_ASAP7_75t_R hold685 (.A(net2409),
    .Y(net2809));
 BUFx2_ASAP7_75t_R hold686 (.A(net2546),
    .Y(net2810));
 BUFx2_ASAP7_75t_R hold687 (.A(net119),
    .Y(net2811));
 BUFx2_ASAP7_75t_R hold688 (.A(net2547),
    .Y(net2812));
 BUFx2_ASAP7_75t_R hold689 (.A(net2410),
    .Y(net2813));
 BUFx2_ASAP7_75t_R hold690 (.A(net2548),
    .Y(net2814));
 BUFx2_ASAP7_75t_R hold691 (.A(instr_rdata_i[13]),
    .Y(net2815));
 BUFx2_ASAP7_75t_R hold692 (.A(net2630),
    .Y(net2816));
 BUFx2_ASAP7_75t_R hold693 (.A(net2499),
    .Y(net2817));
 BUFx2_ASAP7_75t_R hold694 (.A(net2631),
    .Y(net2818));
 BUFx2_ASAP7_75t_R hold695 (.A(net100),
    .Y(net2819));
 BUFx2_ASAP7_75t_R hold696 (.A(net2632),
    .Y(net2820));
 BUFx2_ASAP7_75t_R hold697 (.A(net2500),
    .Y(net2821));
 BUFx2_ASAP7_75t_R hold698 (.A(net2633),
    .Y(net2822));
 BUFx2_ASAP7_75t_R hold699 (.A(instr_rdata_i[14]),
    .Y(net2823));
 BUFx2_ASAP7_75t_R hold700 (.A(net2555),
    .Y(net2824));
 BUFx2_ASAP7_75t_R hold701 (.A(net2427),
    .Y(net2825));
 BUFx2_ASAP7_75t_R hold702 (.A(net2556),
    .Y(net2826));
 BUFx2_ASAP7_75t_R hold703 (.A(net101),
    .Y(net2827));
 BUFx2_ASAP7_75t_R hold704 (.A(net2557),
    .Y(net2828));
 BUFx2_ASAP7_75t_R hold705 (.A(net2428),
    .Y(net2829));
 BUFx2_ASAP7_75t_R hold706 (.A(net2558),
    .Y(net2830));
 BUFx2_ASAP7_75t_R hold707 (.A(instr_rdata_i[11]),
    .Y(net2831));
 BUFx2_ASAP7_75t_R hold708 (.A(net2581),
    .Y(net2832));
 BUFx2_ASAP7_75t_R hold709 (.A(net2430),
    .Y(net2833));
 BUFx2_ASAP7_75t_R hold710 (.A(net2582),
    .Y(net2834));
 BUFx2_ASAP7_75t_R hold711 (.A(net98),
    .Y(net2835));
 BUFx2_ASAP7_75t_R hold712 (.A(net2583),
    .Y(net2836));
 BUFx2_ASAP7_75t_R hold713 (.A(net2431),
    .Y(net2837));
 BUFx2_ASAP7_75t_R hold714 (.A(net2584),
    .Y(net2838));
 BUFx2_ASAP7_75t_R hold715 (.A(instr_rdata_i[2]),
    .Y(net2839));
 BUFx2_ASAP7_75t_R hold716 (.A(net2577),
    .Y(net2840));
 BUFx2_ASAP7_75t_R hold717 (.A(net2424),
    .Y(net2841));
 BUFx2_ASAP7_75t_R hold718 (.A(net2578),
    .Y(net2842));
 BUFx2_ASAP7_75t_R hold719 (.A(net118),
    .Y(net2843));
 BUFx2_ASAP7_75t_R hold720 (.A(net2579),
    .Y(net2844));
 BUFx2_ASAP7_75t_R hold721 (.A(net2425),
    .Y(net2845));
 BUFx2_ASAP7_75t_R hold722 (.A(net2580),
    .Y(net2846));
 BUFx2_ASAP7_75t_R hold723 (.A(instr_rdata_i[27]),
    .Y(net2847));
 BUFx2_ASAP7_75t_R hold724 (.A(net2592),
    .Y(net2848));
 BUFx2_ASAP7_75t_R hold725 (.A(net2454),
    .Y(net2849));
 BUFx2_ASAP7_75t_R hold726 (.A(net2593),
    .Y(net2850));
 BUFx2_ASAP7_75t_R hold727 (.A(net115),
    .Y(net2851));
 BUFx2_ASAP7_75t_R hold728 (.A(net2594),
    .Y(net2852));
 BUFx2_ASAP7_75t_R hold729 (.A(net2455),
    .Y(net2853));
 BUFx2_ASAP7_75t_R hold730 (.A(net2595),
    .Y(net2854));
 BUFx2_ASAP7_75t_R hold731 (.A(instr_rdata_i[31]),
    .Y(net2855));
 BUFx2_ASAP7_75t_R hold732 (.A(net2534),
    .Y(net2856));
 BUFx2_ASAP7_75t_R hold733 (.A(net2442),
    .Y(net2857));
 BUFx2_ASAP7_75t_R hold734 (.A(net2535),
    .Y(net2858));
 BUFx2_ASAP7_75t_R hold735 (.A(net120),
    .Y(net2859));
 BUFx2_ASAP7_75t_R hold736 (.A(net2536),
    .Y(net2860));
 BUFx2_ASAP7_75t_R hold737 (.A(net2443),
    .Y(net2861));
 BUFx2_ASAP7_75t_R hold738 (.A(net2537),
    .Y(net2862));
 BUFx2_ASAP7_75t_R hold739 (.A(instr_rdata_i[7]),
    .Y(net2863));
 BUFx2_ASAP7_75t_R hold740 (.A(net2604),
    .Y(net2864));
 BUFx2_ASAP7_75t_R hold741 (.A(net2469),
    .Y(net2865));
 BUFx2_ASAP7_75t_R hold742 (.A(net2605),
    .Y(net2866));
 BUFx2_ASAP7_75t_R hold743 (.A(net125),
    .Y(net2867));
 BUFx2_ASAP7_75t_R hold744 (.A(net2606),
    .Y(net2868));
 BUFx2_ASAP7_75t_R hold745 (.A(net2470),
    .Y(net2869));
 BUFx2_ASAP7_75t_R hold746 (.A(net2607),
    .Y(net2870));
 BUFx2_ASAP7_75t_R hold747 (.A(instr_rdata_i[21]),
    .Y(net2871));
 BUFx2_ASAP7_75t_R hold748 (.A(net2596),
    .Y(net2872));
 BUFx2_ASAP7_75t_R hold749 (.A(net2445),
    .Y(net2873));
 BUFx2_ASAP7_75t_R hold750 (.A(net2597),
    .Y(net2874));
 BUFx2_ASAP7_75t_R hold751 (.A(net109),
    .Y(net2875));
 BUFx2_ASAP7_75t_R hold752 (.A(net2598),
    .Y(net2876));
 BUFx2_ASAP7_75t_R hold753 (.A(net2446),
    .Y(net2877));
 BUFx2_ASAP7_75t_R hold754 (.A(net2599),
    .Y(net2878));
 BUFx2_ASAP7_75t_R hold755 (.A(instr_rdata_i[5]),
    .Y(net2879));
 BUFx2_ASAP7_75t_R hold756 (.A(net2600),
    .Y(net2880));
 BUFx2_ASAP7_75t_R hold757 (.A(net2451),
    .Y(net2881));
 BUFx2_ASAP7_75t_R hold758 (.A(net2601),
    .Y(net2882));
 BUFx2_ASAP7_75t_R hold759 (.A(net123),
    .Y(net2883));
 BUFx2_ASAP7_75t_R hold760 (.A(net2602),
    .Y(net2884));
 BUFx2_ASAP7_75t_R hold761 (.A(net2452),
    .Y(net2885));
 BUFx2_ASAP7_75t_R hold762 (.A(net2603),
    .Y(net2886));
 BUFx2_ASAP7_75t_R hold763 (.A(instr_rdata_i[18]),
    .Y(net2887));
 BUFx2_ASAP7_75t_R hold764 (.A(net2615),
    .Y(net2888));
 BUFx2_ASAP7_75t_R hold765 (.A(net2463),
    .Y(net2889));
 BUFx2_ASAP7_75t_R hold766 (.A(net2616),
    .Y(net2890));
 BUFx2_ASAP7_75t_R hold767 (.A(net105),
    .Y(net2891));
 BUFx2_ASAP7_75t_R hold768 (.A(net2617),
    .Y(net2892));
 BUFx2_ASAP7_75t_R hold769 (.A(net2464),
    .Y(net2893));
 BUFx2_ASAP7_75t_R hold770 (.A(net2618),
    .Y(net2894));
 BUFx2_ASAP7_75t_R hold771 (.A(instr_rdata_i[17]),
    .Y(net2895));
 BUFx2_ASAP7_75t_R hold772 (.A(net2622),
    .Y(net2896));
 BUFx2_ASAP7_75t_R hold773 (.A(net2472),
    .Y(net2897));
 BUFx2_ASAP7_75t_R hold774 (.A(net2623),
    .Y(net2898));
 BUFx2_ASAP7_75t_R hold775 (.A(net104),
    .Y(net2899));
 BUFx2_ASAP7_75t_R hold776 (.A(net2624),
    .Y(net2900));
 BUFx2_ASAP7_75t_R hold777 (.A(net2473),
    .Y(net2901));
 BUFx2_ASAP7_75t_R hold778 (.A(net2625),
    .Y(net2902));
 BUFx2_ASAP7_75t_R hold779 (.A(instr_rdata_i[29]),
    .Y(net2903));
 BUFx2_ASAP7_75t_R hold780 (.A(net2634),
    .Y(net2904));
 BUFx2_ASAP7_75t_R hold781 (.A(net2490),
    .Y(net2905));
 BUFx2_ASAP7_75t_R hold782 (.A(net2635),
    .Y(net2906));
 BUFx2_ASAP7_75t_R hold783 (.A(net117),
    .Y(net2907));
 BUFx2_ASAP7_75t_R hold784 (.A(net2636),
    .Y(net2908));
 BUFx2_ASAP7_75t_R hold785 (.A(net2491),
    .Y(net2909));
 BUFx2_ASAP7_75t_R hold786 (.A(net2637),
    .Y(net2910));
 BUFx2_ASAP7_75t_R hold787 (.A(instr_rdata_i[25]),
    .Y(net2911));
 BUFx2_ASAP7_75t_R hold788 (.A(net2645),
    .Y(net2912));
 BUFx2_ASAP7_75t_R hold789 (.A(net2484),
    .Y(net2913));
 BUFx2_ASAP7_75t_R hold790 (.A(net2646),
    .Y(net2914));
 BUFx2_ASAP7_75t_R hold791 (.A(net113),
    .Y(net2915));
 BUFx2_ASAP7_75t_R hold792 (.A(net2647),
    .Y(net2916));
 BUFx2_ASAP7_75t_R hold793 (.A(net2485),
    .Y(net2917));
 BUFx2_ASAP7_75t_R hold794 (.A(net2648),
    .Y(net2918));
 BUFx2_ASAP7_75t_R hold795 (.A(net3277),
    .Y(net2919));
 BUFx2_ASAP7_75t_R hold796 (.A(net3279),
    .Y(net2920));
 BUFx2_ASAP7_75t_R hold797 (.A(net3281),
    .Y(net2921));
 BUFx2_ASAP7_75t_R hold798 (.A(net3283),
    .Y(net2922));
 BUFx2_ASAP7_75t_R hold799 (.A(_06406_),
    .Y(net2923));
 BUFx2_ASAP7_75t_R hold800 (.A(instr_rdata_i[23]),
    .Y(net2924));
 BUFx2_ASAP7_75t_R hold801 (.A(net2638),
    .Y(net2925));
 BUFx2_ASAP7_75t_R hold802 (.A(net2506),
    .Y(net2926));
 BUFx2_ASAP7_75t_R hold803 (.A(net2639),
    .Y(net2927));
 BUFx2_ASAP7_75t_R hold804 (.A(net111),
    .Y(net2928));
 BUFx2_ASAP7_75t_R hold805 (.A(net2640),
    .Y(net2929));
 BUFx2_ASAP7_75t_R hold806 (.A(net2507),
    .Y(net2930));
 BUFx2_ASAP7_75t_R hold807 (.A(net2641),
    .Y(net2931));
 BUFx2_ASAP7_75t_R hold808 (.A(net2962),
    .Y(net2932));
 BUFx2_ASAP7_75t_R hold809 (.A(net2964),
    .Y(net2933));
 BUFx2_ASAP7_75t_R hold810 (.A(net2966),
    .Y(net2934));
 BUFx2_ASAP7_75t_R hold811 (.A(net2968),
    .Y(net2935));
 BUFx2_ASAP7_75t_R hold812 (.A(_06591_),
    .Y(net2936));
 BUFx2_ASAP7_75t_R hold813 (.A(_12673_),
    .Y(net2937));
 BUFx2_ASAP7_75t_R hold814 (.A(instr_rdata_i[26]),
    .Y(net2938));
 BUFx2_ASAP7_75t_R hold815 (.A(net2659),
    .Y(net2939));
 BUFx2_ASAP7_75t_R hold816 (.A(net2512),
    .Y(net2940));
 BUFx2_ASAP7_75t_R hold817 (.A(net2660),
    .Y(net2941));
 BUFx2_ASAP7_75t_R hold818 (.A(net114),
    .Y(net2942));
 BUFx2_ASAP7_75t_R hold819 (.A(net2661),
    .Y(net2943));
 BUFx2_ASAP7_75t_R hold820 (.A(net2513),
    .Y(net2944));
 BUFx2_ASAP7_75t_R hold821 (.A(net2662),
    .Y(net2945));
 BUFx2_ASAP7_75t_R hold822 (.A(instr_rdata_i[10]),
    .Y(net2946));
 BUFx2_ASAP7_75t_R hold823 (.A(net2655),
    .Y(net2947));
 BUFx2_ASAP7_75t_R hold824 (.A(net2515),
    .Y(net2948));
 BUFx2_ASAP7_75t_R hold825 (.A(net2656),
    .Y(net2949));
 BUFx2_ASAP7_75t_R hold826 (.A(net97),
    .Y(net2950));
 BUFx2_ASAP7_75t_R hold827 (.A(net2657),
    .Y(net2951));
 BUFx2_ASAP7_75t_R hold828 (.A(net2516),
    .Y(net2952));
 BUFx2_ASAP7_75t_R hold829 (.A(net2658),
    .Y(net2953));
 BUFx2_ASAP7_75t_R hold830 (.A(instr_rdata_i[3]),
    .Y(net2954));
 BUFx2_ASAP7_75t_R hold831 (.A(net2667),
    .Y(net2955));
 BUFx2_ASAP7_75t_R hold832 (.A(net2542),
    .Y(net2956));
 BUFx2_ASAP7_75t_R hold833 (.A(net2668),
    .Y(net2957));
 BUFx2_ASAP7_75t_R hold834 (.A(net121),
    .Y(net2958));
 BUFx2_ASAP7_75t_R hold835 (.A(net2669),
    .Y(net2959));
 BUFx2_ASAP7_75t_R hold836 (.A(net2543),
    .Y(net2960));
 BUFx2_ASAP7_75t_R hold837 (.A(net2670),
    .Y(net2961));
 BUFx2_ASAP7_75t_R hold838 (.A(instr_err_i),
    .Y(net2962));
 BUFx2_ASAP7_75t_R hold839 (.A(net2932),
    .Y(net2963));
 BUFx2_ASAP7_75t_R hold840 (.A(net2528),
    .Y(net2964));
 BUFx2_ASAP7_75t_R hold841 (.A(net2933),
    .Y(net2965));
 BUFx2_ASAP7_75t_R hold842 (.A(net94),
    .Y(net2966));
 BUFx2_ASAP7_75t_R hold843 (.A(net2934),
    .Y(net2967));
 BUFx2_ASAP7_75t_R hold844 (.A(net2529),
    .Y(net2968));
 BUFx2_ASAP7_75t_R hold845 (.A(instr_rvalid_i),
    .Y(net2969));
 BUFx2_ASAP7_75t_R hold846 (.A(net2736),
    .Y(net2970));
 BUFx2_ASAP7_75t_R hold847 (.A(net2713),
    .Y(net2971));
 BUFx2_ASAP7_75t_R hold848 (.A(net2737),
    .Y(net2972));
 BUFx2_ASAP7_75t_R hold849 (.A(net128),
    .Y(net2973));
 BUFx2_ASAP7_75t_R hold850 (.A(net2738),
    .Y(net2974));
 BUFx2_ASAP7_75t_R hold851 (.A(net2714),
    .Y(net2975));
 BUFx2_ASAP7_75t_R hold852 (.A(_06577_),
    .Y(net2976));
 BUFx2_ASAP7_75t_R hold853 (.A(_06578_),
    .Y(net2977));
 BUFx2_ASAP7_75t_R hold854 (.A(\if_stage_i.gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .Y(net2978));
 BUFx2_ASAP7_75t_R hold855 (.A(instr_rdata_i[8]),
    .Y(net2979));
 BUFx2_ASAP7_75t_R hold856 (.A(net2679),
    .Y(net2980));
 BUFx2_ASAP7_75t_R hold857 (.A(net2559),
    .Y(net2981));
 BUFx2_ASAP7_75t_R hold858 (.A(net2680),
    .Y(net2982));
 BUFx2_ASAP7_75t_R hold859 (.A(net126),
    .Y(net2983));
 BUFx2_ASAP7_75t_R hold860 (.A(net2681),
    .Y(net2984));
 BUFx2_ASAP7_75t_R hold861 (.A(net2560),
    .Y(net2985));
 BUFx2_ASAP7_75t_R hold862 (.A(net2682),
    .Y(net2986));
 BUFx2_ASAP7_75t_R hold863 (.A(instr_rdata_i[16]),
    .Y(net2987));
 BUFx2_ASAP7_75t_R hold864 (.A(net2689),
    .Y(net2988));
 BUFx2_ASAP7_75t_R hold865 (.A(net2608),
    .Y(net2989));
 BUFx2_ASAP7_75t_R hold866 (.A(net2690),
    .Y(net2990));
 BUFx2_ASAP7_75t_R hold867 (.A(net103),
    .Y(net2991));
 BUFx2_ASAP7_75t_R hold868 (.A(net2691),
    .Y(net2992));
 BUFx2_ASAP7_75t_R hold869 (.A(net2609),
    .Y(net2993));
 BUFx2_ASAP7_75t_R hold870 (.A(net2692),
    .Y(net2994));
 BUFx2_ASAP7_75t_R hold871 (.A(instr_rdata_i[0]),
    .Y(net2995));
 BUFx2_ASAP7_75t_R hold872 (.A(net2685),
    .Y(net2996));
 BUFx2_ASAP7_75t_R hold873 (.A(net2574),
    .Y(net2997));
 BUFx2_ASAP7_75t_R hold874 (.A(net2686),
    .Y(net2998));
 BUFx2_ASAP7_75t_R hold875 (.A(net96),
    .Y(net2999));
 BUFx2_ASAP7_75t_R hold876 (.A(net2687),
    .Y(net3000));
 BUFx2_ASAP7_75t_R hold877 (.A(net2575),
    .Y(net3001));
 BUFx2_ASAP7_75t_R hold878 (.A(net2688),
    .Y(net3002));
 BUFx2_ASAP7_75t_R hold879 (.A(instr_rdata_i[19]),
    .Y(net3003));
 BUFx2_ASAP7_75t_R hold880 (.A(net2649),
    .Y(net3004));
 BUFx2_ASAP7_75t_R hold881 (.A(net2585),
    .Y(net3005));
 BUFx2_ASAP7_75t_R hold882 (.A(net2650),
    .Y(net3006));
 BUFx2_ASAP7_75t_R hold883 (.A(net106),
    .Y(net3007));
 BUFx2_ASAP7_75t_R hold884 (.A(net2651),
    .Y(net3008));
 BUFx2_ASAP7_75t_R hold885 (.A(net2586),
    .Y(net3009));
 BUFx2_ASAP7_75t_R hold886 (.A(net2652),
    .Y(net3010));
 BUFx2_ASAP7_75t_R hold887 (.A(net3337),
    .Y(net3011));
 BUFx2_ASAP7_75t_R hold888 (.A(net3339),
    .Y(net3012));
 BUFx2_ASAP7_75t_R hold889 (.A(net3341),
    .Y(net3013));
 BUFx2_ASAP7_75t_R hold890 (.A(net3343),
    .Y(net3014));
 BUFx2_ASAP7_75t_R hold891 (.A(instr_rdata_i[1]),
    .Y(net3015));
 BUFx2_ASAP7_75t_R hold892 (.A(net2693),
    .Y(net3016));
 BUFx2_ASAP7_75t_R hold893 (.A(net2552),
    .Y(net3017));
 BUFx2_ASAP7_75t_R hold894 (.A(net2694),
    .Y(net3018));
 BUFx2_ASAP7_75t_R hold895 (.A(net107),
    .Y(net3019));
 BUFx2_ASAP7_75t_R hold896 (.A(net2695),
    .Y(net3020));
 BUFx2_ASAP7_75t_R hold897 (.A(net2553),
    .Y(net3021));
 BUFx2_ASAP7_75t_R hold898 (.A(net2696),
    .Y(net3022));
 BUFx2_ASAP7_75t_R hold899 (.A(net3284),
    .Y(net3023));
 BUFx2_ASAP7_75t_R hold900 (.A(net3286),
    .Y(net3024));
 BUFx2_ASAP7_75t_R hold901 (.A(net3288),
    .Y(net3025));
 BUFx2_ASAP7_75t_R hold902 (.A(net3290),
    .Y(net3026));
 BUFx2_ASAP7_75t_R hold903 (.A(net3045),
    .Y(net3027));
 BUFx2_ASAP7_75t_R hold904 (.A(net3047),
    .Y(net3028));
 BUFx2_ASAP7_75t_R hold905 (.A(net3049),
    .Y(net3029));
 BUFx2_ASAP7_75t_R hold906 (.A(net3051),
    .Y(net3030));
 BUFx2_ASAP7_75t_R hold907 (.A(_09301_),
    .Y(net3031));
 BUFx2_ASAP7_75t_R hold908 (.A(_02827_),
    .Y(net3032));
 BUFx2_ASAP7_75t_R hold909 (.A(net3726),
    .Y(net3033));
 BUFx2_ASAP7_75t_R hold910 (.A(net3728),
    .Y(net3034));
 BUFx2_ASAP7_75t_R hold911 (.A(net25),
    .Y(net3035));
 BUFx2_ASAP7_75t_R hold912 (.A(net2732),
    .Y(net3036));
 BUFx2_ASAP7_75t_R hold913 (.A(_05551_),
    .Y(net3037));
 BUFx2_ASAP7_75t_R hold914 (.A(net3057),
    .Y(net3038));
 BUFx2_ASAP7_75t_R hold915 (.A(\id_stage_i.controller_i.load_err_d ),
    .Y(net3039));
 BUFx2_ASAP7_75t_R hold916 (.A(net3313),
    .Y(net3040));
 BUFx2_ASAP7_75t_R hold917 (.A(net3315),
    .Y(net3041));
 BUFx2_ASAP7_75t_R hold918 (.A(net3317),
    .Y(net3042));
 BUFx2_ASAP7_75t_R hold919 (.A(net3319),
    .Y(net3043));
 BUFx2_ASAP7_75t_R hold920 (.A(_06449_),
    .Y(net3044));
 BUFx2_ASAP7_75t_R hold921 (.A(data_gnt_i),
    .Y(net3045));
 BUFx2_ASAP7_75t_R hold922 (.A(net3027),
    .Y(net3046));
 BUFx2_ASAP7_75t_R hold923 (.A(net2727),
    .Y(net3047));
 BUFx2_ASAP7_75t_R hold924 (.A(net3028),
    .Y(net3048));
 BUFx2_ASAP7_75t_R hold925 (.A(net26),
    .Y(net3049));
 BUFx2_ASAP7_75t_R hold926 (.A(net3029),
    .Y(net3050));
 BUFx2_ASAP7_75t_R hold927 (.A(net2728),
    .Y(net3051));
 BUFx2_ASAP7_75t_R hold928 (.A(net3135),
    .Y(net3052));
 BUFx2_ASAP7_75t_R hold929 (.A(net3137),
    .Y(net3053));
 BUFx2_ASAP7_75t_R hold930 (.A(net59),
    .Y(net3054));
 BUFx2_ASAP7_75t_R hold931 (.A(net2804),
    .Y(net3055));
 BUFx2_ASAP7_75t_R hold932 (.A(_05553_),
    .Y(net3056));
 BUFx2_ASAP7_75t_R hold933 (.A(_05554_),
    .Y(net3057));
 BUFx2_ASAP7_75t_R hold934 (.A(net3038),
    .Y(net3058));
 BUFx2_ASAP7_75t_R hold935 (.A(\id_stage_i.controller_i.store_err_d ),
    .Y(net3059));
 BUFx2_ASAP7_75t_R hold936 (.A(net3261),
    .Y(net3060));
 BUFx2_ASAP7_75t_R hold937 (.A(net3263),
    .Y(net3061));
 BUFx2_ASAP7_75t_R hold938 (.A(net3265),
    .Y(net3062));
 BUFx2_ASAP7_75t_R hold939 (.A(net3267),
    .Y(net3063));
 BUFx2_ASAP7_75t_R hold940 (.A(_06552_),
    .Y(net3064));
 BUFx2_ASAP7_75t_R hold941 (.A(_06556_),
    .Y(net3065));
 BUFx2_ASAP7_75t_R hold942 (.A(net3945),
    .Y(net3066));
 BUFx2_ASAP7_75t_R hold943 (.A(net3947),
    .Y(net3067));
 BUFx2_ASAP7_75t_R hold944 (.A(net3949),
    .Y(net3068));
 BUFx2_ASAP7_75t_R hold945 (.A(net3951),
    .Y(net3069));
 BUFx2_ASAP7_75t_R hold946 (.A(instr_rdata_i[6]),
    .Y(net3070));
 BUFx2_ASAP7_75t_R hold947 (.A(net2611),
    .Y(net3071));
 BUFx2_ASAP7_75t_R hold948 (.A(net2466),
    .Y(net3072));
 BUFx2_ASAP7_75t_R hold949 (.A(net2612),
    .Y(net3073));
 BUFx2_ASAP7_75t_R hold950 (.A(net124),
    .Y(net3074));
 BUFx2_ASAP7_75t_R hold951 (.A(net2613),
    .Y(net3075));
 BUFx2_ASAP7_75t_R hold952 (.A(net2467),
    .Y(net3076));
 BUFx2_ASAP7_75t_R hold953 (.A(net2614),
    .Y(net3077));
 BUFx2_ASAP7_75t_R hold954 (.A(instr_rdata_i[22]),
    .Y(net3078));
 BUFx2_ASAP7_75t_R hold955 (.A(net2626),
    .Y(net3079));
 BUFx2_ASAP7_75t_R hold956 (.A(net2478),
    .Y(net3080));
 BUFx2_ASAP7_75t_R hold957 (.A(net2627),
    .Y(net3081));
 BUFx2_ASAP7_75t_R hold958 (.A(net110),
    .Y(net3082));
 BUFx2_ASAP7_75t_R hold959 (.A(net2628),
    .Y(net3083));
 BUFx2_ASAP7_75t_R hold960 (.A(net2479),
    .Y(net3084));
 BUFx2_ASAP7_75t_R hold961 (.A(net2629),
    .Y(net3085));
 BUFx2_ASAP7_75t_R hold962 (.A(net3415),
    .Y(net3086));
 BUFx2_ASAP7_75t_R hold963 (.A(net3417),
    .Y(net3087));
 BUFx2_ASAP7_75t_R hold964 (.A(net3419),
    .Y(net3088));
 BUFx2_ASAP7_75t_R hold965 (.A(net3421),
    .Y(net3089));
 BUFx2_ASAP7_75t_R hold966 (.A(_06389_),
    .Y(net3090));
 BUFx2_ASAP7_75t_R hold967 (.A(instr_rdata_i[20]),
    .Y(net3091));
 BUFx2_ASAP7_75t_R hold968 (.A(net2769),
    .Y(net3092));
 BUFx2_ASAP7_75t_R hold969 (.A(net2653),
    .Y(net3093));
 BUFx2_ASAP7_75t_R hold970 (.A(net2770),
    .Y(net3094));
 BUFx2_ASAP7_75t_R hold971 (.A(net108),
    .Y(net3095));
 BUFx2_ASAP7_75t_R hold972 (.A(net2771),
    .Y(net3096));
 BUFx2_ASAP7_75t_R hold973 (.A(net2654),
    .Y(net3097));
 BUFx2_ASAP7_75t_R hold974 (.A(net2772),
    .Y(net3098));
 BUFx2_ASAP7_75t_R hold975 (.A(net3179),
    .Y(net3099));
 BUFx2_ASAP7_75t_R hold976 (.A(net3181),
    .Y(net3100));
 BUFx2_ASAP7_75t_R hold977 (.A(net3183),
    .Y(net3101));
 BUFx2_ASAP7_75t_R hold978 (.A(net3185),
    .Y(net3102));
 BUFx2_ASAP7_75t_R hold979 (.A(_06670_),
    .Y(net3103));
 BUFx2_ASAP7_75t_R hold980 (.A(_06671_),
    .Y(net3104));
 BUFx2_ASAP7_75t_R hold981 (.A(net3133),
    .Y(net3105));
 BUFx2_ASAP7_75t_R hold982 (.A(_06684_),
    .Y(net3106));
 BUFx2_ASAP7_75t_R hold983 (.A(instr_rdata_i[24]),
    .Y(net3107));
 BUFx2_ASAP7_75t_R hold984 (.A(net2663),
    .Y(net3108));
 BUFx2_ASAP7_75t_R hold985 (.A(net2518),
    .Y(net3109));
 BUFx2_ASAP7_75t_R hold986 (.A(net2664),
    .Y(net3110));
 BUFx2_ASAP7_75t_R hold987 (.A(net112),
    .Y(net3111));
 BUFx2_ASAP7_75t_R hold988 (.A(net2665),
    .Y(net3112));
 BUFx2_ASAP7_75t_R hold989 (.A(net2519),
    .Y(net3113));
 BUFx2_ASAP7_75t_R hold990 (.A(net2666),
    .Y(net3114));
 BUFx2_ASAP7_75t_R hold991 (.A(instr_rdata_i[4]),
    .Y(net3115));
 BUFx2_ASAP7_75t_R hold992 (.A(net2798),
    .Y(net3116));
 BUFx2_ASAP7_75t_R hold993 (.A(net2675),
    .Y(net3117));
 BUFx2_ASAP7_75t_R hold994 (.A(net2799),
    .Y(net3118));
 BUFx2_ASAP7_75t_R hold995 (.A(net122),
    .Y(net3119));
 BUFx2_ASAP7_75t_R hold996 (.A(net2800),
    .Y(net3120));
 BUFx2_ASAP7_75t_R hold997 (.A(net2676),
    .Y(net3121));
 BUFx2_ASAP7_75t_R hold998 (.A(net2801),
    .Y(net3122));
 BUFx2_ASAP7_75t_R hold999 (.A(net3431),
    .Y(net3123));
 BUFx2_ASAP7_75t_R hold1000 (.A(net3433),
    .Y(net3124));
 BUFx2_ASAP7_75t_R hold1001 (.A(net3435),
    .Y(net3125));
 BUFx2_ASAP7_75t_R hold1002 (.A(net3437),
    .Y(net3126));
 BUFx2_ASAP7_75t_R hold1003 (.A(_06394_),
    .Y(net3127));
 BUFx2_ASAP7_75t_R hold1004 (.A(net3753),
    .Y(net3128));
 BUFx2_ASAP7_75t_R hold1005 (.A(net3755),
    .Y(net3129));
 BUFx2_ASAP7_75t_R hold1006 (.A(net3757),
    .Y(net3130));
 BUFx2_ASAP7_75t_R hold1007 (.A(net2643),
    .Y(net3131));
 BUFx2_ASAP7_75t_R hold1008 (.A(_06237_),
    .Y(net3132));
 BUFx2_ASAP7_75t_R hold1009 (.A(_06672_),
    .Y(net3133));
 BUFx2_ASAP7_75t_R hold1010 (.A(net3105),
    .Y(net3134));
 BUFx2_ASAP7_75t_R hold1011 (.A(data_rvalid_i),
    .Y(net3135));
 BUFx2_ASAP7_75t_R hold1012 (.A(net3052),
    .Y(net3136));
 BUFx2_ASAP7_75t_R hold1013 (.A(net2803),
    .Y(net3137));
 BUFx2_ASAP7_75t_R hold1014 (.A(net3053),
    .Y(net3138));
 BUFx2_ASAP7_75t_R hold1015 (.A(net3960),
    .Y(net3139));
 BUFx2_ASAP7_75t_R hold1016 (.A(net3962),
    .Y(net3140));
 BUFx2_ASAP7_75t_R hold1017 (.A(net3964),
    .Y(net3141));
 BUFx2_ASAP7_75t_R hold1018 (.A(net3966),
    .Y(net3142));
 BUFx2_ASAP7_75t_R hold1019 (.A(net3321),
    .Y(net3143));
 BUFx2_ASAP7_75t_R hold1020 (.A(net3323),
    .Y(net3144));
 BUFx2_ASAP7_75t_R hold1021 (.A(net3325),
    .Y(net3145));
 BUFx2_ASAP7_75t_R hold1022 (.A(net3327),
    .Y(net3146));
 BUFx2_ASAP7_75t_R hold1023 (.A(_06525_),
    .Y(net3147));
 BUFx2_ASAP7_75t_R hold1024 (.A(net3238),
    .Y(net3148));
 BUFx2_ASAP7_75t_R hold1025 (.A(net3240),
    .Y(net3149));
 BUFx2_ASAP7_75t_R hold1026 (.A(net3242),
    .Y(net3150));
 BUFx2_ASAP7_75t_R hold1027 (.A(net3244),
    .Y(net3151));
 BUFx2_ASAP7_75t_R hold1028 (.A(_06534_),
    .Y(net3152));
 BUFx2_ASAP7_75t_R hold1029 (.A(net3359),
    .Y(net3153));
 BUFx2_ASAP7_75t_R hold1030 (.A(net3361),
    .Y(net3154));
 BUFx2_ASAP7_75t_R hold1031 (.A(net3363),
    .Y(net3155));
 BUFx2_ASAP7_75t_R hold1032 (.A(net3365),
    .Y(net3156));
 BUFx2_ASAP7_75t_R hold1033 (.A(_06510_),
    .Y(net3157));
 BUFx2_ASAP7_75t_R hold1034 (.A(net3453),
    .Y(net3158));
 BUFx2_ASAP7_75t_R hold1035 (.A(net3455),
    .Y(net3159));
 BUFx2_ASAP7_75t_R hold1036 (.A(net3457),
    .Y(net3160));
 BUFx2_ASAP7_75t_R hold1037 (.A(net3459),
    .Y(net3161));
 BUFx2_ASAP7_75t_R hold1038 (.A(_06419_),
    .Y(net3162));
 BUFx2_ASAP7_75t_R hold1039 (.A(net3468),
    .Y(net3163));
 BUFx2_ASAP7_75t_R hold1040 (.A(net3470),
    .Y(net3164));
 BUFx2_ASAP7_75t_R hold1041 (.A(net3472),
    .Y(net3165));
 BUFx2_ASAP7_75t_R hold1042 (.A(net3474),
    .Y(net3166));
 BUFx2_ASAP7_75t_R hold1043 (.A(_06436_),
    .Y(net3167));
 BUFx2_ASAP7_75t_R hold1044 (.A(_06440_),
    .Y(net3168));
 BUFx2_ASAP7_75t_R hold1045 (.A(net3423),
    .Y(net3169));
 BUFx2_ASAP7_75t_R hold1046 (.A(net3425),
    .Y(net3170));
 BUFx2_ASAP7_75t_R hold1047 (.A(net3427),
    .Y(net3171));
 BUFx2_ASAP7_75t_R hold1048 (.A(net3429),
    .Y(net3172));
 BUFx2_ASAP7_75t_R hold1049 (.A(_06471_),
    .Y(net3173));
 BUFx2_ASAP7_75t_R hold1050 (.A(net3438),
    .Y(net3174));
 BUFx2_ASAP7_75t_R hold1051 (.A(net3440),
    .Y(net3175));
 BUFx2_ASAP7_75t_R hold1052 (.A(net3442),
    .Y(net3176));
 BUFx2_ASAP7_75t_R hold1053 (.A(net3444),
    .Y(net3177));
 BUFx2_ASAP7_75t_R hold1054 (.A(_06505_),
    .Y(net3178));
 BUFx2_ASAP7_75t_R hold1055 (.A(debug_req_i),
    .Y(net3179));
 BUFx2_ASAP7_75t_R hold1056 (.A(net3099),
    .Y(net3180));
 BUFx2_ASAP7_75t_R hold1057 (.A(net2531),
    .Y(net3181));
 BUFx2_ASAP7_75t_R hold1058 (.A(net3100),
    .Y(net3182));
 BUFx2_ASAP7_75t_R hold1059 (.A(net60),
    .Y(net3183));
 BUFx2_ASAP7_75t_R hold1060 (.A(net3101),
    .Y(net3184));
 BUFx2_ASAP7_75t_R hold1061 (.A(net2532),
    .Y(net3185));
 BUFx2_ASAP7_75t_R hold1062 (.A(net3392),
    .Y(net3186));
 BUFx2_ASAP7_75t_R hold1063 (.A(net3394),
    .Y(net3187));
 BUFx2_ASAP7_75t_R hold1064 (.A(net3396),
    .Y(net3188));
 BUFx2_ASAP7_75t_R hold1065 (.A(net3398),
    .Y(net3189));
 BUFx2_ASAP7_75t_R hold1066 (.A(_06540_),
    .Y(net3190));
 BUFx2_ASAP7_75t_R hold1067 (.A(net3445),
    .Y(net3191));
 BUFx2_ASAP7_75t_R hold1068 (.A(net3447),
    .Y(net3192));
 BUFx2_ASAP7_75t_R hold1069 (.A(net3449),
    .Y(net3193));
 BUFx2_ASAP7_75t_R hold1070 (.A(net3451),
    .Y(net3194));
 BUFx2_ASAP7_75t_R hold1071 (.A(_06442_),
    .Y(net3195));
 BUFx2_ASAP7_75t_R hold1072 (.A(net3461),
    .Y(net3196));
 BUFx2_ASAP7_75t_R hold1073 (.A(net3463),
    .Y(net3197));
 BUFx2_ASAP7_75t_R hold1074 (.A(net3465),
    .Y(net3198));
 BUFx2_ASAP7_75t_R hold1075 (.A(net3467),
    .Y(net3199));
 BUFx2_ASAP7_75t_R hold1076 (.A(_06457_),
    .Y(net3200));
 BUFx2_ASAP7_75t_R hold1077 (.A(net3269),
    .Y(net3201));
 BUFx2_ASAP7_75t_R hold1078 (.A(net3271),
    .Y(net3202));
 BUFx2_ASAP7_75t_R hold1079 (.A(net3273),
    .Y(net3203));
 BUFx2_ASAP7_75t_R hold1080 (.A(net3275),
    .Y(net3204));
 BUFx2_ASAP7_75t_R hold1081 (.A(_06478_),
    .Y(net3205));
 BUFx2_ASAP7_75t_R hold1082 (.A(net3656),
    .Y(net3206));
 BUFx2_ASAP7_75t_R hold1083 (.A(net147),
    .Y(net3207));
 BUFx2_ASAP7_75t_R hold1084 (.A(_06268_),
    .Y(net3208));
 BUFx2_ASAP7_75t_R hold1085 (.A(_06269_),
    .Y(net3209));
 BUFx2_ASAP7_75t_R hold1086 (.A(net3357),
    .Y(net3210));
 BUFx2_ASAP7_75t_R hold1087 (.A(_06271_),
    .Y(net3211));
 BUFx2_ASAP7_75t_R hold1088 (.A(net3399),
    .Y(net3212));
 BUFx2_ASAP7_75t_R hold1089 (.A(net3401),
    .Y(net3213));
 BUFx2_ASAP7_75t_R hold1090 (.A(net3403),
    .Y(net3214));
 BUFx2_ASAP7_75t_R hold1091 (.A(net3405),
    .Y(net3215));
 BUFx2_ASAP7_75t_R hold1092 (.A(_06497_),
    .Y(net3216));
 BUFx2_ASAP7_75t_R hold1093 (.A(net3306),
    .Y(net3217));
 BUFx2_ASAP7_75t_R hold1094 (.A(net3308),
    .Y(net3218));
 BUFx2_ASAP7_75t_R hold1095 (.A(net3310),
    .Y(net3219));
 BUFx2_ASAP7_75t_R hold1096 (.A(net3312),
    .Y(net3220));
 BUFx2_ASAP7_75t_R hold1097 (.A(net3246),
    .Y(net3221));
 BUFx2_ASAP7_75t_R hold1098 (.A(net3248),
    .Y(net3222));
 BUFx2_ASAP7_75t_R hold1099 (.A(net3250),
    .Y(net3223));
 BUFx2_ASAP7_75t_R hold1100 (.A(net3252),
    .Y(net3224));
 BUFx2_ASAP7_75t_R hold1101 (.A(_06431_),
    .Y(net3225));
 BUFx2_ASAP7_75t_R hold1102 (.A(net3254),
    .Y(net3226));
 BUFx2_ASAP7_75t_R hold1103 (.A(net3256),
    .Y(net3227));
 BUFx2_ASAP7_75t_R hold1104 (.A(net3258),
    .Y(net3228));
 BUFx2_ASAP7_75t_R hold1105 (.A(net3260),
    .Y(net3229));
 BUFx2_ASAP7_75t_R hold1106 (.A(net3329),
    .Y(net3230));
 BUFx2_ASAP7_75t_R hold1107 (.A(net3331),
    .Y(net3231));
 BUFx2_ASAP7_75t_R hold1108 (.A(net3333),
    .Y(net3232));
 BUFx2_ASAP7_75t_R hold1109 (.A(net3335),
    .Y(net3233));
 BUFx2_ASAP7_75t_R hold1110 (.A(net3345),
    .Y(net3234));
 BUFx2_ASAP7_75t_R hold1111 (.A(net3347),
    .Y(net3235));
 BUFx2_ASAP7_75t_R hold1112 (.A(net3349),
    .Y(net3236));
 BUFx2_ASAP7_75t_R hold1113 (.A(net3351),
    .Y(net3237));
 BUFx2_ASAP7_75t_R hold1114 (.A(boot_addr_i[28]),
    .Y(net3238));
 BUFx2_ASAP7_75t_R hold1115 (.A(net3148),
    .Y(net3239));
 BUFx2_ASAP7_75t_R hold1116 (.A(net2671),
    .Y(net3240));
 BUFx2_ASAP7_75t_R hold1117 (.A(net3149),
    .Y(net3241));
 BUFx2_ASAP7_75t_R hold1118 (.A(net19),
    .Y(net3242));
 BUFx2_ASAP7_75t_R hold1119 (.A(net3150),
    .Y(net3243));
 BUFx2_ASAP7_75t_R hold1120 (.A(net2672),
    .Y(net3244));
 BUFx2_ASAP7_75t_R hold1121 (.A(net3151),
    .Y(net3245));
 BUFx2_ASAP7_75t_R hold1122 (.A(boot_addr_i[13]),
    .Y(net3246));
 BUFx2_ASAP7_75t_R hold1123 (.A(net3221),
    .Y(net3247));
 BUFx2_ASAP7_75t_R hold1124 (.A(net2717),
    .Y(net3248));
 BUFx2_ASAP7_75t_R hold1125 (.A(net3222),
    .Y(net3249));
 BUFx2_ASAP7_75t_R hold1126 (.A(net4),
    .Y(net3250));
 BUFx2_ASAP7_75t_R hold1127 (.A(net3223),
    .Y(net3251));
 BUFx2_ASAP7_75t_R hold1128 (.A(net2718),
    .Y(net3252));
 BUFx2_ASAP7_75t_R hold1129 (.A(net3224),
    .Y(net3253));
 BUFx2_ASAP7_75t_R hold1130 (.A(boot_addr_i[30]),
    .Y(net3254));
 BUFx2_ASAP7_75t_R hold1131 (.A(net3226),
    .Y(net3255));
 BUFx2_ASAP7_75t_R hold1132 (.A(net2743),
    .Y(net3256));
 BUFx2_ASAP7_75t_R hold1133 (.A(net3227),
    .Y(net3257));
 BUFx2_ASAP7_75t_R hold1134 (.A(net21),
    .Y(net3258));
 BUFx2_ASAP7_75t_R hold1135 (.A(net3228),
    .Y(net3259));
 BUFx2_ASAP7_75t_R hold1136 (.A(net2744),
    .Y(net3260));
 BUFx2_ASAP7_75t_R hold1137 (.A(boot_addr_i[31]),
    .Y(net3261));
 BUFx2_ASAP7_75t_R hold1138 (.A(net3060),
    .Y(net3262));
 BUFx2_ASAP7_75t_R hold1139 (.A(net2707),
    .Y(net3263));
 BUFx2_ASAP7_75t_R hold1140 (.A(net3061),
    .Y(net3264));
 BUFx2_ASAP7_75t_R hold1141 (.A(net22),
    .Y(net3265));
 BUFx2_ASAP7_75t_R hold1142 (.A(net3062),
    .Y(net3266));
 BUFx2_ASAP7_75t_R hold1143 (.A(net2708),
    .Y(net3267));
 BUFx2_ASAP7_75t_R hold1144 (.A(net3063),
    .Y(net3268));
 BUFx2_ASAP7_75t_R hold1145 (.A(boot_addr_i[20]),
    .Y(net3269));
 BUFx2_ASAP7_75t_R hold1146 (.A(net3201),
    .Y(net3270));
 BUFx2_ASAP7_75t_R hold1147 (.A(net2705),
    .Y(net3271));
 BUFx2_ASAP7_75t_R hold1148 (.A(net3202),
    .Y(net3272));
 BUFx2_ASAP7_75t_R hold1149 (.A(net11),
    .Y(net3273));
 BUFx2_ASAP7_75t_R hold1150 (.A(net3203),
    .Y(net3274));
 BUFx2_ASAP7_75t_R hold1151 (.A(net2706),
    .Y(net3275));
 BUFx2_ASAP7_75t_R hold1152 (.A(net3204),
    .Y(net3276));
 BUFx2_ASAP7_75t_R hold1153 (.A(boot_addr_i[11]),
    .Y(net3277));
 BUFx2_ASAP7_75t_R hold1154 (.A(net2919),
    .Y(net3278));
 BUFx2_ASAP7_75t_R hold1155 (.A(net2723),
    .Y(net3279));
 BUFx2_ASAP7_75t_R hold1156 (.A(net2920),
    .Y(net3280));
 BUFx2_ASAP7_75t_R hold1157 (.A(net2),
    .Y(net3281));
 BUFx2_ASAP7_75t_R hold1158 (.A(net2921),
    .Y(net3282));
 BUFx2_ASAP7_75t_R hold1159 (.A(net2724),
    .Y(net3283));
 BUFx2_ASAP7_75t_R hold1160 (.A(boot_addr_i[10]),
    .Y(net3284));
 BUFx2_ASAP7_75t_R hold1161 (.A(net3023),
    .Y(net3285));
 BUFx2_ASAP7_75t_R hold1162 (.A(net2753),
    .Y(net3286));
 BUFx2_ASAP7_75t_R hold1163 (.A(net3024),
    .Y(net3287));
 BUFx2_ASAP7_75t_R hold1164 (.A(net1),
    .Y(net3288));
 BUFx2_ASAP7_75t_R hold1165 (.A(net3025),
    .Y(net3289));
 BUFx2_ASAP7_75t_R hold1166 (.A(net2754),
    .Y(net3290));
 BUFx2_ASAP7_75t_R hold1167 (.A(instr_gnt_i),
    .Y(net3291));
 BUFx2_ASAP7_75t_R hold1168 (.A(net2755),
    .Y(net3292));
 BUFx2_ASAP7_75t_R hold1169 (.A(net2460),
    .Y(net3293));
 BUFx2_ASAP7_75t_R hold1170 (.A(net2756),
    .Y(net3294));
 BUFx2_ASAP7_75t_R hold1171 (.A(net95),
    .Y(net3295));
 BUFx2_ASAP7_75t_R hold1172 (.A(net2757),
    .Y(net3296));
 BUFx2_ASAP7_75t_R hold1173 (.A(net2461),
    .Y(net3297));
 BUFx2_ASAP7_75t_R hold1174 (.A(net3669),
    .Y(net3298));
 BUFx2_ASAP7_75t_R hold1175 (.A(net130),
    .Y(net3299));
 BUFx2_ASAP7_75t_R hold1176 (.A(_06250_),
    .Y(net3300));
 BUFx2_ASAP7_75t_R hold1177 (.A(net3494),
    .Y(net3301));
 BUFx2_ASAP7_75t_R hold1178 (.A(_06607_),
    .Y(net3302));
 BUFx2_ASAP7_75t_R hold1179 (.A(_06714_),
    .Y(net3303));
 BUFx2_ASAP7_75t_R hold1180 (.A(_06897_),
    .Y(net3304));
 BUFx2_ASAP7_75t_R hold1181 (.A(_06912_),
    .Y(net3305));
 BUFx2_ASAP7_75t_R hold1182 (.A(boot_addr_i[22]),
    .Y(net3306));
 BUFx2_ASAP7_75t_R hold1183 (.A(net3217),
    .Y(net3307));
 BUFx2_ASAP7_75t_R hold1184 (.A(net2729),
    .Y(net3308));
 BUFx2_ASAP7_75t_R hold1185 (.A(net3218),
    .Y(net3309));
 BUFx2_ASAP7_75t_R hold1186 (.A(net13),
    .Y(net3310));
 BUFx2_ASAP7_75t_R hold1187 (.A(net3219),
    .Y(net3311));
 BUFx2_ASAP7_75t_R hold1188 (.A(net2730),
    .Y(net3312));
 BUFx2_ASAP7_75t_R hold1189 (.A(boot_addr_i[16]),
    .Y(net3313));
 BUFx2_ASAP7_75t_R hold1190 (.A(net3040),
    .Y(net3314));
 BUFx2_ASAP7_75t_R hold1191 (.A(net2721),
    .Y(net3315));
 BUFx2_ASAP7_75t_R hold1192 (.A(net3041),
    .Y(net3316));
 BUFx2_ASAP7_75t_R hold1193 (.A(net7),
    .Y(net3317));
 BUFx2_ASAP7_75t_R hold1194 (.A(net3042),
    .Y(net3318));
 BUFx2_ASAP7_75t_R hold1195 (.A(net2722),
    .Y(net3319));
 BUFx2_ASAP7_75t_R hold1196 (.A(net3043),
    .Y(net3320));
 BUFx2_ASAP7_75t_R hold1197 (.A(boot_addr_i[27]),
    .Y(net3321));
 BUFx2_ASAP7_75t_R hold1198 (.A(net3143),
    .Y(net3322));
 BUFx2_ASAP7_75t_R hold1199 (.A(net2677),
    .Y(net3323));
 BUFx2_ASAP7_75t_R hold1200 (.A(net3144),
    .Y(net3324));
 BUFx2_ASAP7_75t_R hold1201 (.A(net18),
    .Y(net3325));
 BUFx2_ASAP7_75t_R hold1202 (.A(net3145),
    .Y(net3326));
 BUFx2_ASAP7_75t_R hold1203 (.A(net2678),
    .Y(net3327));
 BUFx2_ASAP7_75t_R hold1204 (.A(net3146),
    .Y(net3328));
 BUFx2_ASAP7_75t_R hold1205 (.A(boot_addr_i[18]),
    .Y(net3329));
 BUFx2_ASAP7_75t_R hold1206 (.A(net3230),
    .Y(net3330));
 BUFx2_ASAP7_75t_R hold1207 (.A(net2701),
    .Y(net3331));
 BUFx2_ASAP7_75t_R hold1208 (.A(net3231),
    .Y(net3332));
 BUFx2_ASAP7_75t_R hold1209 (.A(net9),
    .Y(net3333));
 BUFx2_ASAP7_75t_R hold1210 (.A(net3232),
    .Y(net3334));
 BUFx2_ASAP7_75t_R hold1211 (.A(net2702),
    .Y(net3335));
 BUFx2_ASAP7_75t_R hold1212 (.A(net3233),
    .Y(net3336));
 BUFx2_ASAP7_75t_R hold1213 (.A(boot_addr_i[21]),
    .Y(net3337));
 BUFx2_ASAP7_75t_R hold1214 (.A(net3011),
    .Y(net3338));
 BUFx2_ASAP7_75t_R hold1215 (.A(net2703),
    .Y(net3339));
 BUFx2_ASAP7_75t_R hold1216 (.A(net3012),
    .Y(net3340));
 BUFx2_ASAP7_75t_R hold1217 (.A(net12),
    .Y(net3341));
 BUFx2_ASAP7_75t_R hold1218 (.A(net3013),
    .Y(net3342));
 BUFx2_ASAP7_75t_R hold1219 (.A(net2704),
    .Y(net3343));
 BUFx2_ASAP7_75t_R hold1220 (.A(net3014),
    .Y(net3344));
 BUFx2_ASAP7_75t_R hold1221 (.A(boot_addr_i[26]),
    .Y(net3345));
 BUFx2_ASAP7_75t_R hold1222 (.A(net3234),
    .Y(net3346));
 BUFx2_ASAP7_75t_R hold1223 (.A(net2697),
    .Y(net3347));
 BUFx2_ASAP7_75t_R hold1224 (.A(net3235),
    .Y(net3348));
 BUFx2_ASAP7_75t_R hold1225 (.A(net17),
    .Y(net3349));
 BUFx2_ASAP7_75t_R hold1226 (.A(net3236),
    .Y(net3350));
 BUFx2_ASAP7_75t_R hold1227 (.A(net2698),
    .Y(net3351));
 BUFx2_ASAP7_75t_R hold1228 (.A(net3237),
    .Y(net3352));
 BUFx2_ASAP7_75t_R hold1229 (.A(net3484),
    .Y(net3353));
 BUFx2_ASAP7_75t_R hold1230 (.A(net3486),
    .Y(net3354));
 BUFx2_ASAP7_75t_R hold1231 (.A(_06259_),
    .Y(net3355));
 BUFx2_ASAP7_75t_R hold1232 (.A(net3410),
    .Y(net3356));
 BUFx2_ASAP7_75t_R hold1233 (.A(_06270_),
    .Y(net3357));
 BUFx2_ASAP7_75t_R hold1234 (.A(net3210),
    .Y(net3358));
 BUFx2_ASAP7_75t_R hold1235 (.A(boot_addr_i[25]),
    .Y(net3359));
 BUFx2_ASAP7_75t_R hold1236 (.A(net3153),
    .Y(net3360));
 BUFx2_ASAP7_75t_R hold1237 (.A(net2719),
    .Y(net3361));
 BUFx2_ASAP7_75t_R hold1238 (.A(net3154),
    .Y(net3362));
 BUFx2_ASAP7_75t_R hold1239 (.A(net16),
    .Y(net3363));
 BUFx2_ASAP7_75t_R hold1240 (.A(net3155),
    .Y(net3364));
 BUFx2_ASAP7_75t_R hold1241 (.A(net2720),
    .Y(net3365));
 BUFx2_ASAP7_75t_R hold1242 (.A(net3156),
    .Y(net3366));
 BUFx2_ASAP7_75t_R hold1243 (.A(net3624),
    .Y(net3367));
 BUFx2_ASAP7_75t_R hold1244 (.A(net129),
    .Y(net3368));
 BUFx2_ASAP7_75t_R hold1245 (.A(_06265_),
    .Y(net3369));
 BUFx2_ASAP7_75t_R hold1246 (.A(_06266_),
    .Y(net3370));
 BUFx2_ASAP7_75t_R hold1247 (.A(net3548),
    .Y(net3371));
 BUFx2_ASAP7_75t_R hold1248 (.A(net133),
    .Y(net3372));
 BUFx2_ASAP7_75t_R hold1249 (.A(net3550),
    .Y(net3373));
 BUFx2_ASAP7_75t_R hold1250 (.A(_06337_),
    .Y(net3374));
 BUFx2_ASAP7_75t_R hold1251 (.A(net3501),
    .Y(net3375));
 BUFx2_ASAP7_75t_R hold1252 (.A(net3381),
    .Y(net3376));
 BUFx2_ASAP7_75t_R hold1253 (.A(net3383),
    .Y(net3377));
 BUFx2_ASAP7_75t_R hold1254 (.A(_09485_),
    .Y(net3378));
 BUFx2_ASAP7_75t_R hold1255 (.A(_09486_),
    .Y(net3379));
 BUFx2_ASAP7_75t_R hold1256 (.A(_04096_),
    .Y(net3380));
 BUFx2_ASAP7_75t_R hold1257 (.A(hart_id_i[4]),
    .Y(net3381));
 BUFx2_ASAP7_75t_R hold1258 (.A(net3376),
    .Y(net3382));
 BUFx2_ASAP7_75t_R hold1259 (.A(net88),
    .Y(net3383));
 BUFx2_ASAP7_75t_R hold1260 (.A(net3377),
    .Y(net3384));
 BUFx2_ASAP7_75t_R hold1261 (.A(_07598_),
    .Y(net3385));
 BUFx2_ASAP7_75t_R hold1262 (.A(net3623),
    .Y(net3386));
 BUFx2_ASAP7_75t_R hold1263 (.A(net134),
    .Y(net3387));
 BUFx2_ASAP7_75t_R hold1264 (.A(_06292_),
    .Y(net3388));
 BUFx2_ASAP7_75t_R hold1265 (.A(net3488),
    .Y(net3389));
 BUFx2_ASAP7_75t_R hold1266 (.A(net3490),
    .Y(net3390));
 BUFx2_ASAP7_75t_R hold1267 (.A(_06312_),
    .Y(net3391));
 BUFx2_ASAP7_75t_R hold1268 (.A(boot_addr_i[29]),
    .Y(net3392));
 BUFx2_ASAP7_75t_R hold1269 (.A(net3186),
    .Y(net3393));
 BUFx2_ASAP7_75t_R hold1270 (.A(net2749),
    .Y(net3394));
 BUFx2_ASAP7_75t_R hold1271 (.A(net3187),
    .Y(net3395));
 BUFx2_ASAP7_75t_R hold1272 (.A(net20),
    .Y(net3396));
 BUFx2_ASAP7_75t_R hold1273 (.A(net3188),
    .Y(net3397));
 BUFx2_ASAP7_75t_R hold1274 (.A(net2750),
    .Y(net3398));
 BUFx2_ASAP7_75t_R hold1275 (.A(boot_addr_i[23]),
    .Y(net3399));
 BUFx2_ASAP7_75t_R hold1276 (.A(net3212),
    .Y(net3400));
 BUFx2_ASAP7_75t_R hold1277 (.A(net2745),
    .Y(net3401));
 BUFx2_ASAP7_75t_R hold1278 (.A(net3213),
    .Y(net3402));
 BUFx2_ASAP7_75t_R hold1279 (.A(net14),
    .Y(net3403));
 BUFx2_ASAP7_75t_R hold1280 (.A(net3214),
    .Y(net3404));
 BUFx2_ASAP7_75t_R hold1281 (.A(net2746),
    .Y(net3405));
 BUFx2_ASAP7_75t_R hold1282 (.A(irq_fast_i[10]),
    .Y(net3406));
 BUFx2_ASAP7_75t_R hold1283 (.A(net131),
    .Y(net3407));
 BUFx2_ASAP7_75t_R hold1284 (.A(_06253_),
    .Y(net3408));
 BUFx2_ASAP7_75t_R hold1285 (.A(_06254_),
    .Y(net3409));
 BUFx2_ASAP7_75t_R hold1286 (.A(_06263_),
    .Y(net3410));
 BUFx2_ASAP7_75t_R hold1287 (.A(net3356),
    .Y(net3411));
 BUFx2_ASAP7_75t_R hold1288 (.A(_06358_),
    .Y(net3412));
 BUFx2_ASAP7_75t_R hold1289 (.A(_06359_),
    .Y(net3413));
 BUFx2_ASAP7_75t_R hold1290 (.A(_12393_),
    .Y(net3414));
 BUFx2_ASAP7_75t_R hold1291 (.A(boot_addr_i[8]),
    .Y(net3415));
 BUFx2_ASAP7_75t_R hold1292 (.A(net3086),
    .Y(net3416));
 BUFx2_ASAP7_75t_R hold1293 (.A(net2709),
    .Y(net3417));
 BUFx2_ASAP7_75t_R hold1294 (.A(net3087),
    .Y(net3418));
 BUFx2_ASAP7_75t_R hold1295 (.A(net23),
    .Y(net3419));
 BUFx2_ASAP7_75t_R hold1296 (.A(net3088),
    .Y(net3420));
 BUFx2_ASAP7_75t_R hold1297 (.A(net2710),
    .Y(net3421));
 BUFx2_ASAP7_75t_R hold1298 (.A(net3089),
    .Y(net3422));
 BUFx2_ASAP7_75t_R hold1299 (.A(boot_addr_i[19]),
    .Y(net3423));
 BUFx2_ASAP7_75t_R hold1300 (.A(net3169),
    .Y(net3424));
 BUFx2_ASAP7_75t_R hold1301 (.A(net2673),
    .Y(net3425));
 BUFx2_ASAP7_75t_R hold1302 (.A(net3170),
    .Y(net3426));
 BUFx2_ASAP7_75t_R hold1303 (.A(net10),
    .Y(net3427));
 BUFx2_ASAP7_75t_R hold1304 (.A(net3171),
    .Y(net3428));
 BUFx2_ASAP7_75t_R hold1305 (.A(net2674),
    .Y(net3429));
 BUFx2_ASAP7_75t_R hold1306 (.A(net3172),
    .Y(net3430));
 BUFx2_ASAP7_75t_R hold1307 (.A(boot_addr_i[9]),
    .Y(net3431));
 BUFx2_ASAP7_75t_R hold1308 (.A(net3123),
    .Y(net3432));
 BUFx2_ASAP7_75t_R hold1309 (.A(net2751),
    .Y(net3433));
 BUFx2_ASAP7_75t_R hold1310 (.A(net3124),
    .Y(net3434));
 BUFx2_ASAP7_75t_R hold1311 (.A(net24),
    .Y(net3435));
 BUFx2_ASAP7_75t_R hold1312 (.A(net3125),
    .Y(net3436));
 BUFx2_ASAP7_75t_R hold1313 (.A(net2752),
    .Y(net3437));
 BUFx2_ASAP7_75t_R hold1314 (.A(boot_addr_i[24]),
    .Y(net3438));
 BUFx2_ASAP7_75t_R hold1315 (.A(net3174),
    .Y(net3439));
 BUFx2_ASAP7_75t_R hold1316 (.A(net2747),
    .Y(net3440));
 BUFx2_ASAP7_75t_R hold1317 (.A(net3175),
    .Y(net3441));
 BUFx2_ASAP7_75t_R hold1318 (.A(net15),
    .Y(net3442));
 BUFx2_ASAP7_75t_R hold1319 (.A(net3176),
    .Y(net3443));
 BUFx2_ASAP7_75t_R hold1320 (.A(net2748),
    .Y(net3444));
 BUFx2_ASAP7_75t_R hold1321 (.A(boot_addr_i[15]),
    .Y(net3445));
 BUFx2_ASAP7_75t_R hold1322 (.A(net3191),
    .Y(net3446));
 BUFx2_ASAP7_75t_R hold1323 (.A(net2711),
    .Y(net3447));
 BUFx2_ASAP7_75t_R hold1324 (.A(net3192),
    .Y(net3448));
 BUFx2_ASAP7_75t_R hold1325 (.A(net6),
    .Y(net3449));
 BUFx2_ASAP7_75t_R hold1326 (.A(net3193),
    .Y(net3450));
 BUFx2_ASAP7_75t_R hold1327 (.A(net2712),
    .Y(net3451));
 BUFx2_ASAP7_75t_R hold1328 (.A(net3194),
    .Y(net3452));
 BUFx2_ASAP7_75t_R hold1329 (.A(boot_addr_i[12]),
    .Y(net3453));
 BUFx2_ASAP7_75t_R hold1330 (.A(net3158),
    .Y(net3454));
 BUFx2_ASAP7_75t_R hold1331 (.A(net2699),
    .Y(net3455));
 BUFx2_ASAP7_75t_R hold1332 (.A(net3159),
    .Y(net3456));
 BUFx2_ASAP7_75t_R hold1333 (.A(net3),
    .Y(net3457));
 BUFx2_ASAP7_75t_R hold1334 (.A(net3160),
    .Y(net3458));
 BUFx2_ASAP7_75t_R hold1335 (.A(net2700),
    .Y(net3459));
 BUFx2_ASAP7_75t_R hold1336 (.A(net3161),
    .Y(net3460));
 BUFx2_ASAP7_75t_R hold1337 (.A(boot_addr_i[17]),
    .Y(net3461));
 BUFx2_ASAP7_75t_R hold1338 (.A(net3196),
    .Y(net3462));
 BUFx2_ASAP7_75t_R hold1339 (.A(net2725),
    .Y(net3463));
 BUFx2_ASAP7_75t_R hold1340 (.A(net3197),
    .Y(net3464));
 BUFx2_ASAP7_75t_R hold1341 (.A(net8),
    .Y(net3465));
 BUFx2_ASAP7_75t_R hold1342 (.A(net3198),
    .Y(net3466));
 BUFx2_ASAP7_75t_R hold1343 (.A(net2726),
    .Y(net3467));
 BUFx2_ASAP7_75t_R hold1344 (.A(boot_addr_i[14]),
    .Y(net3468));
 BUFx2_ASAP7_75t_R hold1345 (.A(net3163),
    .Y(net3469));
 BUFx2_ASAP7_75t_R hold1346 (.A(net2683),
    .Y(net3470));
 BUFx2_ASAP7_75t_R hold1347 (.A(net3164),
    .Y(net3471));
 BUFx2_ASAP7_75t_R hold1348 (.A(net5),
    .Y(net3472));
 BUFx2_ASAP7_75t_R hold1349 (.A(net3165),
    .Y(net3473));
 BUFx2_ASAP7_75t_R hold1350 (.A(net2684),
    .Y(net3474));
 BUFx2_ASAP7_75t_R hold1351 (.A(net3166),
    .Y(net3475));
 BUFx2_ASAP7_75t_R hold1352 (.A(net3662),
    .Y(net3476));
 BUFx2_ASAP7_75t_R hold1353 (.A(net144),
    .Y(net3477));
 BUFx2_ASAP7_75t_R hold1354 (.A(_06257_),
    .Y(net3478));
 BUFx2_ASAP7_75t_R hold1355 (.A(_06334_),
    .Y(net3479));
 BUFx2_ASAP7_75t_R hold1356 (.A(_06347_),
    .Y(net3480));
 BUFx2_ASAP7_75t_R hold1357 (.A(_06349_),
    .Y(net3481));
 BUFx2_ASAP7_75t_R hold1358 (.A(_06350_),
    .Y(net3482));
 BUFx2_ASAP7_75t_R hold1359 (.A(_06351_),
    .Y(net3483));
 BUFx2_ASAP7_75t_R hold1360 (.A(irq_fast_i[14]),
    .Y(net3484));
 BUFx2_ASAP7_75t_R hold1361 (.A(net3353),
    .Y(net3485));
 BUFx2_ASAP7_75t_R hold1362 (.A(net135),
    .Y(net3486));
 BUFx2_ASAP7_75t_R hold1363 (.A(net3354),
    .Y(net3487));
 BUFx2_ASAP7_75t_R hold1364 (.A(_06294_),
    .Y(net3488));
 BUFx2_ASAP7_75t_R hold1365 (.A(net3389),
    .Y(net3489));
 BUFx2_ASAP7_75t_R hold1366 (.A(_06295_),
    .Y(net3490));
 BUFx2_ASAP7_75t_R hold1367 (.A(net3600),
    .Y(net3491));
 BUFx2_ASAP7_75t_R hold1368 (.A(net142),
    .Y(net3492));
 BUFx2_ASAP7_75t_R hold1369 (.A(_06241_),
    .Y(net3493));
 BUFx2_ASAP7_75t_R hold1370 (.A(_06251_),
    .Y(net3494));
 BUFx2_ASAP7_75t_R hold1371 (.A(net3301),
    .Y(net3495));
 BUFx2_ASAP7_75t_R hold1372 (.A(net3685),
    .Y(net3496));
 BUFx2_ASAP7_75t_R hold1373 (.A(net139),
    .Y(net3497));
 BUFx2_ASAP7_75t_R hold1374 (.A(_06244_),
    .Y(net3498));
 BUFx2_ASAP7_75t_R hold1375 (.A(_06335_),
    .Y(net3499));
 BUFx2_ASAP7_75t_R hold1376 (.A(_06336_),
    .Y(net3500));
 BUFx2_ASAP7_75t_R hold1377 (.A(net3514),
    .Y(net3501));
 BUFx2_ASAP7_75t_R hold1378 (.A(net3375),
    .Y(net3502));
 BUFx2_ASAP7_75t_R hold1379 (.A(_06343_),
    .Y(net3503));
 BUFx2_ASAP7_75t_R hold1380 (.A(net3537),
    .Y(net3504));
 BUFx2_ASAP7_75t_R hold1381 (.A(net132),
    .Y(net3505));
 BUFx2_ASAP7_75t_R hold1382 (.A(_06252_),
    .Y(net3506));
 BUFx2_ASAP7_75t_R hold1383 (.A(_06323_),
    .Y(net3507));
 BUFx2_ASAP7_75t_R hold1384 (.A(net3551),
    .Y(net3508));
 BUFx2_ASAP7_75t_R hold1385 (.A(_06327_),
    .Y(net3509));
 BUFx2_ASAP7_75t_R hold1386 (.A(_06328_),
    .Y(net3510));
 BUFx2_ASAP7_75t_R hold1387 (.A(_06330_),
    .Y(net3511));
 BUFx2_ASAP7_75t_R hold1388 (.A(net3564),
    .Y(net3512));
 BUFx2_ASAP7_75t_R hold1389 (.A(net146),
    .Y(net3513));
 BUFx2_ASAP7_75t_R hold1390 (.A(_06338_),
    .Y(net3514));
 BUFx2_ASAP7_75t_R hold1391 (.A(net3626),
    .Y(net3515));
 BUFx2_ASAP7_75t_R hold1392 (.A(net3628),
    .Y(net3516));
 BUFx2_ASAP7_75t_R hold1393 (.A(_11069_),
    .Y(net3517));
 BUFx2_ASAP7_75t_R hold1394 (.A(_12374_),
    .Y(net3518));
 BUFx2_ASAP7_75t_R hold1395 (.A(_04301_),
    .Y(net3519));
 BUFx2_ASAP7_75t_R hold1396 (.A(net3546),
    .Y(net3520));
 BUFx2_ASAP7_75t_R hold1397 (.A(net143),
    .Y(net3521));
 BUFx2_ASAP7_75t_R hold1398 (.A(net3534),
    .Y(net3522));
 BUFx2_ASAP7_75t_R hold1399 (.A(net3536),
    .Y(net3523));
 BUFx2_ASAP7_75t_R hold1400 (.A(_07444_),
    .Y(net3524));
 BUFx2_ASAP7_75t_R hold1401 (.A(_07462_),
    .Y(net3525));
 BUFx2_ASAP7_75t_R hold1402 (.A(_09472_),
    .Y(net3526));
 BUFx2_ASAP7_75t_R hold1403 (.A(_09473_),
    .Y(net3527));
 BUFx2_ASAP7_75t_R hold1404 (.A(_02866_),
    .Y(net3528));
 BUFx2_ASAP7_75t_R hold1405 (.A(net3587),
    .Y(net3529));
 BUFx2_ASAP7_75t_R hold1406 (.A(net3589),
    .Y(net3530));
 BUFx2_ASAP7_75t_R hold1407 (.A(_09643_),
    .Y(net3531));
 BUFx2_ASAP7_75t_R hold1408 (.A(irq_fast_i[5]),
    .Y(net3532));
 BUFx2_ASAP7_75t_R hold1409 (.A(net140),
    .Y(net3533));
 BUFx2_ASAP7_75t_R hold1410 (.A(hart_id_i[2]),
    .Y(net3534));
 BUFx2_ASAP7_75t_R hold1411 (.A(net3522),
    .Y(net3535));
 BUFx2_ASAP7_75t_R hold1412 (.A(net84),
    .Y(net3536));
 BUFx2_ASAP7_75t_R hold1413 (.A(irq_fast_i[11]),
    .Y(net3537));
 BUFx2_ASAP7_75t_R hold1414 (.A(net3504),
    .Y(net3538));
 BUFx2_ASAP7_75t_R hold1415 (.A(net3583),
    .Y(net3539));
 BUFx2_ASAP7_75t_R hold1416 (.A(net3585),
    .Y(net3540));
 BUFx2_ASAP7_75t_R hold1417 (.A(_09566_),
    .Y(net3541));
 BUFx2_ASAP7_75t_R hold1418 (.A(net3559),
    .Y(net3542));
 BUFx2_ASAP7_75t_R hold1419 (.A(net3561),
    .Y(net3543));
 BUFx2_ASAP7_75t_R hold1420 (.A(_09477_),
    .Y(net3544));
 BUFx2_ASAP7_75t_R hold1421 (.A(_04268_),
    .Y(net3545));
 BUFx2_ASAP7_75t_R hold1422 (.A(irq_fast_i[8]),
    .Y(net3546));
 BUFx2_ASAP7_75t_R hold1423 (.A(net3520),
    .Y(net3547));
 BUFx2_ASAP7_75t_R hold1424 (.A(irq_fast_i[12]),
    .Y(net3548));
 BUFx2_ASAP7_75t_R hold1425 (.A(net3371),
    .Y(net3549));
 BUFx2_ASAP7_75t_R hold1426 (.A(_06262_),
    .Y(net3550));
 BUFx2_ASAP7_75t_R hold1427 (.A(_06326_),
    .Y(net3551));
 BUFx2_ASAP7_75t_R hold1428 (.A(net3567),
    .Y(net3552));
 BUFx2_ASAP7_75t_R hold1429 (.A(net3569),
    .Y(net3553));
 BUFx2_ASAP7_75t_R hold1430 (.A(net3576),
    .Y(net3554));
 BUFx2_ASAP7_75t_R hold1431 (.A(net137),
    .Y(net3555));
 BUFx2_ASAP7_75t_R hold1432 (.A(_09600_),
    .Y(net3556));
 BUFx2_ASAP7_75t_R hold1433 (.A(net3572),
    .Y(net3557));
 BUFx2_ASAP7_75t_R hold1434 (.A(_04253_),
    .Y(net3558));
 BUFx2_ASAP7_75t_R hold1435 (.A(hart_id_i[3]),
    .Y(net3559));
 BUFx2_ASAP7_75t_R hold1436 (.A(net3542),
    .Y(net3560));
 BUFx2_ASAP7_75t_R hold1437 (.A(net87),
    .Y(net3561));
 BUFx2_ASAP7_75t_R hold1438 (.A(_07540_),
    .Y(net3562));
 BUFx2_ASAP7_75t_R hold1439 (.A(net3544),
    .Y(net3563));
 BUFx2_ASAP7_75t_R hold1440 (.A(irq_software_i),
    .Y(net3564));
 BUFx2_ASAP7_75t_R hold1441 (.A(net3692),
    .Y(net3565));
 BUFx2_ASAP7_75t_R hold1442 (.A(net141),
    .Y(net3566));
 BUFx2_ASAP7_75t_R hold1443 (.A(hart_id_i[18]),
    .Y(net3567));
 BUFx2_ASAP7_75t_R hold1444 (.A(net3552),
    .Y(net3568));
 BUFx2_ASAP7_75t_R hold1445 (.A(net71),
    .Y(net3569));
 BUFx2_ASAP7_75t_R hold1446 (.A(net3553),
    .Y(net3570));
 BUFx2_ASAP7_75t_R hold1447 (.A(net3556),
    .Y(net3571));
 BUFx2_ASAP7_75t_R hold1448 (.A(_09601_),
    .Y(net3572));
 BUFx2_ASAP7_75t_R hold1449 (.A(net3557),
    .Y(net3573));
 BUFx2_ASAP7_75t_R hold1450 (.A(hart_id_i[31]),
    .Y(net3574));
 BUFx2_ASAP7_75t_R hold1451 (.A(net86),
    .Y(net3575));
 BUFx2_ASAP7_75t_R hold1452 (.A(irq_fast_i[2]),
    .Y(net3576));
 BUFx2_ASAP7_75t_R hold1453 (.A(net3554),
    .Y(net3577));
 BUFx2_ASAP7_75t_R hold1454 (.A(net3596),
    .Y(net3578));
 BUFx2_ASAP7_75t_R hold1455 (.A(net3598),
    .Y(net3579));
 BUFx2_ASAP7_75t_R hold1456 (.A(_09637_),
    .Y(net3580));
 BUFx2_ASAP7_75t_R hold1457 (.A(_12112_),
    .Y(net3581));
 BUFx2_ASAP7_75t_R hold1458 (.A(_04208_),
    .Y(net3582));
 BUFx2_ASAP7_75t_R hold1459 (.A(hart_id_i[14]),
    .Y(net3583));
 BUFx2_ASAP7_75t_R hold1460 (.A(net3539),
    .Y(net3584));
 BUFx2_ASAP7_75t_R hold1461 (.A(net67),
    .Y(net3585));
 BUFx2_ASAP7_75t_R hold1462 (.A(net3540),
    .Y(net3586));
 BUFx2_ASAP7_75t_R hold1463 (.A(hart_id_i[24]),
    .Y(net3587));
 BUFx2_ASAP7_75t_R hold1464 (.A(net3529),
    .Y(net3588));
 BUFx2_ASAP7_75t_R hold1465 (.A(net78),
    .Y(net3589));
 BUFx2_ASAP7_75t_R hold1466 (.A(net3530),
    .Y(net3590));
 BUFx2_ASAP7_75t_R hold1467 (.A(net3616),
    .Y(net3591));
 BUFx2_ASAP7_75t_R hold1468 (.A(net3618),
    .Y(net3592));
 BUFx2_ASAP7_75t_R hold1469 (.A(_08531_),
    .Y(net3593));
 BUFx2_ASAP7_75t_R hold1470 (.A(_09668_),
    .Y(net3594));
 BUFx2_ASAP7_75t_R hold1471 (.A(_04262_),
    .Y(net3595));
 BUFx2_ASAP7_75t_R hold1472 (.A(hart_id_i[23]),
    .Y(net3596));
 BUFx2_ASAP7_75t_R hold1473 (.A(net3578),
    .Y(net3597));
 BUFx2_ASAP7_75t_R hold1474 (.A(net77),
    .Y(net3598));
 BUFx2_ASAP7_75t_R hold1475 (.A(net3580),
    .Y(net3599));
 BUFx2_ASAP7_75t_R hold1476 (.A(irq_fast_i[7]),
    .Y(net3600));
 BUFx2_ASAP7_75t_R hold1477 (.A(net3619),
    .Y(net3601));
 BUFx2_ASAP7_75t_R hold1478 (.A(net3621),
    .Y(net3602));
 BUFx2_ASAP7_75t_R hold1479 (.A(_08138_),
    .Y(net3603));
 BUFx2_ASAP7_75t_R hold1480 (.A(net3622),
    .Y(net3604));
 BUFx2_ASAP7_75t_R hold1481 (.A(_04251_),
    .Y(net3605));
 BUFx2_ASAP7_75t_R hold1482 (.A(hart_id_i[29]),
    .Y(net3606));
 BUFx2_ASAP7_75t_R hold1483 (.A(net83),
    .Y(net3607));
 BUFx2_ASAP7_75t_R hold1484 (.A(_08586_),
    .Y(net3608));
 BUFx2_ASAP7_75t_R hold1485 (.A(_08587_),
    .Y(net3609));
 BUFx2_ASAP7_75t_R hold1486 (.A(_08588_),
    .Y(net3610));
 BUFx2_ASAP7_75t_R hold1487 (.A(_09683_),
    .Y(net3611));
 BUFx2_ASAP7_75t_R hold1488 (.A(net3651),
    .Y(net3612));
 BUFx2_ASAP7_75t_R hold1489 (.A(net3653),
    .Y(net3613));
 BUFx2_ASAP7_75t_R hold1490 (.A(_07742_),
    .Y(net3614));
 BUFx2_ASAP7_75t_R hold1491 (.A(_09512_),
    .Y(net3615));
 BUFx2_ASAP7_75t_R hold1492 (.A(hart_id_i[27]),
    .Y(net3616));
 BUFx2_ASAP7_75t_R hold1493 (.A(net3591),
    .Y(net3617));
 BUFx2_ASAP7_75t_R hold1494 (.A(net81),
    .Y(net3618));
 BUFx2_ASAP7_75t_R hold1495 (.A(hart_id_i[16]),
    .Y(net3619));
 BUFx2_ASAP7_75t_R hold1496 (.A(net3601),
    .Y(net3620));
 BUFx2_ASAP7_75t_R hold1497 (.A(net69),
    .Y(net3621));
 BUFx2_ASAP7_75t_R hold1498 (.A(_09585_),
    .Y(net3622));
 BUFx2_ASAP7_75t_R hold1499 (.A(irq_fast_i[13]),
    .Y(net3623));
 BUFx2_ASAP7_75t_R hold1500 (.A(irq_external_i),
    .Y(net3624));
 BUFx2_ASAP7_75t_R hold1501 (.A(net3367),
    .Y(net3625));
 BUFx2_ASAP7_75t_R hold1502 (.A(hart_id_i[0]),
    .Y(net3626));
 BUFx2_ASAP7_75t_R hold1503 (.A(net3515),
    .Y(net3627));
 BUFx2_ASAP7_75t_R hold1504 (.A(net62),
    .Y(net3628));
 BUFx2_ASAP7_75t_R hold1505 (.A(net3634),
    .Y(net3629));
 BUFx2_ASAP7_75t_R hold1506 (.A(net89),
    .Y(net3630));
 BUFx2_ASAP7_75t_R hold1507 (.A(_07652_),
    .Y(net3631));
 BUFx2_ASAP7_75t_R hold1508 (.A(_09493_),
    .Y(net3632));
 BUFx2_ASAP7_75t_R hold1509 (.A(_02869_),
    .Y(net3633));
 BUFx2_ASAP7_75t_R hold1510 (.A(hart_id_i[5]),
    .Y(net3634));
 BUFx2_ASAP7_75t_R hold1511 (.A(net3629),
    .Y(net3635));
 BUFx2_ASAP7_75t_R hold1512 (.A(net3641),
    .Y(net3636));
 BUFx2_ASAP7_75t_R hold1513 (.A(net79),
    .Y(net3637));
 BUFx2_ASAP7_75t_R hold1514 (.A(_08471_),
    .Y(net3638));
 BUFx2_ASAP7_75t_R hold1515 (.A(net3643),
    .Y(net3639));
 BUFx2_ASAP7_75t_R hold1516 (.A(_04210_),
    .Y(net3640));
 BUFx2_ASAP7_75t_R hold1517 (.A(hart_id_i[25]),
    .Y(net3641));
 BUFx2_ASAP7_75t_R hold1518 (.A(net3636),
    .Y(net3642));
 BUFx2_ASAP7_75t_R hold1519 (.A(_09653_),
    .Y(net3643));
 BUFx2_ASAP7_75t_R hold1520 (.A(net3639),
    .Y(net3644));
 BUFx2_ASAP7_75t_R hold1521 (.A(net3649),
    .Y(net3645));
 BUFx2_ASAP7_75t_R hold1522 (.A(net73),
    .Y(net3646));
 BUFx2_ASAP7_75t_R hold1523 (.A(_09452_),
    .Y(net3647));
 BUFx2_ASAP7_75t_R hold1524 (.A(_04093_),
    .Y(net3648));
 BUFx2_ASAP7_75t_R hold1525 (.A(hart_id_i[1]),
    .Y(net3649));
 BUFx2_ASAP7_75t_R hold1526 (.A(net3645),
    .Y(net3650));
 BUFx2_ASAP7_75t_R hold1527 (.A(hart_id_i[7]),
    .Y(net3651));
 BUFx2_ASAP7_75t_R hold1528 (.A(net3612),
    .Y(net3652));
 BUFx2_ASAP7_75t_R hold1529 (.A(net91),
    .Y(net3653));
 BUFx2_ASAP7_75t_R hold1530 (.A(net3615),
    .Y(net3654));
 BUFx2_ASAP7_75t_R hold1531 (.A(_04267_),
    .Y(net3655));
 BUFx2_ASAP7_75t_R hold1532 (.A(irq_timer_i),
    .Y(net3656));
 BUFx2_ASAP7_75t_R hold1533 (.A(hart_id_i[17]),
    .Y(net3657));
 BUFx2_ASAP7_75t_R hold1534 (.A(net70),
    .Y(net3658));
 BUFx2_ASAP7_75t_R hold1535 (.A(_08168_),
    .Y(net3659));
 BUFx2_ASAP7_75t_R hold1536 (.A(net3668),
    .Y(net3660));
 BUFx2_ASAP7_75t_R hold1537 (.A(_04252_),
    .Y(net3661));
 BUFx2_ASAP7_75t_R hold1538 (.A(irq_fast_i[9]),
    .Y(net3662));
 BUFx2_ASAP7_75t_R hold1539 (.A(net3476),
    .Y(net3663));
 BUFx2_ASAP7_75t_R hold1540 (.A(irq_fast_i[1]),
    .Y(net3664));
 BUFx2_ASAP7_75t_R hold1541 (.A(net136),
    .Y(net3665));
 BUFx2_ASAP7_75t_R hold1542 (.A(_08170_),
    .Y(net3666));
 BUFx2_ASAP7_75t_R hold1543 (.A(_08173_),
    .Y(net3667));
 BUFx2_ASAP7_75t_R hold1544 (.A(_09592_),
    .Y(net3668));
 BUFx2_ASAP7_75t_R hold1545 (.A(irq_fast_i[0]),
    .Y(net3669));
 BUFx2_ASAP7_75t_R hold1546 (.A(net3693),
    .Y(net3670));
 BUFx2_ASAP7_75t_R hold1547 (.A(net65),
    .Y(net3671));
 BUFx2_ASAP7_75t_R hold1548 (.A(_07980_),
    .Y(net3672));
 BUFx2_ASAP7_75t_R hold1549 (.A(_09548_),
    .Y(net3673));
 BUFx2_ASAP7_75t_R hold1550 (.A(net3684),
    .Y(net3674));
 BUFx2_ASAP7_75t_R hold1551 (.A(net75),
    .Y(net3675));
 BUFx2_ASAP7_75t_R hold1552 (.A(_08317_),
    .Y(net3676));
 BUFx2_ASAP7_75t_R hold1553 (.A(_08319_),
    .Y(net3677));
 BUFx2_ASAP7_75t_R hold1554 (.A(_09623_),
    .Y(net3678));
 BUFx2_ASAP7_75t_R hold1555 (.A(hart_id_i[20]),
    .Y(net3679));
 BUFx2_ASAP7_75t_R hold1556 (.A(net74),
    .Y(net3680));
 BUFx2_ASAP7_75t_R hold1557 (.A(net3686),
    .Y(net3681));
 BUFx2_ASAP7_75t_R hold1558 (.A(_09615_),
    .Y(net3682));
 BUFx2_ASAP7_75t_R hold1559 (.A(_09616_),
    .Y(net3683));
 BUFx2_ASAP7_75t_R hold1560 (.A(hart_id_i[21]),
    .Y(net3684));
 BUFx2_ASAP7_75t_R hold1561 (.A(irq_fast_i[4]),
    .Y(net3685));
 BUFx2_ASAP7_75t_R hold1562 (.A(_08285_),
    .Y(net3686));
 BUFx2_ASAP7_75t_R hold1563 (.A(hart_id_i[22]),
    .Y(net3687));
 BUFx2_ASAP7_75t_R hold1564 (.A(net76),
    .Y(net3688));
 BUFx2_ASAP7_75t_R hold1565 (.A(_08356_),
    .Y(net3689));
 BUFx2_ASAP7_75t_R hold1566 (.A(_08358_),
    .Y(net3690));
 BUFx2_ASAP7_75t_R hold1567 (.A(_09631_),
    .Y(net3691));
 BUFx2_ASAP7_75t_R hold1568 (.A(irq_fast_i[6]),
    .Y(net3692));
 BUFx2_ASAP7_75t_R hold1569 (.A(hart_id_i[12]),
    .Y(net3693));
 BUFx2_ASAP7_75t_R hold1570 (.A(net3699),
    .Y(net3694));
 BUFx2_ASAP7_75t_R hold1571 (.A(net85),
    .Y(net3695));
 BUFx2_ASAP7_75t_R hold1572 (.A(_08599_),
    .Y(net3696));
 BUFx2_ASAP7_75t_R hold1573 (.A(_08607_),
    .Y(net3697));
 BUFx2_ASAP7_75t_R hold1574 (.A(_09691_),
    .Y(net3698));
 BUFx2_ASAP7_75t_R hold1575 (.A(hart_id_i[30]),
    .Y(net3699));
 BUFx2_ASAP7_75t_R hold1576 (.A(hart_id_i[11]),
    .Y(net3700));
 BUFx2_ASAP7_75t_R hold1577 (.A(net64),
    .Y(net3701));
 BUFx2_ASAP7_75t_R hold1578 (.A(_07933_),
    .Y(net3702));
 BUFx2_ASAP7_75t_R hold1579 (.A(net3748),
    .Y(net3703));
 BUFx2_ASAP7_75t_R hold1580 (.A(net138),
    .Y(net3704));
 BUFx2_ASAP7_75t_R hold1581 (.A(net3730),
    .Y(net3705));
 BUFx2_ASAP7_75t_R hold1582 (.A(net3732),
    .Y(net3706));
 BUFx2_ASAP7_75t_R hold1583 (.A(_09556_),
    .Y(net3707));
 BUFx2_ASAP7_75t_R hold1584 (.A(_11835_),
    .Y(net3708));
 BUFx2_ASAP7_75t_R hold1585 (.A(net3717),
    .Y(net3709));
 BUFx2_ASAP7_75t_R hold1586 (.A(net3719),
    .Y(net3710));
 BUFx2_ASAP7_75t_R hold1587 (.A(_09607_),
    .Y(net3711));
 BUFx2_ASAP7_75t_R hold1588 (.A(_04254_),
    .Y(net3712));
 BUFx2_ASAP7_75t_R hold1589 (.A(net3737),
    .Y(net3713));
 BUFx2_ASAP7_75t_R hold1590 (.A(net93),
    .Y(net3714));
 BUFx2_ASAP7_75t_R hold1591 (.A(_07851_),
    .Y(net3715));
 BUFx2_ASAP7_75t_R hold1592 (.A(_09524_),
    .Y(net3716));
 BUFx2_ASAP7_75t_R hold1593 (.A(hart_id_i[19]),
    .Y(net3717));
 BUFx2_ASAP7_75t_R hold1594 (.A(net3709),
    .Y(net3718));
 BUFx2_ASAP7_75t_R hold1595 (.A(net72),
    .Y(net3719));
 BUFx2_ASAP7_75t_R hold1596 (.A(_08256_),
    .Y(net3720));
 BUFx2_ASAP7_75t_R hold1597 (.A(net3711),
    .Y(net3721));
 BUFx2_ASAP7_75t_R hold1598 (.A(net3738),
    .Y(net3722));
 BUFx2_ASAP7_75t_R hold1599 (.A(net92),
    .Y(net3723));
 BUFx2_ASAP7_75t_R hold1600 (.A(_07795_),
    .Y(net3724));
 BUFx2_ASAP7_75t_R hold1601 (.A(_09518_),
    .Y(net3725));
 BUFx2_ASAP7_75t_R hold1602 (.A(data_err_i),
    .Y(net3726));
 BUFx2_ASAP7_75t_R hold1603 (.A(net3033),
    .Y(net3727));
 BUFx2_ASAP7_75t_R hold1604 (.A(net2731),
    .Y(net3728));
 BUFx2_ASAP7_75t_R hold1605 (.A(net3034),
    .Y(net3729));
 BUFx2_ASAP7_75t_R hold1606 (.A(hart_id_i[13]),
    .Y(net3730));
 BUFx2_ASAP7_75t_R hold1607 (.A(net3705),
    .Y(net3731));
 BUFx2_ASAP7_75t_R hold1608 (.A(net66),
    .Y(net3732));
 BUFx2_ASAP7_75t_R hold1609 (.A(hart_id_i[10]),
    .Y(net3733));
 BUFx2_ASAP7_75t_R hold1610 (.A(net63),
    .Y(net3734));
 BUFx2_ASAP7_75t_R hold1611 (.A(_07882_),
    .Y(net3735));
 BUFx2_ASAP7_75t_R hold1612 (.A(_09531_),
    .Y(net3736));
 BUFx2_ASAP7_75t_R hold1613 (.A(hart_id_i[9]),
    .Y(net3737));
 BUFx2_ASAP7_75t_R hold1614 (.A(hart_id_i[8]),
    .Y(net3738));
 BUFx2_ASAP7_75t_R hold1615 (.A(hart_id_i[28]),
    .Y(net3739));
 BUFx2_ASAP7_75t_R hold1616 (.A(net82),
    .Y(net3740));
 BUFx2_ASAP7_75t_R hold1617 (.A(_08556_),
    .Y(net3741));
 BUFx2_ASAP7_75t_R hold1618 (.A(_08558_),
    .Y(net3742));
 BUFx2_ASAP7_75t_R hold1619 (.A(hart_id_i[6]),
    .Y(net3743));
 BUFx2_ASAP7_75t_R hold1620 (.A(net90),
    .Y(net3744));
 BUFx2_ASAP7_75t_R hold1621 (.A(net3766),
    .Y(net3745));
 BUFx2_ASAP7_75t_R hold1622 (.A(net68),
    .Y(net3746));
 BUFx2_ASAP7_75t_R hold1623 (.A(_09575_),
    .Y(net3747));
 BUFx2_ASAP7_75t_R hold1624 (.A(irq_fast_i[3]),
    .Y(net3748));
 BUFx2_ASAP7_75t_R hold1625 (.A(hart_id_i[26]),
    .Y(net3749));
 BUFx2_ASAP7_75t_R hold1626 (.A(net80),
    .Y(net3750));
 BUFx2_ASAP7_75t_R hold1627 (.A(_08497_),
    .Y(net3751));
 BUFx2_ASAP7_75t_R hold1628 (.A(_08503_),
    .Y(net3752));
 BUFx2_ASAP7_75t_R hold1629 (.A(irq_nm_i),
    .Y(net3753));
 BUFx2_ASAP7_75t_R hold1630 (.A(net3128),
    .Y(net3754));
 BUFx2_ASAP7_75t_R hold1631 (.A(net2642),
    .Y(net3755));
 BUFx2_ASAP7_75t_R hold1632 (.A(net3129),
    .Y(net3756));
 BUFx2_ASAP7_75t_R hold1633 (.A(net145),
    .Y(net3757));
 BUFx2_ASAP7_75t_R hold1634 (.A(net3130),
    .Y(net3758));
 BUFx2_ASAP7_75t_R hold1635 (.A(net3929),
    .Y(net3759));
 BUFx2_ASAP7_75t_R hold1636 (.A(net3931),
    .Y(net3760));
 BUFx2_ASAP7_75t_R hold1637 (.A(net3933),
    .Y(net3761));
 BUFx2_ASAP7_75t_R hold1638 (.A(net3765),
    .Y(net3762));
 BUFx2_ASAP7_75t_R hold1639 (.A(net56),
    .Y(net3763));
 BUFx2_ASAP7_75t_R hold1640 (.A(_07758_),
    .Y(net3764));
 BUFx2_ASAP7_75t_R hold1641 (.A(data_rdata_i[7]),
    .Y(net3765));
 BUFx2_ASAP7_75t_R hold1642 (.A(hart_id_i[15]),
    .Y(net3766));
 BUFx2_ASAP7_75t_R hold1643 (.A(net3745),
    .Y(net3767));
 BUFx2_ASAP7_75t_R hold1644 (.A(data_rdata_i[6]),
    .Y(net3768));
 BUFx2_ASAP7_75t_R hold1645 (.A(net55),
    .Y(net3769));
 BUFx2_ASAP7_75t_R hold1646 (.A(_07671_),
    .Y(net3770));
 BUFx2_ASAP7_75t_R hold1647 (.A(data_rdata_i[2]),
    .Y(net3771));
 BUFx2_ASAP7_75t_R hold1648 (.A(net49),
    .Y(net3772));
 BUFx2_ASAP7_75t_R hold1649 (.A(_07470_),
    .Y(net3773));
 BUFx2_ASAP7_75t_R hold1650 (.A(data_rdata_i[5]),
    .Y(net3774));
 BUFx2_ASAP7_75t_R hold1651 (.A(net3953),
    .Y(net3775));
 BUFx2_ASAP7_75t_R hold1652 (.A(net3955),
    .Y(net3776));
 BUFx2_ASAP7_75t_R hold1653 (.A(net3957),
    .Y(net3777));
 BUFx2_ASAP7_75t_R hold1654 (.A(net3959),
    .Y(net3778));
 BUFx2_ASAP7_75t_R hold1655 (.A(data_rdata_i[0]),
    .Y(net3779));
 BUFx2_ASAP7_75t_R hold1656 (.A(net27),
    .Y(net3780));
 BUFx2_ASAP7_75t_R hold1657 (.A(net3937),
    .Y(net3781));
 BUFx2_ASAP7_75t_R hold1658 (.A(net3939),
    .Y(net3782));
 BUFx2_ASAP7_75t_R hold1659 (.A(net3941),
    .Y(net3783));
 BUFx2_ASAP7_75t_R hold1660 (.A(net3943),
    .Y(net3784));
 BUFx2_ASAP7_75t_R hold1661 (.A(data_rdata_i[4]),
    .Y(net3785));
 BUFx2_ASAP7_75t_R hold1662 (.A(data_rdata_i[1]),
    .Y(net3786));
 BUFx2_ASAP7_75t_R hold1663 (.A(net3904),
    .Y(net3787));
 BUFx2_ASAP7_75t_R hold1664 (.A(net3906),
    .Y(net3788));
 BUFx2_ASAP7_75t_R hold1665 (.A(net3908),
    .Y(net3789));
 BUFx2_ASAP7_75t_R hold1666 (.A(net3921),
    .Y(net3790));
 BUFx2_ASAP7_75t_R hold1667 (.A(net3923),
    .Y(net3791));
 BUFx2_ASAP7_75t_R hold1668 (.A(net3925),
    .Y(net3792));
 BUFx2_ASAP7_75t_R hold1669 (.A(net3913),
    .Y(net3793));
 BUFx2_ASAP7_75t_R hold1670 (.A(net3915),
    .Y(net3794));
 BUFx2_ASAP7_75t_R hold1671 (.A(net3917),
    .Y(net3795));
 BUFx2_ASAP7_75t_R hold1672 (.A(net3967),
    .Y(net3796));
 BUFx2_ASAP7_75t_R hold1673 (.A(net3969),
    .Y(net3797));
 BUFx2_ASAP7_75t_R hold1674 (.A(net3971),
    .Y(net3798));
 BUFx2_ASAP7_75t_R hold1675 (.A(net2395),
    .Y(net3799));
 BUFx2_ASAP7_75t_R hold1676 (.A(_04364_),
    .Y(net3800));
 BUFx2_ASAP7_75t_R hold1677 (.A(net2396),
    .Y(net3801));
 BUFx2_ASAP7_75t_R hold1678 (.A(net3973),
    .Y(net3802));
 BUFx2_ASAP7_75t_R hold1679 (.A(net3975),
    .Y(net3803));
 BUFx2_ASAP7_75t_R hold1680 (.A(net3977),
    .Y(net3804));
 BUFx2_ASAP7_75t_R hold1681 (.A(net2413),
    .Y(net3805));
 BUFx2_ASAP7_75t_R hold1682 (.A(_04350_),
    .Y(net3806));
 BUFx2_ASAP7_75t_R hold1683 (.A(net2414),
    .Y(net3807));
 BUFx2_ASAP7_75t_R hold1684 (.A(net3985),
    .Y(net3808));
 BUFx2_ASAP7_75t_R hold1685 (.A(net3987),
    .Y(net3809));
 BUFx2_ASAP7_75t_R hold1686 (.A(net3989),
    .Y(net3810));
 BUFx2_ASAP7_75t_R hold1687 (.A(net2419),
    .Y(net3811));
 BUFx2_ASAP7_75t_R hold1688 (.A(_04368_),
    .Y(net3812));
 BUFx2_ASAP7_75t_R hold1689 (.A(net2420),
    .Y(net3813));
 BUFx2_ASAP7_75t_R hold1690 (.A(net3979),
    .Y(net3814));
 BUFx2_ASAP7_75t_R hold1691 (.A(net3981),
    .Y(net3815));
 BUFx2_ASAP7_75t_R hold1692 (.A(net3983),
    .Y(net3816));
 BUFx2_ASAP7_75t_R hold1693 (.A(net2416),
    .Y(net3817));
 BUFx2_ASAP7_75t_R hold1694 (.A(_04346_),
    .Y(net3818));
 BUFx2_ASAP7_75t_R hold1695 (.A(net2417),
    .Y(net3819));
 BUFx2_ASAP7_75t_R hold1696 (.A(net3990),
    .Y(net3820));
 BUFx2_ASAP7_75t_R hold1697 (.A(net3992),
    .Y(net3821));
 BUFx2_ASAP7_75t_R hold1698 (.A(net3994),
    .Y(net3822));
 BUFx2_ASAP7_75t_R hold1699 (.A(net2422),
    .Y(net3823));
 BUFx2_ASAP7_75t_R hold1700 (.A(_04348_),
    .Y(net3824));
 BUFx2_ASAP7_75t_R hold1701 (.A(net2423),
    .Y(net3825));
 BUFx2_ASAP7_75t_R hold1702 (.A(net4005),
    .Y(net3826));
 BUFx2_ASAP7_75t_R hold1703 (.A(net4007),
    .Y(net3827));
 BUFx2_ASAP7_75t_R hold1704 (.A(net4009),
    .Y(net3828));
 BUFx2_ASAP7_75t_R hold1705 (.A(net2440),
    .Y(net3829));
 BUFx2_ASAP7_75t_R hold1706 (.A(_04352_),
    .Y(net3830));
 BUFx2_ASAP7_75t_R hold1707 (.A(net2441),
    .Y(net3831));
 BUFx2_ASAP7_75t_R hold1708 (.A(net3995),
    .Y(net3832));
 BUFx2_ASAP7_75t_R hold1709 (.A(net3997),
    .Y(net3833));
 BUFx2_ASAP7_75t_R hold1710 (.A(net3999),
    .Y(net3834));
 BUFx2_ASAP7_75t_R hold1711 (.A(net2437),
    .Y(net3835));
 BUFx2_ASAP7_75t_R hold1712 (.A(_04363_),
    .Y(net3836));
 BUFx2_ASAP7_75t_R hold1713 (.A(net2438),
    .Y(net3837));
 BUFx2_ASAP7_75t_R hold1714 (.A(net4000),
    .Y(net3838));
 BUFx2_ASAP7_75t_R hold1715 (.A(net4002),
    .Y(net3839));
 BUFx2_ASAP7_75t_R hold1716 (.A(net4004),
    .Y(net3840));
 BUFx2_ASAP7_75t_R hold1717 (.A(net2458),
    .Y(net3841));
 BUFx2_ASAP7_75t_R hold1718 (.A(_04365_),
    .Y(net3842));
 BUFx2_ASAP7_75t_R hold1719 (.A(net2459),
    .Y(net3843));
 BUFx2_ASAP7_75t_R hold1720 (.A(net4010),
    .Y(net3844));
 BUFx2_ASAP7_75t_R hold1721 (.A(net4012),
    .Y(net3845));
 BUFx2_ASAP7_75t_R hold1722 (.A(net4014),
    .Y(net3846));
 BUFx2_ASAP7_75t_R hold1723 (.A(net2497),
    .Y(net3847));
 BUFx2_ASAP7_75t_R hold1724 (.A(_04356_),
    .Y(net3848));
 BUFx2_ASAP7_75t_R hold1725 (.A(net2498),
    .Y(net3849));
 BUFx2_ASAP7_75t_R hold1726 (.A(net4015),
    .Y(net3850));
 BUFx2_ASAP7_75t_R hold1727 (.A(net4017),
    .Y(net3851));
 BUFx2_ASAP7_75t_R hold1728 (.A(net4019),
    .Y(net3852));
 BUFx2_ASAP7_75t_R hold1729 (.A(net2482),
    .Y(net3853));
 BUFx2_ASAP7_75t_R hold1730 (.A(_04359_),
    .Y(net3854));
 BUFx2_ASAP7_75t_R hold1731 (.A(net2483),
    .Y(net3855));
 BUFx2_ASAP7_75t_R hold1732 (.A(net4020),
    .Y(net3856));
 BUFx2_ASAP7_75t_R hold1733 (.A(net4022),
    .Y(net3857));
 BUFx2_ASAP7_75t_R hold1734 (.A(net4024),
    .Y(net3858));
 BUFx2_ASAP7_75t_R hold1735 (.A(net2494),
    .Y(net3859));
 BUFx2_ASAP7_75t_R hold1736 (.A(_04354_),
    .Y(net3860));
 BUFx2_ASAP7_75t_R hold1737 (.A(net2495),
    .Y(net3861));
 BUFx2_ASAP7_75t_R hold1738 (.A(net4035),
    .Y(net3862));
 BUFx2_ASAP7_75t_R hold1739 (.A(net4037),
    .Y(net3863));
 BUFx2_ASAP7_75t_R hold1740 (.A(net4039),
    .Y(net3864));
 BUFx2_ASAP7_75t_R hold1741 (.A(net2510),
    .Y(net3865));
 BUFx2_ASAP7_75t_R hold1742 (.A(_04369_),
    .Y(net3866));
 BUFx2_ASAP7_75t_R hold1743 (.A(net2511),
    .Y(net3867));
 BUFx2_ASAP7_75t_R hold1744 (.A(net4030),
    .Y(net3868));
 BUFx2_ASAP7_75t_R hold1745 (.A(net4032),
    .Y(net3869));
 BUFx2_ASAP7_75t_R hold1746 (.A(net4034),
    .Y(net3870));
 BUFx2_ASAP7_75t_R hold1747 (.A(net2526),
    .Y(net3871));
 BUFx2_ASAP7_75t_R hold1748 (.A(_04347_),
    .Y(net3872));
 BUFx2_ASAP7_75t_R hold1749 (.A(net2527),
    .Y(net3873));
 BUFx2_ASAP7_75t_R hold1750 (.A(net4025),
    .Y(net3874));
 BUFx2_ASAP7_75t_R hold1751 (.A(net4027),
    .Y(net3875));
 BUFx2_ASAP7_75t_R hold1752 (.A(net4029),
    .Y(net3876));
 BUFx2_ASAP7_75t_R hold1753 (.A(net2550),
    .Y(net3877));
 BUFx2_ASAP7_75t_R hold1754 (.A(_04349_),
    .Y(net3878));
 BUFx2_ASAP7_75t_R hold1755 (.A(net2551),
    .Y(net3879));
 BUFx2_ASAP7_75t_R hold1756 (.A(net4040),
    .Y(net3880));
 BUFx2_ASAP7_75t_R hold1757 (.A(net4042),
    .Y(net3881));
 BUFx2_ASAP7_75t_R hold1758 (.A(net4044),
    .Y(net3882));
 BUFx2_ASAP7_75t_R hold1759 (.A(net2563),
    .Y(net3883));
 BUFx2_ASAP7_75t_R hold1760 (.A(_04360_),
    .Y(net3884));
 BUFx2_ASAP7_75t_R hold1761 (.A(net2564),
    .Y(net3885));
 BUFx2_ASAP7_75t_R hold1762 (.A(net4050),
    .Y(net3886));
 BUFx2_ASAP7_75t_R hold1763 (.A(net4052),
    .Y(net3887));
 BUFx2_ASAP7_75t_R hold1764 (.A(net4054),
    .Y(net3888));
 BUFx2_ASAP7_75t_R hold1765 (.A(net2569),
    .Y(net3889));
 BUFx2_ASAP7_75t_R hold1766 (.A(_04353_),
    .Y(net3890));
 BUFx2_ASAP7_75t_R hold1767 (.A(net2570),
    .Y(net3891));
 BUFx2_ASAP7_75t_R hold1768 (.A(net4045),
    .Y(net3892));
 BUFx2_ASAP7_75t_R hold1769 (.A(net4047),
    .Y(net3893));
 BUFx2_ASAP7_75t_R hold1770 (.A(net4049),
    .Y(net3894));
 BUFx2_ASAP7_75t_R hold1771 (.A(net2572),
    .Y(net3895));
 BUFx2_ASAP7_75t_R hold1772 (.A(_04355_),
    .Y(net3896));
 BUFx2_ASAP7_75t_R hold1773 (.A(net2573),
    .Y(net3897));
 BUFx2_ASAP7_75t_R hold1774 (.A(net4055),
    .Y(net3898));
 BUFx2_ASAP7_75t_R hold1775 (.A(net4057),
    .Y(net3899));
 BUFx2_ASAP7_75t_R hold1776 (.A(net4059),
    .Y(net3900));
 BUFx2_ASAP7_75t_R hold1777 (.A(net2620),
    .Y(net3901));
 BUFx2_ASAP7_75t_R hold1778 (.A(_04357_),
    .Y(net3902));
 BUFx2_ASAP7_75t_R hold1779 (.A(net2621),
    .Y(net3903));
 BUFx2_ASAP7_75t_R hold1780 (.A(data_rdata_i[28]),
    .Y(net3904));
 BUFx2_ASAP7_75t_R hold1781 (.A(net3787),
    .Y(net3905));
 BUFx2_ASAP7_75t_R hold1782 (.A(net2397),
    .Y(net3906));
 BUFx2_ASAP7_75t_R hold1783 (.A(net3788),
    .Y(net3907));
 BUFx2_ASAP7_75t_R hold1784 (.A(net47),
    .Y(net3908));
 BUFx2_ASAP7_75t_R hold1785 (.A(net3789),
    .Y(net3909));
 BUFx2_ASAP7_75t_R hold1786 (.A(net2398),
    .Y(net3910));
 BUFx2_ASAP7_75t_R hold1787 (.A(_04366_),
    .Y(net3911));
 BUFx2_ASAP7_75t_R hold1788 (.A(net2399),
    .Y(net3912));
 BUFx2_ASAP7_75t_R hold1789 (.A(data_rdata_i[13]),
    .Y(net3913));
 BUFx2_ASAP7_75t_R hold1790 (.A(net3793),
    .Y(net3914));
 BUFx2_ASAP7_75t_R hold1791 (.A(net2433),
    .Y(net3915));
 BUFx2_ASAP7_75t_R hold1792 (.A(net3794),
    .Y(net3916));
 BUFx2_ASAP7_75t_R hold1793 (.A(net31),
    .Y(net3917));
 BUFx2_ASAP7_75t_R hold1794 (.A(net3795),
    .Y(net3918));
 BUFx2_ASAP7_75t_R hold1795 (.A(net2434),
    .Y(net3919));
 BUFx2_ASAP7_75t_R hold1796 (.A(_04351_),
    .Y(net3920));
 BUFx2_ASAP7_75t_R hold1797 (.A(data_rdata_i[20]),
    .Y(net3921));
 BUFx2_ASAP7_75t_R hold1798 (.A(net3790),
    .Y(net3922));
 BUFx2_ASAP7_75t_R hold1799 (.A(net2487),
    .Y(net3923));
 BUFx2_ASAP7_75t_R hold1800 (.A(net3791),
    .Y(net3924));
 BUFx2_ASAP7_75t_R hold1801 (.A(net39),
    .Y(net3925));
 BUFx2_ASAP7_75t_R hold1802 (.A(net3792),
    .Y(net3926));
 BUFx2_ASAP7_75t_R hold1803 (.A(net2488),
    .Y(net3927));
 BUFx2_ASAP7_75t_R hold1804 (.A(_04358_),
    .Y(net3928));
 BUFx2_ASAP7_75t_R hold1805 (.A(data_rdata_i[23]),
    .Y(net3929));
 BUFx2_ASAP7_75t_R hold1806 (.A(net3759),
    .Y(net3930));
 BUFx2_ASAP7_75t_R hold1807 (.A(net2565),
    .Y(net3931));
 BUFx2_ASAP7_75t_R hold1808 (.A(net3760),
    .Y(net3932));
 BUFx2_ASAP7_75t_R hold1809 (.A(net42),
    .Y(net3933));
 BUFx2_ASAP7_75t_R hold1810 (.A(net3761),
    .Y(net3934));
 BUFx2_ASAP7_75t_R hold1811 (.A(net2566),
    .Y(net3935));
 BUFx2_ASAP7_75t_R hold1812 (.A(_04361_),
    .Y(net3936));
 BUFx2_ASAP7_75t_R hold1813 (.A(data_rdata_i[24]),
    .Y(net3937));
 BUFx2_ASAP7_75t_R hold1814 (.A(net3781),
    .Y(net3938));
 BUFx2_ASAP7_75t_R hold1815 (.A(net2391),
    .Y(net3939));
 BUFx2_ASAP7_75t_R hold1816 (.A(net3782),
    .Y(net3940));
 BUFx2_ASAP7_75t_R hold1817 (.A(net43),
    .Y(net3941));
 BUFx2_ASAP7_75t_R hold1818 (.A(net3783),
    .Y(net3942));
 BUFx2_ASAP7_75t_R hold1819 (.A(net2392),
    .Y(net3943));
 BUFx2_ASAP7_75t_R hold1820 (.A(net3784),
    .Y(net3944));
 BUFx2_ASAP7_75t_R hold1821 (.A(fetch_enable_i),
    .Y(net3945));
 BUFx2_ASAP7_75t_R hold1822 (.A(net3066),
    .Y(net3946));
 BUFx2_ASAP7_75t_R hold1823 (.A(net61),
    .Y(net3947));
 BUFx2_ASAP7_75t_R hold1824 (.A(net3067),
    .Y(net3948));
 BUFx2_ASAP7_75t_R hold1825 (.A(_12717_),
    .Y(net3949));
 BUFx2_ASAP7_75t_R hold1826 (.A(net3068),
    .Y(net3950));
 BUFx2_ASAP7_75t_R hold1827 (.A(_04470_),
    .Y(net3951));
 BUFx2_ASAP7_75t_R hold1828 (.A(net3069),
    .Y(net3952));
 BUFx2_ASAP7_75t_R hold1829 (.A(data_rdata_i[29]),
    .Y(net3953));
 BUFx2_ASAP7_75t_R hold1830 (.A(net3775),
    .Y(net3954));
 BUFx2_ASAP7_75t_R hold1831 (.A(net2475),
    .Y(net3955));
 BUFx2_ASAP7_75t_R hold1832 (.A(net3776),
    .Y(net3956));
 BUFx2_ASAP7_75t_R hold1833 (.A(net48),
    .Y(net3957));
 BUFx2_ASAP7_75t_R hold1834 (.A(net3777),
    .Y(net3958));
 BUFx2_ASAP7_75t_R hold1835 (.A(net2476),
    .Y(net3959));
 BUFx2_ASAP7_75t_R hold1836 (.A(test_en_i),
    .Y(net3960));
 BUFx2_ASAP7_75t_R hold1837 (.A(net3139),
    .Y(net3961));
 BUFx2_ASAP7_75t_R hold1838 (.A(net149),
    .Y(net3962));
 BUFx2_ASAP7_75t_R hold1839 (.A(net3140),
    .Y(net3963));
 BUFx2_ASAP7_75t_R hold1840 (.A(_06717_),
    .Y(net3964));
 BUFx2_ASAP7_75t_R hold1841 (.A(net3141),
    .Y(net3965));
 BUFx2_ASAP7_75t_R hold1842 (.A(_00008_),
    .Y(net3966));
 BUFx2_ASAP7_75t_R hold1843 (.A(data_rdata_i[26]),
    .Y(net3967));
 BUFx2_ASAP7_75t_R hold1844 (.A(net3796),
    .Y(net3968));
 BUFx2_ASAP7_75t_R hold1845 (.A(net2394),
    .Y(net3969));
 BUFx2_ASAP7_75t_R hold1846 (.A(net3797),
    .Y(net3970));
 BUFx2_ASAP7_75t_R hold1847 (.A(net45),
    .Y(net3971));
 BUFx2_ASAP7_75t_R hold1848 (.A(net3798),
    .Y(net3972));
 BUFx2_ASAP7_75t_R hold1849 (.A(data_rdata_i[12]),
    .Y(net3973));
 BUFx2_ASAP7_75t_R hold1850 (.A(net3802),
    .Y(net3974));
 BUFx2_ASAP7_75t_R hold1851 (.A(net2412),
    .Y(net3975));
 BUFx2_ASAP7_75t_R hold1852 (.A(net3803),
    .Y(net3976));
 BUFx2_ASAP7_75t_R hold1853 (.A(net30),
    .Y(net3977));
 BUFx2_ASAP7_75t_R hold1854 (.A(net3804),
    .Y(net3978));
 BUFx2_ASAP7_75t_R hold1855 (.A(data_rdata_i[8]),
    .Y(net3979));
 BUFx2_ASAP7_75t_R hold1856 (.A(net3814),
    .Y(net3980));
 BUFx2_ASAP7_75t_R hold1857 (.A(net2415),
    .Y(net3981));
 BUFx2_ASAP7_75t_R hold1858 (.A(net3815),
    .Y(net3982));
 BUFx2_ASAP7_75t_R hold1859 (.A(net57),
    .Y(net3983));
 BUFx2_ASAP7_75t_R hold1860 (.A(net3816),
    .Y(net3984));
 BUFx2_ASAP7_75t_R hold1861 (.A(data_rdata_i[30]),
    .Y(net3985));
 BUFx2_ASAP7_75t_R hold1862 (.A(net3808),
    .Y(net3986));
 BUFx2_ASAP7_75t_R hold1863 (.A(net2418),
    .Y(net3987));
 BUFx2_ASAP7_75t_R hold1864 (.A(net3809),
    .Y(net3988));
 BUFx2_ASAP7_75t_R hold1865 (.A(net50),
    .Y(net3989));
 BUFx2_ASAP7_75t_R hold1866 (.A(data_rdata_i[10]),
    .Y(net3990));
 BUFx2_ASAP7_75t_R hold1867 (.A(net3820),
    .Y(net3991));
 BUFx2_ASAP7_75t_R hold1868 (.A(net2421),
    .Y(net3992));
 BUFx2_ASAP7_75t_R hold1869 (.A(net3821),
    .Y(net3993));
 BUFx2_ASAP7_75t_R hold1870 (.A(net28),
    .Y(net3994));
 BUFx2_ASAP7_75t_R hold1871 (.A(data_rdata_i[25]),
    .Y(net3995));
 BUFx2_ASAP7_75t_R hold1872 (.A(net3832),
    .Y(net3996));
 BUFx2_ASAP7_75t_R hold1873 (.A(net2436),
    .Y(net3997));
 BUFx2_ASAP7_75t_R hold1874 (.A(net3833),
    .Y(net3998));
 BUFx2_ASAP7_75t_R hold1875 (.A(net44),
    .Y(net3999));
 BUFx2_ASAP7_75t_R hold1876 (.A(data_rdata_i[27]),
    .Y(net4000));
 BUFx2_ASAP7_75t_R hold1877 (.A(net3838),
    .Y(net4001));
 BUFx2_ASAP7_75t_R hold1878 (.A(net2457),
    .Y(net4002));
 BUFx2_ASAP7_75t_R hold1879 (.A(net3839),
    .Y(net4003));
 BUFx2_ASAP7_75t_R hold1880 (.A(net46),
    .Y(net4004));
 BUFx2_ASAP7_75t_R hold1881 (.A(data_rdata_i[14]),
    .Y(net4005));
 BUFx2_ASAP7_75t_R hold1882 (.A(net3826),
    .Y(net4006));
 BUFx2_ASAP7_75t_R hold1883 (.A(net2439),
    .Y(net4007));
 BUFx2_ASAP7_75t_R hold1884 (.A(net3827),
    .Y(net4008));
 BUFx2_ASAP7_75t_R hold1885 (.A(net32),
    .Y(net4009));
 BUFx2_ASAP7_75t_R hold1886 (.A(data_rdata_i[18]),
    .Y(net4010));
 BUFx2_ASAP7_75t_R hold1887 (.A(net3844),
    .Y(net4011));
 BUFx2_ASAP7_75t_R hold1888 (.A(net2496),
    .Y(net4012));
 BUFx2_ASAP7_75t_R hold1889 (.A(net3845),
    .Y(net4013));
 BUFx2_ASAP7_75t_R hold1890 (.A(net36),
    .Y(net4014));
 BUFx2_ASAP7_75t_R hold1891 (.A(data_rdata_i[21]),
    .Y(net4015));
 BUFx2_ASAP7_75t_R hold1892 (.A(net3850),
    .Y(net4016));
 BUFx2_ASAP7_75t_R hold1893 (.A(net2481),
    .Y(net4017));
 BUFx2_ASAP7_75t_R hold1894 (.A(net3851),
    .Y(net4018));
 BUFx2_ASAP7_75t_R hold1895 (.A(net40),
    .Y(net4019));
 BUFx2_ASAP7_75t_R hold1896 (.A(data_rdata_i[16]),
    .Y(net4020));
 BUFx2_ASAP7_75t_R hold1897 (.A(net3856),
    .Y(net4021));
 BUFx2_ASAP7_75t_R hold1898 (.A(net2493),
    .Y(net4022));
 BUFx2_ASAP7_75t_R hold1899 (.A(net3857),
    .Y(net4023));
 BUFx2_ASAP7_75t_R hold1900 (.A(net34),
    .Y(net4024));
 BUFx2_ASAP7_75t_R hold1901 (.A(data_rdata_i[11]),
    .Y(net4025));
 BUFx2_ASAP7_75t_R hold1902 (.A(net3874),
    .Y(net4026));
 BUFx2_ASAP7_75t_R hold1903 (.A(net2549),
    .Y(net4027));
 BUFx2_ASAP7_75t_R hold1904 (.A(net3875),
    .Y(net4028));
 BUFx2_ASAP7_75t_R hold1905 (.A(net29),
    .Y(net4029));
 BUFx2_ASAP7_75t_R hold1906 (.A(data_rdata_i[9]),
    .Y(net4030));
 BUFx2_ASAP7_75t_R hold1907 (.A(net3868),
    .Y(net4031));
 BUFx2_ASAP7_75t_R hold1908 (.A(net2525),
    .Y(net4032));
 BUFx2_ASAP7_75t_R hold1909 (.A(net3869),
    .Y(net4033));
 BUFx2_ASAP7_75t_R hold1910 (.A(net58),
    .Y(net4034));
 BUFx2_ASAP7_75t_R hold1911 (.A(data_rdata_i[31]),
    .Y(net4035));
 BUFx2_ASAP7_75t_R hold1912 (.A(net3862),
    .Y(net4036));
 BUFx2_ASAP7_75t_R hold1913 (.A(net2509),
    .Y(net4037));
 BUFx2_ASAP7_75t_R hold1914 (.A(net3863),
    .Y(net4038));
 BUFx2_ASAP7_75t_R hold1915 (.A(net51),
    .Y(net4039));
 BUFx2_ASAP7_75t_R hold1916 (.A(data_rdata_i[22]),
    .Y(net4040));
 BUFx2_ASAP7_75t_R hold1917 (.A(net3880),
    .Y(net4041));
 BUFx2_ASAP7_75t_R hold1918 (.A(net2562),
    .Y(net4042));
 BUFx2_ASAP7_75t_R hold1919 (.A(net3881),
    .Y(net4043));
 BUFx2_ASAP7_75t_R hold1920 (.A(net41),
    .Y(net4044));
 BUFx2_ASAP7_75t_R hold1921 (.A(data_rdata_i[17]),
    .Y(net4045));
 BUFx2_ASAP7_75t_R hold1922 (.A(net3892),
    .Y(net4046));
 BUFx2_ASAP7_75t_R hold1923 (.A(net2571),
    .Y(net4047));
 BUFx2_ASAP7_75t_R hold1924 (.A(net3893),
    .Y(net4048));
 BUFx2_ASAP7_75t_R hold1925 (.A(net35),
    .Y(net4049));
 BUFx2_ASAP7_75t_R hold1926 (.A(data_rdata_i[15]),
    .Y(net4050));
 BUFx2_ASAP7_75t_R hold1927 (.A(net3886),
    .Y(net4051));
 BUFx2_ASAP7_75t_R hold1928 (.A(net2568),
    .Y(net4052));
 BUFx2_ASAP7_75t_R hold1929 (.A(net3887),
    .Y(net4053));
 BUFx2_ASAP7_75t_R hold1930 (.A(net33),
    .Y(net4054));
 BUFx2_ASAP7_75t_R hold1931 (.A(data_rdata_i[19]),
    .Y(net4055));
 BUFx2_ASAP7_75t_R hold1932 (.A(net3898),
    .Y(net4056));
 BUFx2_ASAP7_75t_R hold1933 (.A(net2619),
    .Y(net4057));
 BUFx2_ASAP7_75t_R hold1934 (.A(net3899),
    .Y(net4058));
 BUFx2_ASAP7_75t_R hold1935 (.A(net37),
    .Y(net4059));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx10_ASAP7_75t_R FILLER_0_134 ();
 DECAPx10_ASAP7_75t_R FILLER_0_156 ();
 DECAPx10_ASAP7_75t_R FILLER_0_178 ();
 DECAPx10_ASAP7_75t_R FILLER_0_200 ();
 DECAPx10_ASAP7_75t_R FILLER_0_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_505 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_0_546 ();
 DECAPx1_ASAP7_75t_R FILLER_0_625 ();
 DECAPx10_ASAP7_75t_R FILLER_0_790 ();
 DECAPx10_ASAP7_75t_R FILLER_0_812 ();
 DECAPx10_ASAP7_75t_R FILLER_0_834 ();
 DECAPx10_ASAP7_75t_R FILLER_0_856 ();
 DECAPx10_ASAP7_75t_R FILLER_0_878 ();
 DECAPx10_ASAP7_75t_R FILLER_0_900 ();
 FILLER_ASAP7_75t_R FILLER_0_922 ();
 DECAPx2_ASAP7_75t_R FILLER_0_926 ();
 FILLER_ASAP7_75t_R FILLER_0_932 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx10_ASAP7_75t_R FILLER_1_134 ();
 DECAPx10_ASAP7_75t_R FILLER_1_156 ();
 DECAPx10_ASAP7_75t_R FILLER_1_178 ();
 DECAPx10_ASAP7_75t_R FILLER_1_200 ();
 DECAPx10_ASAP7_75t_R FILLER_1_222 ();
 DECAPx2_ASAP7_75t_R FILLER_1_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_250 ();
 FILLER_ASAP7_75t_R FILLER_1_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_443 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_472 ();
 DECAPx1_ASAP7_75t_R FILLER_1_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_561 ();
 FILLER_ASAP7_75t_R FILLER_1_569 ();
 FILLER_ASAP7_75t_R FILLER_1_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_600 ();
 FILLER_ASAP7_75t_R FILLER_1_612 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_686 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_720 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_730 ();
 FILLER_ASAP7_75t_R FILLER_1_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_748 ();
 DECAPx10_ASAP7_75t_R FILLER_1_776 ();
 DECAPx10_ASAP7_75t_R FILLER_1_798 ();
 DECAPx10_ASAP7_75t_R FILLER_1_820 ();
 DECAPx10_ASAP7_75t_R FILLER_1_842 ();
 DECAPx10_ASAP7_75t_R FILLER_1_864 ();
 DECAPx10_ASAP7_75t_R FILLER_1_886 ();
 DECAPx6_ASAP7_75t_R FILLER_1_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_1_922 ();
 DECAPx2_ASAP7_75t_R FILLER_1_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_933 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx10_ASAP7_75t_R FILLER_2_134 ();
 DECAPx10_ASAP7_75t_R FILLER_2_156 ();
 DECAPx10_ASAP7_75t_R FILLER_2_178 ();
 DECAPx10_ASAP7_75t_R FILLER_2_200 ();
 DECAPx10_ASAP7_75t_R FILLER_2_222 ();
 DECAPx6_ASAP7_75t_R FILLER_2_244 ();
 DECAPx1_ASAP7_75t_R FILLER_2_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_2_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_512 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_520 ();
 FILLER_ASAP7_75t_R FILLER_2_588 ();
 FILLER_ASAP7_75t_R FILLER_2_610 ();
 DECAPx1_ASAP7_75t_R FILLER_2_668 ();
 FILLER_ASAP7_75t_R FILLER_2_679 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_2_701 ();
 DECAPx10_ASAP7_75t_R FILLER_2_769 ();
 DECAPx10_ASAP7_75t_R FILLER_2_791 ();
 DECAPx10_ASAP7_75t_R FILLER_2_813 ();
 DECAPx10_ASAP7_75t_R FILLER_2_835 ();
 DECAPx10_ASAP7_75t_R FILLER_2_857 ();
 DECAPx10_ASAP7_75t_R FILLER_2_879 ();
 DECAPx10_ASAP7_75t_R FILLER_2_901 ();
 DECAPx4_ASAP7_75t_R FILLER_2_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_933 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx10_ASAP7_75t_R FILLER_3_134 ();
 DECAPx10_ASAP7_75t_R FILLER_3_156 ();
 DECAPx10_ASAP7_75t_R FILLER_3_178 ();
 DECAPx4_ASAP7_75t_R FILLER_3_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_217 ();
 DECAPx10_ASAP7_75t_R FILLER_3_224 ();
 DECAPx2_ASAP7_75t_R FILLER_3_246 ();
 FILLER_ASAP7_75t_R FILLER_3_252 ();
 DECAPx2_ASAP7_75t_R FILLER_3_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_263 ();
 FILLER_ASAP7_75t_R FILLER_3_292 ();
 FILLER_ASAP7_75t_R FILLER_3_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_455 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_3_467 ();
 FILLER_ASAP7_75t_R FILLER_3_491 ();
 DECAPx1_ASAP7_75t_R FILLER_3_504 ();
 FILLER_ASAP7_75t_R FILLER_3_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_598 ();
 DECAPx1_ASAP7_75t_R FILLER_3_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_691 ();
 DECAPx10_ASAP7_75t_R FILLER_3_755 ();
 DECAPx10_ASAP7_75t_R FILLER_3_777 ();
 DECAPx10_ASAP7_75t_R FILLER_3_799 ();
 DECAPx10_ASAP7_75t_R FILLER_3_821 ();
 DECAPx10_ASAP7_75t_R FILLER_3_843 ();
 DECAPx10_ASAP7_75t_R FILLER_3_865 ();
 DECAPx10_ASAP7_75t_R FILLER_3_887 ();
 DECAPx6_ASAP7_75t_R FILLER_3_909 ();
 FILLER_ASAP7_75t_R FILLER_3_923 ();
 DECAPx2_ASAP7_75t_R FILLER_3_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_933 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx10_ASAP7_75t_R FILLER_4_134 ();
 DECAPx10_ASAP7_75t_R FILLER_4_156 ();
 DECAPx10_ASAP7_75t_R FILLER_4_178 ();
 DECAPx1_ASAP7_75t_R FILLER_4_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_230 ();
 FILLER_ASAP7_75t_R FILLER_4_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_265 ();
 DECAPx1_ASAP7_75t_R FILLER_4_272 ();
 FILLER_ASAP7_75t_R FILLER_4_308 ();
 FILLER_ASAP7_75t_R FILLER_4_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_392 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_512 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_4_620 ();
 DECAPx1_ASAP7_75t_R FILLER_4_676 ();
 DECAPx1_ASAP7_75t_R FILLER_4_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_703 ();
 DECAPx10_ASAP7_75t_R FILLER_4_739 ();
 DECAPx10_ASAP7_75t_R FILLER_4_761 ();
 DECAPx4_ASAP7_75t_R FILLER_4_783 ();
 FILLER_ASAP7_75t_R FILLER_4_793 ();
 DECAPx1_ASAP7_75t_R FILLER_4_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_806 ();
 DECAPx10_ASAP7_75t_R FILLER_4_813 ();
 DECAPx10_ASAP7_75t_R FILLER_4_835 ();
 DECAPx10_ASAP7_75t_R FILLER_4_857 ();
 DECAPx10_ASAP7_75t_R FILLER_4_879 ();
 DECAPx10_ASAP7_75t_R FILLER_4_901 ();
 DECAPx4_ASAP7_75t_R FILLER_4_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_933 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx10_ASAP7_75t_R FILLER_5_134 ();
 DECAPx10_ASAP7_75t_R FILLER_5_156 ();
 DECAPx6_ASAP7_75t_R FILLER_5_178 ();
 FILLER_ASAP7_75t_R FILLER_5_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_200 ();
 DECAPx4_ASAP7_75t_R FILLER_5_207 ();
 FILLER_ASAP7_75t_R FILLER_5_217 ();
 FILLER_ASAP7_75t_R FILLER_5_251 ();
 DECAPx4_ASAP7_75t_R FILLER_5_279 ();
 FILLER_ASAP7_75t_R FILLER_5_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_441 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_5_470 ();
 DECAPx1_ASAP7_75t_R FILLER_5_493 ();
 DECAPx1_ASAP7_75t_R FILLER_5_505 ();
 DECAPx1_ASAP7_75t_R FILLER_5_542 ();
 FILLER_ASAP7_75t_R FILLER_5_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_5_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_691 ();
 DECAPx10_ASAP7_75t_R FILLER_5_725 ();
 DECAPx10_ASAP7_75t_R FILLER_5_747 ();
 FILLER_ASAP7_75t_R FILLER_5_769 ();
 DECAPx2_ASAP7_75t_R FILLER_5_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_790 ();
 DECAPx10_ASAP7_75t_R FILLER_5_817 ();
 DECAPx10_ASAP7_75t_R FILLER_5_839 ();
 DECAPx10_ASAP7_75t_R FILLER_5_861 ();
 DECAPx10_ASAP7_75t_R FILLER_5_883 ();
 DECAPx6_ASAP7_75t_R FILLER_5_905 ();
 DECAPx2_ASAP7_75t_R FILLER_5_919 ();
 DECAPx2_ASAP7_75t_R FILLER_5_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_933 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx10_ASAP7_75t_R FILLER_6_134 ();
 DECAPx10_ASAP7_75t_R FILLER_6_156 ();
 DECAPx4_ASAP7_75t_R FILLER_6_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_188 ();
 DECAPx6_ASAP7_75t_R FILLER_6_215 ();
 DECAPx2_ASAP7_75t_R FILLER_6_229 ();
 FILLER_ASAP7_75t_R FILLER_6_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_258 ();
 DECAPx10_ASAP7_75t_R FILLER_6_271 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_407 ();
 FILLER_ASAP7_75t_R FILLER_6_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_606 ();
 FILLER_ASAP7_75t_R FILLER_6_618 ();
 DECAPx2_ASAP7_75t_R FILLER_6_696 ();
 FILLER_ASAP7_75t_R FILLER_6_707 ();
 DECAPx6_ASAP7_75t_R FILLER_6_715 ();
 DECAPx1_ASAP7_75t_R FILLER_6_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_733 ();
 DECAPx1_ASAP7_75t_R FILLER_6_747 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_758 ();
 DECAPx6_ASAP7_75t_R FILLER_6_787 ();
 DECAPx10_ASAP7_75t_R FILLER_6_807 ();
 DECAPx10_ASAP7_75t_R FILLER_6_829 ();
 DECAPx10_ASAP7_75t_R FILLER_6_851 ();
 DECAPx10_ASAP7_75t_R FILLER_6_873 ();
 DECAPx10_ASAP7_75t_R FILLER_6_895 ();
 DECAPx6_ASAP7_75t_R FILLER_6_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_6_931 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx10_ASAP7_75t_R FILLER_7_134 ();
 DECAPx6_ASAP7_75t_R FILLER_7_156 ();
 DECAPx2_ASAP7_75t_R FILLER_7_170 ();
 FILLER_ASAP7_75t_R FILLER_7_182 ();
 DECAPx2_ASAP7_75t_R FILLER_7_193 ();
 DECAPx1_ASAP7_75t_R FILLER_7_208 ();
 DECAPx10_ASAP7_75t_R FILLER_7_215 ();
 DECAPx2_ASAP7_75t_R FILLER_7_237 ();
 DECAPx10_ASAP7_75t_R FILLER_7_246 ();
 DECAPx6_ASAP7_75t_R FILLER_7_268 ();
 DECAPx6_ASAP7_75t_R FILLER_7_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_302 ();
 FILLER_ASAP7_75t_R FILLER_7_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_408 ();
 FILLER_ASAP7_75t_R FILLER_7_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_457 ();
 FILLER_ASAP7_75t_R FILLER_7_484 ();
 FILLER_ASAP7_75t_R FILLER_7_502 ();
 DECAPx4_ASAP7_75t_R FILLER_7_514 ();
 FILLER_ASAP7_75t_R FILLER_7_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_532 ();
 DECAPx1_ASAP7_75t_R FILLER_7_539 ();
 FILLER_ASAP7_75t_R FILLER_7_554 ();
 DECAPx1_ASAP7_75t_R FILLER_7_668 ();
 FILLER_ASAP7_75t_R FILLER_7_679 ();
 DECAPx10_ASAP7_75t_R FILLER_7_692 ();
 DECAPx6_ASAP7_75t_R FILLER_7_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_728 ();
 FILLER_ASAP7_75t_R FILLER_7_775 ();
 DECAPx10_ASAP7_75t_R FILLER_7_789 ();
 DECAPx10_ASAP7_75t_R FILLER_7_811 ();
 DECAPx10_ASAP7_75t_R FILLER_7_833 ();
 DECAPx10_ASAP7_75t_R FILLER_7_855 ();
 DECAPx10_ASAP7_75t_R FILLER_7_877 ();
 DECAPx10_ASAP7_75t_R FILLER_7_899 ();
 DECAPx1_ASAP7_75t_R FILLER_7_921 ();
 DECAPx2_ASAP7_75t_R FILLER_7_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_933 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx10_ASAP7_75t_R FILLER_8_134 ();
 DECAPx4_ASAP7_75t_R FILLER_8_156 ();
 FILLER_ASAP7_75t_R FILLER_8_166 ();
 DECAPx10_ASAP7_75t_R FILLER_8_232 ();
 DECAPx6_ASAP7_75t_R FILLER_8_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_412 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_430 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_464 ();
 DECAPx10_ASAP7_75t_R FILLER_8_482 ();
 DECAPx2_ASAP7_75t_R FILLER_8_504 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_510 ();
 DECAPx1_ASAP7_75t_R FILLER_8_527 ();
 FILLER_ASAP7_75t_R FILLER_8_561 ();
 FILLER_ASAP7_75t_R FILLER_8_569 ();
 FILLER_ASAP7_75t_R FILLER_8_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_667 ();
 DECAPx1_ASAP7_75t_R FILLER_8_694 ();
 DECAPx1_ASAP7_75t_R FILLER_8_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_715 ();
 DECAPx2_ASAP7_75t_R FILLER_8_735 ();
 FILLER_ASAP7_75t_R FILLER_8_741 ();
 DECAPx10_ASAP7_75t_R FILLER_8_763 ();
 DECAPx10_ASAP7_75t_R FILLER_8_785 ();
 DECAPx10_ASAP7_75t_R FILLER_8_807 ();
 DECAPx10_ASAP7_75t_R FILLER_8_829 ();
 DECAPx10_ASAP7_75t_R FILLER_8_851 ();
 DECAPx10_ASAP7_75t_R FILLER_8_873 ();
 DECAPx10_ASAP7_75t_R FILLER_8_895 ();
 DECAPx6_ASAP7_75t_R FILLER_8_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_8_931 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx10_ASAP7_75t_R FILLER_9_134 ();
 DECAPx10_ASAP7_75t_R FILLER_9_156 ();
 DECAPx2_ASAP7_75t_R FILLER_9_178 ();
 DECAPx6_ASAP7_75t_R FILLER_9_187 ();
 DECAPx1_ASAP7_75t_R FILLER_9_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_241 ();
 DECAPx1_ASAP7_75t_R FILLER_9_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_390 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_411 ();
 FILLER_ASAP7_75t_R FILLER_9_470 ();
 DECAPx6_ASAP7_75t_R FILLER_9_489 ();
 DECAPx1_ASAP7_75t_R FILLER_9_503 ();
 DECAPx2_ASAP7_75t_R FILLER_9_532 ();
 FILLER_ASAP7_75t_R FILLER_9_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_587 ();
 DECAPx4_ASAP7_75t_R FILLER_9_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_676 ();
 DECAPx4_ASAP7_75t_R FILLER_9_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_693 ();
 DECAPx1_ASAP7_75t_R FILLER_9_714 ();
 DECAPx10_ASAP7_75t_R FILLER_9_738 ();
 DECAPx10_ASAP7_75t_R FILLER_9_760 ();
 DECAPx10_ASAP7_75t_R FILLER_9_782 ();
 DECAPx10_ASAP7_75t_R FILLER_9_804 ();
 DECAPx2_ASAP7_75t_R FILLER_9_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_839 ();
 DECAPx10_ASAP7_75t_R FILLER_9_846 ();
 DECAPx10_ASAP7_75t_R FILLER_9_868 ();
 DECAPx10_ASAP7_75t_R FILLER_9_890 ();
 DECAPx4_ASAP7_75t_R FILLER_9_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_9_922 ();
 DECAPx2_ASAP7_75t_R FILLER_9_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_933 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx10_ASAP7_75t_R FILLER_10_134 ();
 DECAPx10_ASAP7_75t_R FILLER_10_156 ();
 DECAPx10_ASAP7_75t_R FILLER_10_178 ();
 DECAPx10_ASAP7_75t_R FILLER_10_200 ();
 DECAPx2_ASAP7_75t_R FILLER_10_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_228 ();
 FILLER_ASAP7_75t_R FILLER_10_258 ();
 FILLER_ASAP7_75t_R FILLER_10_269 ();
 DECAPx4_ASAP7_75t_R FILLER_10_274 ();
 DECAPx2_ASAP7_75t_R FILLER_10_287 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_293 ();
 DECAPx10_ASAP7_75t_R FILLER_10_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_327 ();
 DECAPx1_ASAP7_75t_R FILLER_10_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_394 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_420 ();
 DECAPx2_ASAP7_75t_R FILLER_10_442 ();
 FILLER_ASAP7_75t_R FILLER_10_460 ();
 DECAPx2_ASAP7_75t_R FILLER_10_467 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_473 ();
 DECAPx2_ASAP7_75t_R FILLER_10_507 ();
 DECAPx1_ASAP7_75t_R FILLER_10_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_611 ();
 FILLER_ASAP7_75t_R FILLER_10_638 ();
 DECAPx10_ASAP7_75t_R FILLER_10_661 ();
 DECAPx2_ASAP7_75t_R FILLER_10_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_689 ();
 DECAPx4_ASAP7_75t_R FILLER_10_697 ();
 FILLER_ASAP7_75t_R FILLER_10_707 ();
 DECAPx10_ASAP7_75t_R FILLER_10_736 ();
 FILLER_ASAP7_75t_R FILLER_10_758 ();
 DECAPx2_ASAP7_75t_R FILLER_10_773 ();
 FILLER_ASAP7_75t_R FILLER_10_779 ();
 FILLER_ASAP7_75t_R FILLER_10_788 ();
 DECAPx10_ASAP7_75t_R FILLER_10_796 ();
 DECAPx2_ASAP7_75t_R FILLER_10_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_10_824 ();
 DECAPx10_ASAP7_75t_R FILLER_10_853 ();
 DECAPx10_ASAP7_75t_R FILLER_10_875 ();
 DECAPx10_ASAP7_75t_R FILLER_10_897 ();
 DECAPx6_ASAP7_75t_R FILLER_10_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_933 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx6_ASAP7_75t_R FILLER_11_134 ();
 DECAPx2_ASAP7_75t_R FILLER_11_148 ();
 DECAPx10_ASAP7_75t_R FILLER_11_180 ();
 DECAPx10_ASAP7_75t_R FILLER_11_202 ();
 DECAPx4_ASAP7_75t_R FILLER_11_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_234 ();
 DECAPx1_ASAP7_75t_R FILLER_11_243 ();
 DECAPx2_ASAP7_75t_R FILLER_11_250 ();
 DECAPx10_ASAP7_75t_R FILLER_11_262 ();
 DECAPx10_ASAP7_75t_R FILLER_11_284 ();
 DECAPx2_ASAP7_75t_R FILLER_11_306 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_312 ();
 DECAPx2_ASAP7_75t_R FILLER_11_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_347 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_401 ();
 DECAPx1_ASAP7_75t_R FILLER_11_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_416 ();
 DECAPx1_ASAP7_75t_R FILLER_11_433 ();
 DECAPx2_ASAP7_75t_R FILLER_11_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_448 ();
 DECAPx4_ASAP7_75t_R FILLER_11_456 ();
 FILLER_ASAP7_75t_R FILLER_11_466 ();
 FILLER_ASAP7_75t_R FILLER_11_480 ();
 DECAPx1_ASAP7_75t_R FILLER_11_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_497 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_521 ();
 FILLER_ASAP7_75t_R FILLER_11_547 ();
 DECAPx1_ASAP7_75t_R FILLER_11_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_614 ();
 DECAPx1_ASAP7_75t_R FILLER_11_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_645 ();
 DECAPx10_ASAP7_75t_R FILLER_11_654 ();
 DECAPx2_ASAP7_75t_R FILLER_11_676 ();
 DECAPx10_ASAP7_75t_R FILLER_11_708 ();
 DECAPx10_ASAP7_75t_R FILLER_11_730 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_752 ();
 FILLER_ASAP7_75t_R FILLER_11_775 ();
 DECAPx10_ASAP7_75t_R FILLER_11_803 ();
 DECAPx6_ASAP7_75t_R FILLER_11_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_839 ();
 DECAPx10_ASAP7_75t_R FILLER_11_846 ();
 DECAPx10_ASAP7_75t_R FILLER_11_868 ();
 DECAPx10_ASAP7_75t_R FILLER_11_890 ();
 DECAPx4_ASAP7_75t_R FILLER_11_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_11_922 ();
 DECAPx2_ASAP7_75t_R FILLER_11_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_933 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx10_ASAP7_75t_R FILLER_12_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_156 ();
 DECAPx2_ASAP7_75t_R FILLER_12_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_225 ();
 DECAPx4_ASAP7_75t_R FILLER_12_234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_244 ();
 DECAPx6_ASAP7_75t_R FILLER_12_253 ();
 DECAPx2_ASAP7_75t_R FILLER_12_273 ();
 FILLER_ASAP7_75t_R FILLER_12_279 ();
 DECAPx2_ASAP7_75t_R FILLER_12_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_308 ();
 FILLER_ASAP7_75t_R FILLER_12_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_322 ();
 DECAPx10_ASAP7_75t_R FILLER_12_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_354 ();
 DECAPx1_ASAP7_75t_R FILLER_12_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_396 ();
 DECAPx10_ASAP7_75t_R FILLER_12_407 ();
 FILLER_ASAP7_75t_R FILLER_12_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_441 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_454 ();
 DECAPx1_ASAP7_75t_R FILLER_12_458 ();
 DECAPx2_ASAP7_75t_R FILLER_12_464 ();
 FILLER_ASAP7_75t_R FILLER_12_470 ();
 DECAPx2_ASAP7_75t_R FILLER_12_478 ();
 FILLER_ASAP7_75t_R FILLER_12_484 ();
 DECAPx2_ASAP7_75t_R FILLER_12_492 ();
 DECAPx10_ASAP7_75t_R FILLER_12_510 ();
 DECAPx6_ASAP7_75t_R FILLER_12_532 ();
 DECAPx2_ASAP7_75t_R FILLER_12_551 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_562 ();
 DECAPx1_ASAP7_75t_R FILLER_12_611 ();
 FILLER_ASAP7_75t_R FILLER_12_621 ();
 DECAPx10_ASAP7_75t_R FILLER_12_636 ();
 DECAPx10_ASAP7_75t_R FILLER_12_658 ();
 DECAPx6_ASAP7_75t_R FILLER_12_680 ();
 DECAPx10_ASAP7_75t_R FILLER_12_706 ();
 DECAPx6_ASAP7_75t_R FILLER_12_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_742 ();
 DECAPx2_ASAP7_75t_R FILLER_12_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_764 ();
 DECAPx4_ASAP7_75t_R FILLER_12_777 ();
 DECAPx10_ASAP7_75t_R FILLER_12_793 ();
 DECAPx10_ASAP7_75t_R FILLER_12_815 ();
 DECAPx10_ASAP7_75t_R FILLER_12_837 ();
 DECAPx10_ASAP7_75t_R FILLER_12_859 ();
 DECAPx10_ASAP7_75t_R FILLER_12_881 ();
 DECAPx10_ASAP7_75t_R FILLER_12_903 ();
 DECAPx2_ASAP7_75t_R FILLER_12_925 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_12_931 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx4_ASAP7_75t_R FILLER_13_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_144 ();
 DECAPx2_ASAP7_75t_R FILLER_13_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_165 ();
 DECAPx1_ASAP7_75t_R FILLER_13_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_227 ();
 DECAPx1_ASAP7_75t_R FILLER_13_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_238 ();
 DECAPx4_ASAP7_75t_R FILLER_13_255 ();
 FILLER_ASAP7_75t_R FILLER_13_265 ();
 FILLER_ASAP7_75t_R FILLER_13_273 ();
 DECAPx1_ASAP7_75t_R FILLER_13_289 ();
 DECAPx1_ASAP7_75t_R FILLER_13_301 ();
 DECAPx6_ASAP7_75t_R FILLER_13_331 ();
 DECAPx2_ASAP7_75t_R FILLER_13_345 ();
 DECAPx4_ASAP7_75t_R FILLER_13_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_408 ();
 DECAPx4_ASAP7_75t_R FILLER_13_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_441 ();
 DECAPx1_ASAP7_75t_R FILLER_13_465 ();
 DECAPx6_ASAP7_75t_R FILLER_13_472 ();
 DECAPx1_ASAP7_75t_R FILLER_13_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_496 ();
 DECAPx10_ASAP7_75t_R FILLER_13_502 ();
 DECAPx6_ASAP7_75t_R FILLER_13_524 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_546 ();
 DECAPx1_ASAP7_75t_R FILLER_13_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_600 ();
 DECAPx4_ASAP7_75t_R FILLER_13_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_621 ();
 DECAPx1_ASAP7_75t_R FILLER_13_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_646 ();
 DECAPx6_ASAP7_75t_R FILLER_13_652 ();
 DECAPx1_ASAP7_75t_R FILLER_13_666 ();
 DECAPx10_ASAP7_75t_R FILLER_13_683 ();
 DECAPx10_ASAP7_75t_R FILLER_13_705 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_727 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_13_737 ();
 DECAPx10_ASAP7_75t_R FILLER_13_760 ();
 DECAPx10_ASAP7_75t_R FILLER_13_782 ();
 DECAPx10_ASAP7_75t_R FILLER_13_804 ();
 DECAPx10_ASAP7_75t_R FILLER_13_826 ();
 DECAPx10_ASAP7_75t_R FILLER_13_848 ();
 DECAPx10_ASAP7_75t_R FILLER_13_870 ();
 DECAPx10_ASAP7_75t_R FILLER_13_892 ();
 DECAPx4_ASAP7_75t_R FILLER_13_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_924 ();
 DECAPx2_ASAP7_75t_R FILLER_13_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_933 ();
 DECAPx10_ASAP7_75t_R FILLER_14_2 ();
 DECAPx10_ASAP7_75t_R FILLER_14_24 ();
 DECAPx10_ASAP7_75t_R FILLER_14_46 ();
 DECAPx10_ASAP7_75t_R FILLER_14_68 ();
 DECAPx10_ASAP7_75t_R FILLER_14_90 ();
 DECAPx10_ASAP7_75t_R FILLER_14_112 ();
 DECAPx4_ASAP7_75t_R FILLER_14_134 ();
 FILLER_ASAP7_75t_R FILLER_14_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_191 ();
 DECAPx2_ASAP7_75t_R FILLER_14_207 ();
 FILLER_ASAP7_75t_R FILLER_14_213 ();
 DECAPx1_ASAP7_75t_R FILLER_14_223 ();
 DECAPx6_ASAP7_75t_R FILLER_14_249 ();
 DECAPx1_ASAP7_75t_R FILLER_14_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_267 ();
 DECAPx1_ASAP7_75t_R FILLER_14_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_294 ();
 DECAPx1_ASAP7_75t_R FILLER_14_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_307 ();
 DECAPx6_ASAP7_75t_R FILLER_14_314 ();
 DECAPx2_ASAP7_75t_R FILLER_14_328 ();
 DECAPx10_ASAP7_75t_R FILLER_14_340 ();
 DECAPx2_ASAP7_75t_R FILLER_14_362 ();
 FILLER_ASAP7_75t_R FILLER_14_368 ();
 FILLER_ASAP7_75t_R FILLER_14_382 ();
 DECAPx2_ASAP7_75t_R FILLER_14_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_459 ();
 DECAPx10_ASAP7_75t_R FILLER_14_470 ();
 FILLER_ASAP7_75t_R FILLER_14_492 ();
 DECAPx6_ASAP7_75t_R FILLER_14_511 ();
 DECAPx1_ASAP7_75t_R FILLER_14_525 ();
 DECAPx1_ASAP7_75t_R FILLER_14_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_573 ();
 DECAPx4_ASAP7_75t_R FILLER_14_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_589 ();
 FILLER_ASAP7_75t_R FILLER_14_597 ();
 DECAPx10_ASAP7_75t_R FILLER_14_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_626 ();
 DECAPx10_ASAP7_75t_R FILLER_14_638 ();
 DECAPx1_ASAP7_75t_R FILLER_14_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_664 ();
 DECAPx6_ASAP7_75t_R FILLER_14_691 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_705 ();
 DECAPx1_ASAP7_75t_R FILLER_14_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_724 ();
 DECAPx10_ASAP7_75t_R FILLER_14_767 ();
 DECAPx10_ASAP7_75t_R FILLER_14_789 ();
 DECAPx10_ASAP7_75t_R FILLER_14_811 ();
 DECAPx10_ASAP7_75t_R FILLER_14_833 ();
 DECAPx10_ASAP7_75t_R FILLER_14_855 ();
 DECAPx10_ASAP7_75t_R FILLER_14_877 ();
 DECAPx10_ASAP7_75t_R FILLER_14_899 ();
 DECAPx4_ASAP7_75t_R FILLER_14_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_14_931 ();
 DECAPx10_ASAP7_75t_R FILLER_15_2 ();
 DECAPx10_ASAP7_75t_R FILLER_15_24 ();
 DECAPx10_ASAP7_75t_R FILLER_15_46 ();
 DECAPx10_ASAP7_75t_R FILLER_15_68 ();
 DECAPx6_ASAP7_75t_R FILLER_15_90 ();
 FILLER_ASAP7_75t_R FILLER_15_104 ();
 DECAPx6_ASAP7_75t_R FILLER_15_144 ();
 DECAPx10_ASAP7_75t_R FILLER_15_161 ();
 DECAPx10_ASAP7_75t_R FILLER_15_183 ();
 DECAPx10_ASAP7_75t_R FILLER_15_205 ();
 DECAPx1_ASAP7_75t_R FILLER_15_239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_249 ();
 DECAPx10_ASAP7_75t_R FILLER_15_286 ();
 DECAPx6_ASAP7_75t_R FILLER_15_308 ();
 DECAPx2_ASAP7_75t_R FILLER_15_322 ();
 FILLER_ASAP7_75t_R FILLER_15_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_384 ();
 DECAPx1_ASAP7_75t_R FILLER_15_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_412 ();
 DECAPx10_ASAP7_75t_R FILLER_15_433 ();
 DECAPx1_ASAP7_75t_R FILLER_15_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_516 ();
 FILLER_ASAP7_75t_R FILLER_15_520 ();
 DECAPx4_ASAP7_75t_R FILLER_15_525 ();
 FILLER_ASAP7_75t_R FILLER_15_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_561 ();
 DECAPx6_ASAP7_75t_R FILLER_15_567 ();
 DECAPx2_ASAP7_75t_R FILLER_15_586 ();
 FILLER_ASAP7_75t_R FILLER_15_592 ();
 DECAPx4_ASAP7_75t_R FILLER_15_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_624 ();
 DECAPx10_ASAP7_75t_R FILLER_15_632 ();
 DECAPx10_ASAP7_75t_R FILLER_15_654 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_15_676 ();
 DECAPx6_ASAP7_75t_R FILLER_15_685 ();
 DECAPx1_ASAP7_75t_R FILLER_15_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_703 ();
 FILLER_ASAP7_75t_R FILLER_15_733 ();
 DECAPx10_ASAP7_75t_R FILLER_15_747 ();
 DECAPx2_ASAP7_75t_R FILLER_15_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_775 ();
 DECAPx10_ASAP7_75t_R FILLER_15_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_826 ();
 DECAPx10_ASAP7_75t_R FILLER_15_833 ();
 DECAPx10_ASAP7_75t_R FILLER_15_855 ();
 DECAPx10_ASAP7_75t_R FILLER_15_877 ();
 DECAPx10_ASAP7_75t_R FILLER_15_899 ();
 DECAPx1_ASAP7_75t_R FILLER_15_921 ();
 DECAPx2_ASAP7_75t_R FILLER_15_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_933 ();
 DECAPx10_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_24 ();
 DECAPx10_ASAP7_75t_R FILLER_16_46 ();
 DECAPx10_ASAP7_75t_R FILLER_16_68 ();
 DECAPx10_ASAP7_75t_R FILLER_16_90 ();
 DECAPx2_ASAP7_75t_R FILLER_16_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_118 ();
 DECAPx10_ASAP7_75t_R FILLER_16_147 ();
 DECAPx10_ASAP7_75t_R FILLER_16_169 ();
 DECAPx10_ASAP7_75t_R FILLER_16_191 ();
 DECAPx6_ASAP7_75t_R FILLER_16_213 ();
 DECAPx2_ASAP7_75t_R FILLER_16_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_233 ();
 DECAPx10_ASAP7_75t_R FILLER_16_266 ();
 DECAPx4_ASAP7_75t_R FILLER_16_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_298 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_325 ();
 DECAPx6_ASAP7_75t_R FILLER_16_363 ();
 DECAPx1_ASAP7_75t_R FILLER_16_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_381 ();
 DECAPx10_ASAP7_75t_R FILLER_16_387 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_415 ();
 DECAPx2_ASAP7_75t_R FILLER_16_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_439 ();
 DECAPx6_ASAP7_75t_R FILLER_16_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_459 ();
 DECAPx2_ASAP7_75t_R FILLER_16_464 ();
 FILLER_ASAP7_75t_R FILLER_16_502 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_513 ();
 DECAPx10_ASAP7_75t_R FILLER_16_536 ();
 DECAPx2_ASAP7_75t_R FILLER_16_558 ();
 FILLER_ASAP7_75t_R FILLER_16_581 ();
 DECAPx2_ASAP7_75t_R FILLER_16_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_596 ();
 FILLER_ASAP7_75t_R FILLER_16_604 ();
 DECAPx6_ASAP7_75t_R FILLER_16_618 ();
 DECAPx2_ASAP7_75t_R FILLER_16_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_638 ();
 DECAPx2_ASAP7_75t_R FILLER_16_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_652 ();
 DECAPx10_ASAP7_75t_R FILLER_16_658 ();
 DECAPx6_ASAP7_75t_R FILLER_16_680 ();
 DECAPx1_ASAP7_75t_R FILLER_16_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_698 ();
 DECAPx1_ASAP7_75t_R FILLER_16_713 ();
 DECAPx10_ASAP7_75t_R FILLER_16_729 ();
 DECAPx4_ASAP7_75t_R FILLER_16_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_16_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_776 ();
 DECAPx6_ASAP7_75t_R FILLER_16_794 ();
 DECAPx2_ASAP7_75t_R FILLER_16_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_814 ();
 DECAPx10_ASAP7_75t_R FILLER_16_841 ();
 DECAPx10_ASAP7_75t_R FILLER_16_863 ();
 DECAPx10_ASAP7_75t_R FILLER_16_885 ();
 DECAPx10_ASAP7_75t_R FILLER_16_907 ();
 DECAPx1_ASAP7_75t_R FILLER_16_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_933 ();
 DECAPx10_ASAP7_75t_R FILLER_17_2 ();
 DECAPx10_ASAP7_75t_R FILLER_17_24 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx4_ASAP7_75t_R FILLER_17_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_122 ();
 DECAPx1_ASAP7_75t_R FILLER_17_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_144 ();
 DECAPx6_ASAP7_75t_R FILLER_17_171 ();
 DECAPx2_ASAP7_75t_R FILLER_17_185 ();
 DECAPx6_ASAP7_75t_R FILLER_17_217 ();
 DECAPx2_ASAP7_75t_R FILLER_17_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_237 ();
 DECAPx1_ASAP7_75t_R FILLER_17_244 ();
 DECAPx10_ASAP7_75t_R FILLER_17_251 ();
 DECAPx10_ASAP7_75t_R FILLER_17_273 ();
 DECAPx2_ASAP7_75t_R FILLER_17_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_313 ();
 FILLER_ASAP7_75t_R FILLER_17_342 ();
 DECAPx10_ASAP7_75t_R FILLER_17_352 ();
 FILLER_ASAP7_75t_R FILLER_17_374 ();
 DECAPx10_ASAP7_75t_R FILLER_17_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_421 ();
 DECAPx4_ASAP7_75t_R FILLER_17_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_461 ();
 DECAPx1_ASAP7_75t_R FILLER_17_469 ();
 DECAPx6_ASAP7_75t_R FILLER_17_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_495 ();
 DECAPx2_ASAP7_75t_R FILLER_17_501 ();
 DECAPx10_ASAP7_75t_R FILLER_17_533 ();
 FILLER_ASAP7_75t_R FILLER_17_555 ();
 DECAPx4_ASAP7_75t_R FILLER_17_589 ();
 FILLER_ASAP7_75t_R FILLER_17_599 ();
 FILLER_ASAP7_75t_R FILLER_17_611 ();
 FILLER_ASAP7_75t_R FILLER_17_631 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_17_639 ();
 DECAPx2_ASAP7_75t_R FILLER_17_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_686 ();
 FILLER_ASAP7_75t_R FILLER_17_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_721 ();
 DECAPx10_ASAP7_75t_R FILLER_17_728 ();
 DECAPx4_ASAP7_75t_R FILLER_17_750 ();
 FILLER_ASAP7_75t_R FILLER_17_760 ();
 DECAPx1_ASAP7_75t_R FILLER_17_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_786 ();
 DECAPx10_ASAP7_75t_R FILLER_17_795 ();
 DECAPx2_ASAP7_75t_R FILLER_17_817 ();
 FILLER_ASAP7_75t_R FILLER_17_823 ();
 DECAPx10_ASAP7_75t_R FILLER_17_831 ();
 DECAPx2_ASAP7_75t_R FILLER_17_853 ();
 FILLER_ASAP7_75t_R FILLER_17_859 ();
 DECAPx10_ASAP7_75t_R FILLER_17_867 ();
 DECAPx10_ASAP7_75t_R FILLER_17_889 ();
 DECAPx6_ASAP7_75t_R FILLER_17_911 ();
 DECAPx2_ASAP7_75t_R FILLER_17_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_933 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx6_ASAP7_75t_R FILLER_18_112 ();
 DECAPx2_ASAP7_75t_R FILLER_18_126 ();
 DECAPx1_ASAP7_75t_R FILLER_18_144 ();
 FILLER_ASAP7_75t_R FILLER_18_154 ();
 FILLER_ASAP7_75t_R FILLER_18_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_170 ();
 DECAPx1_ASAP7_75t_R FILLER_18_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_196 ();
 DECAPx10_ASAP7_75t_R FILLER_18_231 ();
 DECAPx4_ASAP7_75t_R FILLER_18_253 ();
 FILLER_ASAP7_75t_R FILLER_18_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_271 ();
 DECAPx6_ASAP7_75t_R FILLER_18_300 ();
 DECAPx1_ASAP7_75t_R FILLER_18_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_321 ();
 FILLER_ASAP7_75t_R FILLER_18_328 ();
 DECAPx10_ASAP7_75t_R FILLER_18_333 ();
 DECAPx4_ASAP7_75t_R FILLER_18_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_371 ();
 DECAPx1_ASAP7_75t_R FILLER_18_392 ();
 DECAPx2_ASAP7_75t_R FILLER_18_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_433 ();
 FILLER_ASAP7_75t_R FILLER_18_439 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_459 ();
 DECAPx1_ASAP7_75t_R FILLER_18_464 ();
 DECAPx10_ASAP7_75t_R FILLER_18_498 ();
 DECAPx2_ASAP7_75t_R FILLER_18_520 ();
 DECAPx2_ASAP7_75t_R FILLER_18_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_540 ();
 DECAPx6_ASAP7_75t_R FILLER_18_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_591 ();
 DECAPx1_ASAP7_75t_R FILLER_18_609 ();
 DECAPx6_ASAP7_75t_R FILLER_18_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_659 ();
 DECAPx1_ASAP7_75t_R FILLER_18_665 ();
 DECAPx1_ASAP7_75t_R FILLER_18_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_676 ();
 FILLER_ASAP7_75t_R FILLER_18_705 ();
 DECAPx6_ASAP7_75t_R FILLER_18_713 ();
 DECAPx1_ASAP7_75t_R FILLER_18_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_731 ();
 DECAPx4_ASAP7_75t_R FILLER_18_740 ();
 FILLER_ASAP7_75t_R FILLER_18_750 ();
 DECAPx2_ASAP7_75t_R FILLER_18_759 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_18_765 ();
 FILLER_ASAP7_75t_R FILLER_18_780 ();
 DECAPx10_ASAP7_75t_R FILLER_18_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_810 ();
 DECAPx6_ASAP7_75t_R FILLER_18_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_835 ();
 DECAPx10_ASAP7_75t_R FILLER_18_876 ();
 DECAPx10_ASAP7_75t_R FILLER_18_898 ();
 DECAPx6_ASAP7_75t_R FILLER_18_920 ();
 DECAPx10_ASAP7_75t_R FILLER_19_2 ();
 DECAPx10_ASAP7_75t_R FILLER_19_24 ();
 DECAPx10_ASAP7_75t_R FILLER_19_46 ();
 DECAPx10_ASAP7_75t_R FILLER_19_68 ();
 DECAPx6_ASAP7_75t_R FILLER_19_90 ();
 DECAPx2_ASAP7_75t_R FILLER_19_104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_136 ();
 DECAPx1_ASAP7_75t_R FILLER_19_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_191 ();
 DECAPx2_ASAP7_75t_R FILLER_19_217 ();
 FILLER_ASAP7_75t_R FILLER_19_229 ();
 DECAPx2_ASAP7_75t_R FILLER_19_237 ();
 DECAPx1_ASAP7_75t_R FILLER_19_255 ();
 DECAPx1_ASAP7_75t_R FILLER_19_265 ();
 DECAPx1_ASAP7_75t_R FILLER_19_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_311 ();
 DECAPx4_ASAP7_75t_R FILLER_19_324 ();
 DECAPx6_ASAP7_75t_R FILLER_19_340 ();
 DECAPx2_ASAP7_75t_R FILLER_19_354 ();
 DECAPx6_ASAP7_75t_R FILLER_19_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_380 ();
 FILLER_ASAP7_75t_R FILLER_19_387 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_429 ();
 DECAPx2_ASAP7_75t_R FILLER_19_438 ();
 DECAPx1_ASAP7_75t_R FILLER_19_452 ();
 DECAPx10_ASAP7_75t_R FILLER_19_462 ();
 DECAPx1_ASAP7_75t_R FILLER_19_484 ();
 DECAPx6_ASAP7_75t_R FILLER_19_500 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_19_514 ();
 DECAPx6_ASAP7_75t_R FILLER_19_523 ();
 DECAPx1_ASAP7_75t_R FILLER_19_537 ();
 DECAPx6_ASAP7_75t_R FILLER_19_567 ();
 FILLER_ASAP7_75t_R FILLER_19_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_591 ();
 DECAPx1_ASAP7_75t_R FILLER_19_615 ();
 DECAPx1_ASAP7_75t_R FILLER_19_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_626 ();
 DECAPx6_ASAP7_75t_R FILLER_19_635 ();
 DECAPx2_ASAP7_75t_R FILLER_19_649 ();
 DECAPx1_ASAP7_75t_R FILLER_19_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_685 ();
 DECAPx1_ASAP7_75t_R FILLER_19_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_726 ();
 DECAPx10_ASAP7_75t_R FILLER_19_767 ();
 DECAPx1_ASAP7_75t_R FILLER_19_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_793 ();
 DECAPx10_ASAP7_75t_R FILLER_19_808 ();
 DECAPx1_ASAP7_75t_R FILLER_19_830 ();
 DECAPx10_ASAP7_75t_R FILLER_19_867 ();
 DECAPx10_ASAP7_75t_R FILLER_19_889 ();
 DECAPx6_ASAP7_75t_R FILLER_19_911 ();
 DECAPx2_ASAP7_75t_R FILLER_19_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_933 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_112 ();
 DECAPx1_ASAP7_75t_R FILLER_20_174 ();
 DECAPx10_ASAP7_75t_R FILLER_20_191 ();
 DECAPx10_ASAP7_75t_R FILLER_20_213 ();
 FILLER_ASAP7_75t_R FILLER_20_235 ();
 DECAPx2_ASAP7_75t_R FILLER_20_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_284 ();
 DECAPx6_ASAP7_75t_R FILLER_20_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_310 ();
 DECAPx2_ASAP7_75t_R FILLER_20_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_354 ();
 DECAPx1_ASAP7_75t_R FILLER_20_363 ();
 DECAPx2_ASAP7_75t_R FILLER_20_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_401 ();
 FILLER_ASAP7_75t_R FILLER_20_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_433 ();
 DECAPx4_ASAP7_75t_R FILLER_20_452 ();
 DECAPx6_ASAP7_75t_R FILLER_20_464 ();
 DECAPx1_ASAP7_75t_R FILLER_20_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_482 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_503 ();
 FILLER_ASAP7_75t_R FILLER_20_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_528 ();
 DECAPx6_ASAP7_75t_R FILLER_20_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_555 ();
 DECAPx2_ASAP7_75t_R FILLER_20_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_568 ();
 DECAPx2_ASAP7_75t_R FILLER_20_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_587 ();
 DECAPx1_ASAP7_75t_R FILLER_20_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_598 ();
 DECAPx6_ASAP7_75t_R FILLER_20_604 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_618 ();
 DECAPx1_ASAP7_75t_R FILLER_20_672 ();
 DECAPx10_ASAP7_75t_R FILLER_20_682 ();
 DECAPx2_ASAP7_75t_R FILLER_20_704 ();
 DECAPx6_ASAP7_75t_R FILLER_20_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_732 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_20_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_756 ();
 DECAPx6_ASAP7_75t_R FILLER_20_763 ();
 DECAPx1_ASAP7_75t_R FILLER_20_777 ();
 DECAPx1_ASAP7_75t_R FILLER_20_787 ();
 FILLER_ASAP7_75t_R FILLER_20_811 ();
 DECAPx10_ASAP7_75t_R FILLER_20_820 ();
 DECAPx10_ASAP7_75t_R FILLER_20_842 ();
 DECAPx10_ASAP7_75t_R FILLER_20_864 ();
 DECAPx10_ASAP7_75t_R FILLER_20_886 ();
 DECAPx10_ASAP7_75t_R FILLER_20_908 ();
 DECAPx1_ASAP7_75t_R FILLER_20_930 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx4_ASAP7_75t_R FILLER_21_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_122 ();
 DECAPx2_ASAP7_75t_R FILLER_21_143 ();
 FILLER_ASAP7_75t_R FILLER_21_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_157 ();
 DECAPx2_ASAP7_75t_R FILLER_21_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_170 ();
 DECAPx10_ASAP7_75t_R FILLER_21_192 ();
 DECAPx10_ASAP7_75t_R FILLER_21_214 ();
 DECAPx6_ASAP7_75t_R FILLER_21_236 ();
 FILLER_ASAP7_75t_R FILLER_21_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_264 ();
 DECAPx10_ASAP7_75t_R FILLER_21_271 ();
 DECAPx10_ASAP7_75t_R FILLER_21_293 ();
 DECAPx6_ASAP7_75t_R FILLER_21_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_335 ();
 DECAPx4_ASAP7_75t_R FILLER_21_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_392 ();
 DECAPx6_ASAP7_75t_R FILLER_21_400 ();
 DECAPx2_ASAP7_75t_R FILLER_21_414 ();
 FILLER_ASAP7_75t_R FILLER_21_426 ();
 DECAPx6_ASAP7_75t_R FILLER_21_438 ();
 FILLER_ASAP7_75t_R FILLER_21_452 ();
 DECAPx1_ASAP7_75t_R FILLER_21_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_463 ();
 DECAPx1_ASAP7_75t_R FILLER_21_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_473 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_497 ();
 DECAPx2_ASAP7_75t_R FILLER_21_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_514 ();
 FILLER_ASAP7_75t_R FILLER_21_529 ();
 DECAPx10_ASAP7_75t_R FILLER_21_537 ();
 DECAPx2_ASAP7_75t_R FILLER_21_559 ();
 FILLER_ASAP7_75t_R FILLER_21_565 ();
 DECAPx10_ASAP7_75t_R FILLER_21_575 ();
 DECAPx10_ASAP7_75t_R FILLER_21_597 ();
 DECAPx4_ASAP7_75t_R FILLER_21_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_629 ();
 DECAPx2_ASAP7_75t_R FILLER_21_636 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_642 ();
 DECAPx1_ASAP7_75t_R FILLER_21_671 ();
 DECAPx6_ASAP7_75t_R FILLER_21_701 ();
 DECAPx1_ASAP7_75t_R FILLER_21_715 ();
 DECAPx10_ASAP7_75t_R FILLER_21_725 ();
 DECAPx6_ASAP7_75t_R FILLER_21_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_761 ();
 DECAPx2_ASAP7_75t_R FILLER_21_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_21_782 ();
 DECAPx2_ASAP7_75t_R FILLER_21_791 ();
 FILLER_ASAP7_75t_R FILLER_21_797 ();
 FILLER_ASAP7_75t_R FILLER_21_807 ();
 DECAPx1_ASAP7_75t_R FILLER_21_829 ();
 DECAPx2_ASAP7_75t_R FILLER_21_842 ();
 DECAPx1_ASAP7_75t_R FILLER_21_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_858 ();
 DECAPx10_ASAP7_75t_R FILLER_21_867 ();
 DECAPx10_ASAP7_75t_R FILLER_21_889 ();
 DECAPx6_ASAP7_75t_R FILLER_21_911 ();
 DECAPx2_ASAP7_75t_R FILLER_21_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_933 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx10_ASAP7_75t_R FILLER_22_134 ();
 DECAPx10_ASAP7_75t_R FILLER_22_156 ();
 DECAPx6_ASAP7_75t_R FILLER_22_185 ();
 DECAPx2_ASAP7_75t_R FILLER_22_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_205 ();
 FILLER_ASAP7_75t_R FILLER_22_232 ();
 DECAPx6_ASAP7_75t_R FILLER_22_246 ();
 FILLER_ASAP7_75t_R FILLER_22_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_270 ();
 DECAPx10_ASAP7_75t_R FILLER_22_277 ();
 DECAPx10_ASAP7_75t_R FILLER_22_299 ();
 DECAPx10_ASAP7_75t_R FILLER_22_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_343 ();
 FILLER_ASAP7_75t_R FILLER_22_364 ();
 FILLER_ASAP7_75t_R FILLER_22_372 ();
 DECAPx10_ASAP7_75t_R FILLER_22_402 ();
 DECAPx4_ASAP7_75t_R FILLER_22_424 ();
 DECAPx2_ASAP7_75t_R FILLER_22_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_450 ();
 DECAPx2_ASAP7_75t_R FILLER_22_456 ();
 DECAPx10_ASAP7_75t_R FILLER_22_476 ();
 FILLER_ASAP7_75t_R FILLER_22_504 ();
 DECAPx10_ASAP7_75t_R FILLER_22_514 ();
 DECAPx4_ASAP7_75t_R FILLER_22_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_552 ();
 DECAPx4_ASAP7_75t_R FILLER_22_587 ();
 FILLER_ASAP7_75t_R FILLER_22_597 ();
 DECAPx6_ASAP7_75t_R FILLER_22_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_630 ();
 DECAPx6_ASAP7_75t_R FILLER_22_637 ();
 DECAPx1_ASAP7_75t_R FILLER_22_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_655 ();
 DECAPx4_ASAP7_75t_R FILLER_22_662 ();
 FILLER_ASAP7_75t_R FILLER_22_672 ();
 DECAPx1_ASAP7_75t_R FILLER_22_685 ();
 DECAPx4_ASAP7_75t_R FILLER_22_692 ();
 FILLER_ASAP7_75t_R FILLER_22_702 ();
 FILLER_ASAP7_75t_R FILLER_22_721 ();
 DECAPx10_ASAP7_75t_R FILLER_22_746 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_768 ();
 FILLER_ASAP7_75t_R FILLER_22_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_785 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_874 ();
 DECAPx10_ASAP7_75t_R FILLER_22_881 ();
 DECAPx10_ASAP7_75t_R FILLER_22_903 ();
 DECAPx2_ASAP7_75t_R FILLER_22_925 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_22_931 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx4_ASAP7_75t_R FILLER_23_134 ();
 FILLER_ASAP7_75t_R FILLER_23_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_152 ();
 DECAPx2_ASAP7_75t_R FILLER_23_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_165 ();
 DECAPx1_ASAP7_75t_R FILLER_23_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_188 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_195 ();
 DECAPx10_ASAP7_75t_R FILLER_23_256 ();
 FILLER_ASAP7_75t_R FILLER_23_278 ();
 DECAPx1_ASAP7_75t_R FILLER_23_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_299 ();
 FILLER_ASAP7_75t_R FILLER_23_320 ();
 DECAPx10_ASAP7_75t_R FILLER_23_325 ();
 DECAPx2_ASAP7_75t_R FILLER_23_347 ();
 FILLER_ASAP7_75t_R FILLER_23_353 ();
 DECAPx1_ASAP7_75t_R FILLER_23_367 ();
 FILLER_ASAP7_75t_R FILLER_23_391 ();
 DECAPx10_ASAP7_75t_R FILLER_23_407 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_488 ();
 DECAPx10_ASAP7_75t_R FILLER_23_495 ();
 DECAPx10_ASAP7_75t_R FILLER_23_517 ();
 DECAPx2_ASAP7_75t_R FILLER_23_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_595 ();
 DECAPx1_ASAP7_75t_R FILLER_23_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_638 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_657 ();
 FILLER_ASAP7_75t_R FILLER_23_673 ();
 DECAPx4_ASAP7_75t_R FILLER_23_681 ();
 DECAPx4_ASAP7_75t_R FILLER_23_694 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_781 ();
 DECAPx10_ASAP7_75t_R FILLER_23_796 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_23_818 ();
 DECAPx1_ASAP7_75t_R FILLER_23_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_831 ();
 DECAPx6_ASAP7_75t_R FILLER_23_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_860 ();
 DECAPx10_ASAP7_75t_R FILLER_23_901 ();
 FILLER_ASAP7_75t_R FILLER_23_923 ();
 DECAPx2_ASAP7_75t_R FILLER_23_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_933 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx2_ASAP7_75t_R FILLER_24_112 ();
 FILLER_ASAP7_75t_R FILLER_24_124 ();
 DECAPx4_ASAP7_75t_R FILLER_24_132 ();
 FILLER_ASAP7_75t_R FILLER_24_149 ();
 DECAPx1_ASAP7_75t_R FILLER_24_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_209 ();
 DECAPx1_ASAP7_75t_R FILLER_24_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_230 ();
 DECAPx1_ASAP7_75t_R FILLER_24_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_241 ();
 DECAPx10_ASAP7_75t_R FILLER_24_245 ();
 DECAPx2_ASAP7_75t_R FILLER_24_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_273 ();
 DECAPx2_ASAP7_75t_R FILLER_24_309 ();
 FILLER_ASAP7_75t_R FILLER_24_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_343 ();
 DECAPx10_ASAP7_75t_R FILLER_24_352 ();
 DECAPx1_ASAP7_75t_R FILLER_24_374 ();
 FILLER_ASAP7_75t_R FILLER_24_384 ();
 DECAPx1_ASAP7_75t_R FILLER_24_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_470 ();
 DECAPx4_ASAP7_75t_R FILLER_24_478 ();
 DECAPx4_ASAP7_75t_R FILLER_24_500 ();
 DECAPx4_ASAP7_75t_R FILLER_24_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_523 ();
 DECAPx2_ASAP7_75t_R FILLER_24_539 ();
 DECAPx1_ASAP7_75t_R FILLER_24_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_557 ();
 DECAPx1_ASAP7_75t_R FILLER_24_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_700 ();
 DECAPx2_ASAP7_75t_R FILLER_24_720 ();
 DECAPx1_ASAP7_75t_R FILLER_24_742 ();
 DECAPx10_ASAP7_75t_R FILLER_24_766 ();
 DECAPx10_ASAP7_75t_R FILLER_24_788 ();
 DECAPx10_ASAP7_75t_R FILLER_24_810 ();
 DECAPx10_ASAP7_75t_R FILLER_24_832 ();
 DECAPx6_ASAP7_75t_R FILLER_24_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_24_868 ();
 DECAPx1_ASAP7_75t_R FILLER_24_877 ();
 DECAPx10_ASAP7_75t_R FILLER_24_907 ();
 DECAPx1_ASAP7_75t_R FILLER_24_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_933 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx6_ASAP7_75t_R FILLER_25_90 ();
 DECAPx1_ASAP7_75t_R FILLER_25_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_108 ();
 DECAPx1_ASAP7_75t_R FILLER_25_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_139 ();
 DECAPx2_ASAP7_75t_R FILLER_25_166 ();
 FILLER_ASAP7_75t_R FILLER_25_178 ();
 FILLER_ASAP7_75t_R FILLER_25_186 ();
 DECAPx10_ASAP7_75t_R FILLER_25_208 ();
 DECAPx6_ASAP7_75t_R FILLER_25_230 ();
 FILLER_ASAP7_75t_R FILLER_25_244 ();
 DECAPx2_ASAP7_75t_R FILLER_25_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_265 ();
 DECAPx2_ASAP7_75t_R FILLER_25_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_277 ();
 FILLER_ASAP7_75t_R FILLER_25_284 ();
 DECAPx2_ASAP7_75t_R FILLER_25_312 ();
 FILLER_ASAP7_75t_R FILLER_25_318 ();
 FILLER_ASAP7_75t_R FILLER_25_326 ();
 DECAPx6_ASAP7_75t_R FILLER_25_368 ();
 DECAPx1_ASAP7_75t_R FILLER_25_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_386 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_392 ();
 DECAPx2_ASAP7_75t_R FILLER_25_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_412 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_436 ();
 DECAPx10_ASAP7_75t_R FILLER_25_459 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_501 ();
 FILLER_ASAP7_75t_R FILLER_25_516 ();
 DECAPx10_ASAP7_75t_R FILLER_25_524 ();
 DECAPx2_ASAP7_75t_R FILLER_25_546 ();
 DECAPx2_ASAP7_75t_R FILLER_25_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_575 ();
 DECAPx1_ASAP7_75t_R FILLER_25_581 ();
 FILLER_ASAP7_75t_R FILLER_25_599 ();
 DECAPx10_ASAP7_75t_R FILLER_25_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_628 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_648 ();
 DECAPx10_ASAP7_75t_R FILLER_25_700 ();
 DECAPx10_ASAP7_75t_R FILLER_25_722 ();
 DECAPx10_ASAP7_75t_R FILLER_25_765 ();
 DECAPx1_ASAP7_75t_R FILLER_25_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_25_803 ();
 DECAPx6_ASAP7_75t_R FILLER_25_818 ();
 DECAPx1_ASAP7_75t_R FILLER_25_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_836 ();
 DECAPx10_ASAP7_75t_R FILLER_25_845 ();
 DECAPx10_ASAP7_75t_R FILLER_25_867 ();
 DECAPx1_ASAP7_75t_R FILLER_25_889 ();
 DECAPx6_ASAP7_75t_R FILLER_25_906 ();
 DECAPx1_ASAP7_75t_R FILLER_25_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_924 ();
 DECAPx2_ASAP7_75t_R FILLER_25_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_933 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 FILLER_ASAP7_75t_R FILLER_26_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_137 ();
 DECAPx4_ASAP7_75t_R FILLER_26_144 ();
 DECAPx2_ASAP7_75t_R FILLER_26_163 ();
 DECAPx6_ASAP7_75t_R FILLER_26_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_209 ();
 DECAPx10_ASAP7_75t_R FILLER_26_216 ();
 FILLER_ASAP7_75t_R FILLER_26_238 ();
 DECAPx1_ASAP7_75t_R FILLER_26_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_252 ();
 DECAPx2_ASAP7_75t_R FILLER_26_282 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_288 ();
 DECAPx1_ASAP7_75t_R FILLER_26_297 ();
 DECAPx1_ASAP7_75t_R FILLER_26_304 ();
 DECAPx10_ASAP7_75t_R FILLER_26_314 ();
 DECAPx2_ASAP7_75t_R FILLER_26_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_342 ();
 DECAPx1_ASAP7_75t_R FILLER_26_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_353 ();
 DECAPx4_ASAP7_75t_R FILLER_26_357 ();
 FILLER_ASAP7_75t_R FILLER_26_367 ();
 DECAPx2_ASAP7_75t_R FILLER_26_375 ();
 DECAPx10_ASAP7_75t_R FILLER_26_399 ();
 DECAPx6_ASAP7_75t_R FILLER_26_421 ();
 DECAPx2_ASAP7_75t_R FILLER_26_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_441 ();
 DECAPx6_ASAP7_75t_R FILLER_26_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_461 ();
 DECAPx1_ASAP7_75t_R FILLER_26_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_468 ();
 DECAPx4_ASAP7_75t_R FILLER_26_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_491 ();
 DECAPx4_ASAP7_75t_R FILLER_26_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_508 ();
 DECAPx10_ASAP7_75t_R FILLER_26_530 ();
 DECAPx1_ASAP7_75t_R FILLER_26_552 ();
 DECAPx10_ASAP7_75t_R FILLER_26_564 ();
 DECAPx6_ASAP7_75t_R FILLER_26_586 ();
 DECAPx1_ASAP7_75t_R FILLER_26_600 ();
 FILLER_ASAP7_75t_R FILLER_26_611 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_619 ();
 DECAPx4_ASAP7_75t_R FILLER_26_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_638 ();
 DECAPx2_ASAP7_75t_R FILLER_26_648 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_681 ();
 DECAPx10_ASAP7_75t_R FILLER_26_708 ();
 DECAPx10_ASAP7_75t_R FILLER_26_730 ();
 DECAPx4_ASAP7_75t_R FILLER_26_752 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_762 ();
 DECAPx6_ASAP7_75t_R FILLER_26_774 ();
 DECAPx2_ASAP7_75t_R FILLER_26_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_794 ();
 DECAPx6_ASAP7_75t_R FILLER_26_822 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_843 ();
 DECAPx10_ASAP7_75t_R FILLER_26_855 ();
 DECAPx10_ASAP7_75t_R FILLER_26_877 ();
 DECAPx10_ASAP7_75t_R FILLER_26_899 ();
 DECAPx4_ASAP7_75t_R FILLER_26_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_26_931 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx6_ASAP7_75t_R FILLER_27_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_126 ();
 DECAPx1_ASAP7_75t_R FILLER_27_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_147 ();
 DECAPx10_ASAP7_75t_R FILLER_27_155 ();
 DECAPx2_ASAP7_75t_R FILLER_27_177 ();
 DECAPx6_ASAP7_75t_R FILLER_27_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_200 ();
 DECAPx1_ASAP7_75t_R FILLER_27_230 ();
 DECAPx10_ASAP7_75t_R FILLER_27_266 ();
 DECAPx10_ASAP7_75t_R FILLER_27_288 ();
 DECAPx10_ASAP7_75t_R FILLER_27_310 ();
 DECAPx10_ASAP7_75t_R FILLER_27_332 ();
 DECAPx1_ASAP7_75t_R FILLER_27_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_358 ();
 DECAPx1_ASAP7_75t_R FILLER_27_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_402 ();
 DECAPx1_ASAP7_75t_R FILLER_27_409 ();
 DECAPx10_ASAP7_75t_R FILLER_27_436 ();
 DECAPx6_ASAP7_75t_R FILLER_27_458 ();
 DECAPx10_ASAP7_75t_R FILLER_27_484 ();
 DECAPx10_ASAP7_75t_R FILLER_27_506 ();
 DECAPx2_ASAP7_75t_R FILLER_27_528 ();
 DECAPx4_ASAP7_75t_R FILLER_27_541 ();
 DECAPx6_ASAP7_75t_R FILLER_27_580 ();
 DECAPx2_ASAP7_75t_R FILLER_27_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_600 ();
 DECAPx1_ASAP7_75t_R FILLER_27_621 ();
 DECAPx10_ASAP7_75t_R FILLER_27_632 ();
 DECAPx6_ASAP7_75t_R FILLER_27_654 ();
 FILLER_ASAP7_75t_R FILLER_27_673 ();
 FILLER_ASAP7_75t_R FILLER_27_690 ();
 DECAPx1_ASAP7_75t_R FILLER_27_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_704 ();
 FILLER_ASAP7_75t_R FILLER_27_723 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_737 ();
 DECAPx6_ASAP7_75t_R FILLER_27_747 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_761 ();
 DECAPx6_ASAP7_75t_R FILLER_27_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_798 ();
 DECAPx4_ASAP7_75t_R FILLER_27_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_838 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_27_877 ();
 DECAPx10_ASAP7_75t_R FILLER_27_893 ();
 DECAPx4_ASAP7_75t_R FILLER_27_915 ();
 FILLER_ASAP7_75t_R FILLER_27_927 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx6_ASAP7_75t_R FILLER_28_90 ();
 DECAPx1_ASAP7_75t_R FILLER_28_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_108 ();
 DECAPx10_ASAP7_75t_R FILLER_28_130 ();
 DECAPx10_ASAP7_75t_R FILLER_28_152 ();
 DECAPx10_ASAP7_75t_R FILLER_28_174 ();
 DECAPx4_ASAP7_75t_R FILLER_28_196 ();
 DECAPx1_ASAP7_75t_R FILLER_28_212 ();
 DECAPx10_ASAP7_75t_R FILLER_28_251 ();
 DECAPx10_ASAP7_75t_R FILLER_28_273 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_295 ();
 DECAPx1_ASAP7_75t_R FILLER_28_310 ();
 DECAPx1_ASAP7_75t_R FILLER_28_326 ();
 DECAPx1_ASAP7_75t_R FILLER_28_336 ();
 FILLER_ASAP7_75t_R FILLER_28_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_405 ();
 DECAPx6_ASAP7_75t_R FILLER_28_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_435 ();
 DECAPx2_ASAP7_75t_R FILLER_28_454 ();
 FILLER_ASAP7_75t_R FILLER_28_460 ();
 DECAPx4_ASAP7_75t_R FILLER_28_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_474 ();
 DECAPx4_ASAP7_75t_R FILLER_28_506 ();
 DECAPx4_ASAP7_75t_R FILLER_28_522 ();
 DECAPx4_ASAP7_75t_R FILLER_28_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_556 ();
 DECAPx1_ASAP7_75t_R FILLER_28_579 ();
 DECAPx4_ASAP7_75t_R FILLER_28_595 ();
 FILLER_ASAP7_75t_R FILLER_28_605 ();
 DECAPx2_ASAP7_75t_R FILLER_28_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_624 ();
 DECAPx4_ASAP7_75t_R FILLER_28_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_643 ();
 DECAPx6_ASAP7_75t_R FILLER_28_650 ();
 DECAPx1_ASAP7_75t_R FILLER_28_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_668 ();
 DECAPx4_ASAP7_75t_R FILLER_28_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_697 ();
 DECAPx4_ASAP7_75t_R FILLER_28_750 ();
 FILLER_ASAP7_75t_R FILLER_28_760 ();
 DECAPx10_ASAP7_75t_R FILLER_28_790 ();
 DECAPx4_ASAP7_75t_R FILLER_28_812 ();
 DECAPx2_ASAP7_75t_R FILLER_28_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_853 ();
 FILLER_ASAP7_75t_R FILLER_28_862 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_872 ();
 DECAPx10_ASAP7_75t_R FILLER_28_895 ();
 DECAPx6_ASAP7_75t_R FILLER_28_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_28_931 ();
 DECAPx10_ASAP7_75t_R FILLER_29_2 ();
 DECAPx10_ASAP7_75t_R FILLER_29_24 ();
 DECAPx10_ASAP7_75t_R FILLER_29_46 ();
 DECAPx10_ASAP7_75t_R FILLER_29_68 ();
 DECAPx6_ASAP7_75t_R FILLER_29_90 ();
 DECAPx1_ASAP7_75t_R FILLER_29_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_108 ();
 DECAPx6_ASAP7_75t_R FILLER_29_138 ();
 FILLER_ASAP7_75t_R FILLER_29_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_163 ();
 DECAPx10_ASAP7_75t_R FILLER_29_182 ();
 DECAPx10_ASAP7_75t_R FILLER_29_204 ();
 DECAPx2_ASAP7_75t_R FILLER_29_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_239 ();
 DECAPx6_ASAP7_75t_R FILLER_29_243 ();
 FILLER_ASAP7_75t_R FILLER_29_257 ();
 DECAPx1_ASAP7_75t_R FILLER_29_285 ();
 DECAPx10_ASAP7_75t_R FILLER_29_321 ();
 DECAPx1_ASAP7_75t_R FILLER_29_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_347 ();
 DECAPx4_ASAP7_75t_R FILLER_29_366 ();
 FILLER_ASAP7_75t_R FILLER_29_376 ();
 DECAPx1_ASAP7_75t_R FILLER_29_410 ();
 DECAPx4_ASAP7_75t_R FILLER_29_420 ();
 DECAPx1_ASAP7_75t_R FILLER_29_458 ();
 DECAPx1_ASAP7_75t_R FILLER_29_470 ();
 DECAPx6_ASAP7_75t_R FILLER_29_480 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_504 ();
 DECAPx1_ASAP7_75t_R FILLER_29_520 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_538 ();
 FILLER_ASAP7_75t_R FILLER_29_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_609 ();
 DECAPx1_ASAP7_75t_R FILLER_29_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_643 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_29_670 ();
 DECAPx2_ASAP7_75t_R FILLER_29_699 ();
 FILLER_ASAP7_75t_R FILLER_29_705 ();
 FILLER_ASAP7_75t_R FILLER_29_714 ();
 DECAPx1_ASAP7_75t_R FILLER_29_728 ();
 DECAPx2_ASAP7_75t_R FILLER_29_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_751 ();
 DECAPx4_ASAP7_75t_R FILLER_29_764 ();
 FILLER_ASAP7_75t_R FILLER_29_774 ();
 DECAPx2_ASAP7_75t_R FILLER_29_782 ();
 DECAPx10_ASAP7_75t_R FILLER_29_800 ();
 DECAPx10_ASAP7_75t_R FILLER_29_822 ();
 DECAPx10_ASAP7_75t_R FILLER_29_844 ();
 DECAPx4_ASAP7_75t_R FILLER_29_866 ();
 DECAPx10_ASAP7_75t_R FILLER_29_888 ();
 DECAPx6_ASAP7_75t_R FILLER_29_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_924 ();
 DECAPx2_ASAP7_75t_R FILLER_29_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_29_933 ();
 DECAPx10_ASAP7_75t_R FILLER_30_2 ();
 DECAPx10_ASAP7_75t_R FILLER_30_24 ();
 DECAPx10_ASAP7_75t_R FILLER_30_46 ();
 DECAPx10_ASAP7_75t_R FILLER_30_68 ();
 DECAPx10_ASAP7_75t_R FILLER_30_90 ();
 DECAPx2_ASAP7_75t_R FILLER_30_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_118 ();
 DECAPx6_ASAP7_75t_R FILLER_30_128 ();
 FILLER_ASAP7_75t_R FILLER_30_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_150 ();
 FILLER_ASAP7_75t_R FILLER_30_159 ();
 DECAPx1_ASAP7_75t_R FILLER_30_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_215 ();
 DECAPx10_ASAP7_75t_R FILLER_30_229 ();
 DECAPx4_ASAP7_75t_R FILLER_30_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_261 ();
 FILLER_ASAP7_75t_R FILLER_30_269 ();
 FILLER_ASAP7_75t_R FILLER_30_291 ();
 DECAPx2_ASAP7_75t_R FILLER_30_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_318 ();
 DECAPx10_ASAP7_75t_R FILLER_30_347 ();
 FILLER_ASAP7_75t_R FILLER_30_369 ();
 DECAPx10_ASAP7_75t_R FILLER_30_374 ();
 DECAPx6_ASAP7_75t_R FILLER_30_396 ();
 DECAPx1_ASAP7_75t_R FILLER_30_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_476 ();
 DECAPx4_ASAP7_75t_R FILLER_30_483 ();
 DECAPx1_ASAP7_75t_R FILLER_30_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_515 ();
 DECAPx6_ASAP7_75t_R FILLER_30_552 ();
 FILLER_ASAP7_75t_R FILLER_30_571 ();
 DECAPx2_ASAP7_75t_R FILLER_30_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_589 ();
 DECAPx10_ASAP7_75t_R FILLER_30_593 ();
 DECAPx6_ASAP7_75t_R FILLER_30_615 ();
 FILLER_ASAP7_75t_R FILLER_30_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_637 ();
 DECAPx4_ASAP7_75t_R FILLER_30_666 ();
 DECAPx10_ASAP7_75t_R FILLER_30_692 ();
 DECAPx10_ASAP7_75t_R FILLER_30_714 ();
 DECAPx6_ASAP7_75t_R FILLER_30_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_750 ();
 DECAPx10_ASAP7_75t_R FILLER_30_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_791 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_811 ();
 DECAPx1_ASAP7_75t_R FILLER_30_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_830 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_30_846 ();
 DECAPx10_ASAP7_75t_R FILLER_30_862 ();
 DECAPx4_ASAP7_75t_R FILLER_30_884 ();
 DECAPx10_ASAP7_75t_R FILLER_30_907 ();
 DECAPx1_ASAP7_75t_R FILLER_30_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_30_933 ();
 DECAPx10_ASAP7_75t_R FILLER_31_2 ();
 DECAPx10_ASAP7_75t_R FILLER_31_24 ();
 DECAPx10_ASAP7_75t_R FILLER_31_46 ();
 DECAPx10_ASAP7_75t_R FILLER_31_68 ();
 DECAPx10_ASAP7_75t_R FILLER_31_90 ();
 DECAPx6_ASAP7_75t_R FILLER_31_112 ();
 DECAPx1_ASAP7_75t_R FILLER_31_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_130 ();
 DECAPx1_ASAP7_75t_R FILLER_31_209 ();
 DECAPx6_ASAP7_75t_R FILLER_31_245 ();
 FILLER_ASAP7_75t_R FILLER_31_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_267 ();
 FILLER_ASAP7_75t_R FILLER_31_277 ();
 DECAPx6_ASAP7_75t_R FILLER_31_287 ();
 DECAPx1_ASAP7_75t_R FILLER_31_330 ();
 DECAPx4_ASAP7_75t_R FILLER_31_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_358 ();
 DECAPx4_ASAP7_75t_R FILLER_31_381 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_391 ();
 DECAPx10_ASAP7_75t_R FILLER_31_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_421 ();
 DECAPx2_ASAP7_75t_R FILLER_31_430 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_448 ();
 DECAPx2_ASAP7_75t_R FILLER_31_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_489 ();
 DECAPx1_ASAP7_75t_R FILLER_31_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_508 ();
 DECAPx6_ASAP7_75t_R FILLER_31_515 ();
 DECAPx10_ASAP7_75t_R FILLER_31_545 ();
 DECAPx1_ASAP7_75t_R FILLER_31_575 ();
 DECAPx2_ASAP7_75t_R FILLER_31_594 ();
 FILLER_ASAP7_75t_R FILLER_31_600 ();
 DECAPx2_ASAP7_75t_R FILLER_31_605 ();
 DECAPx6_ASAP7_75t_R FILLER_31_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_666 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_678 ();
 DECAPx1_ASAP7_75t_R FILLER_31_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_698 ();
 DECAPx6_ASAP7_75t_R FILLER_31_707 ();
 DECAPx1_ASAP7_75t_R FILLER_31_721 ();
 DECAPx1_ASAP7_75t_R FILLER_31_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_756 ();
 DECAPx2_ASAP7_75t_R FILLER_31_777 ();
 DECAPx1_ASAP7_75t_R FILLER_31_789 ();
 DECAPx4_ASAP7_75t_R FILLER_31_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_829 ();
 DECAPx2_ASAP7_75t_R FILLER_31_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_31_842 ();
 FILLER_ASAP7_75t_R FILLER_31_863 ();
 DECAPx6_ASAP7_75t_R FILLER_31_871 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_885 ();
 DECAPx6_ASAP7_75t_R FILLER_31_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_31_922 ();
 FILLER_ASAP7_75t_R FILLER_31_927 ();
 DECAPx10_ASAP7_75t_R FILLER_32_2 ();
 DECAPx10_ASAP7_75t_R FILLER_32_24 ();
 DECAPx10_ASAP7_75t_R FILLER_32_46 ();
 DECAPx10_ASAP7_75t_R FILLER_32_68 ();
 DECAPx10_ASAP7_75t_R FILLER_32_90 ();
 FILLER_ASAP7_75t_R FILLER_32_112 ();
 FILLER_ASAP7_75t_R FILLER_32_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_184 ();
 DECAPx1_ASAP7_75t_R FILLER_32_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_200 ();
 DECAPx2_ASAP7_75t_R FILLER_32_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_213 ();
 FILLER_ASAP7_75t_R FILLER_32_226 ();
 DECAPx2_ASAP7_75t_R FILLER_32_231 ();
 FILLER_ASAP7_75t_R FILLER_32_237 ();
 DECAPx1_ASAP7_75t_R FILLER_32_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_279 ();
 DECAPx6_ASAP7_75t_R FILLER_32_295 ();
 DECAPx2_ASAP7_75t_R FILLER_32_309 ();
 FILLER_ASAP7_75t_R FILLER_32_318 ();
 DECAPx6_ASAP7_75t_R FILLER_32_333 ();
 DECAPx2_ASAP7_75t_R FILLER_32_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_379 ();
 FILLER_ASAP7_75t_R FILLER_32_398 ();
 DECAPx10_ASAP7_75t_R FILLER_32_405 ();
 DECAPx10_ASAP7_75t_R FILLER_32_433 ();
 DECAPx2_ASAP7_75t_R FILLER_32_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_461 ();
 DECAPx2_ASAP7_75t_R FILLER_32_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_470 ();
 DECAPx4_ASAP7_75t_R FILLER_32_476 ();
 DECAPx10_ASAP7_75t_R FILLER_32_500 ();
 DECAPx10_ASAP7_75t_R FILLER_32_522 ();
 DECAPx6_ASAP7_75t_R FILLER_32_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_558 ();
 DECAPx4_ASAP7_75t_R FILLER_32_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_644 ();
 DECAPx6_ASAP7_75t_R FILLER_32_651 ();
 DECAPx4_ASAP7_75t_R FILLER_32_677 ();
 FILLER_ASAP7_75t_R FILLER_32_687 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_723 ();
 DECAPx6_ASAP7_75t_R FILLER_32_732 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_746 ();
 DECAPx2_ASAP7_75t_R FILLER_32_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_32_779 ();
 DECAPx6_ASAP7_75t_R FILLER_32_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_32_802 ();
 DECAPx2_ASAP7_75t_R FILLER_32_809 ();
 DECAPx10_ASAP7_75t_R FILLER_32_830 ();
 DECAPx1_ASAP7_75t_R FILLER_32_860 ();
 DECAPx2_ASAP7_75t_R FILLER_32_882 ();
 FILLER_ASAP7_75t_R FILLER_32_888 ();
 DECAPx10_ASAP7_75t_R FILLER_32_902 ();
 DECAPx4_ASAP7_75t_R FILLER_32_924 ();
 DECAPx10_ASAP7_75t_R FILLER_33_2 ();
 DECAPx10_ASAP7_75t_R FILLER_33_24 ();
 DECAPx10_ASAP7_75t_R FILLER_33_46 ();
 DECAPx10_ASAP7_75t_R FILLER_33_68 ();
 DECAPx10_ASAP7_75t_R FILLER_33_90 ();
 DECAPx1_ASAP7_75t_R FILLER_33_112 ();
 DECAPx10_ASAP7_75t_R FILLER_33_160 ();
 DECAPx10_ASAP7_75t_R FILLER_33_182 ();
 DECAPx2_ASAP7_75t_R FILLER_33_204 ();
 FILLER_ASAP7_75t_R FILLER_33_239 ();
 FILLER_ASAP7_75t_R FILLER_33_263 ();
 DECAPx6_ASAP7_75t_R FILLER_33_268 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_282 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_291 ();
 DECAPx4_ASAP7_75t_R FILLER_33_300 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_310 ();
 DECAPx4_ASAP7_75t_R FILLER_33_334 ();
 FILLER_ASAP7_75t_R FILLER_33_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_420 ();
 DECAPx6_ASAP7_75t_R FILLER_33_438 ();
 FILLER_ASAP7_75t_R FILLER_33_452 ();
 DECAPx10_ASAP7_75t_R FILLER_33_459 ();
 DECAPx10_ASAP7_75t_R FILLER_33_481 ();
 DECAPx10_ASAP7_75t_R FILLER_33_503 ();
 DECAPx4_ASAP7_75t_R FILLER_33_525 ();
 DECAPx2_ASAP7_75t_R FILLER_33_541 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_547 ();
 DECAPx2_ASAP7_75t_R FILLER_33_558 ();
 FILLER_ASAP7_75t_R FILLER_33_570 ();
 FILLER_ASAP7_75t_R FILLER_33_578 ();
 DECAPx1_ASAP7_75t_R FILLER_33_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_614 ();
 DECAPx10_ASAP7_75t_R FILLER_33_626 ();
 DECAPx4_ASAP7_75t_R FILLER_33_648 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_658 ();
 DECAPx1_ASAP7_75t_R FILLER_33_687 ();
 DECAPx6_ASAP7_75t_R FILLER_33_703 ();
 DECAPx2_ASAP7_75t_R FILLER_33_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_723 ();
 DECAPx1_ASAP7_75t_R FILLER_33_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_740 ();
 DECAPx10_ASAP7_75t_R FILLER_33_746 ();
 DECAPx2_ASAP7_75t_R FILLER_33_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_779 ();
 DECAPx2_ASAP7_75t_R FILLER_33_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_794 ();
 DECAPx4_ASAP7_75t_R FILLER_33_802 ();
 DECAPx10_ASAP7_75t_R FILLER_33_840 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_33_862 ();
 DECAPx10_ASAP7_75t_R FILLER_33_893 ();
 DECAPx4_ASAP7_75t_R FILLER_33_915 ();
 DECAPx2_ASAP7_75t_R FILLER_33_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_33_933 ();
 DECAPx10_ASAP7_75t_R FILLER_34_2 ();
 DECAPx10_ASAP7_75t_R FILLER_34_24 ();
 DECAPx10_ASAP7_75t_R FILLER_34_46 ();
 DECAPx10_ASAP7_75t_R FILLER_34_68 ();
 DECAPx10_ASAP7_75t_R FILLER_34_90 ();
 DECAPx2_ASAP7_75t_R FILLER_34_112 ();
 DECAPx10_ASAP7_75t_R FILLER_34_147 ();
 DECAPx10_ASAP7_75t_R FILLER_34_169 ();
 DECAPx2_ASAP7_75t_R FILLER_34_191 ();
 DECAPx10_ASAP7_75t_R FILLER_34_203 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_255 ();
 DECAPx10_ASAP7_75t_R FILLER_34_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_311 ();
 DECAPx4_ASAP7_75t_R FILLER_34_327 ();
 FILLER_ASAP7_75t_R FILLER_34_337 ();
 DECAPx6_ASAP7_75t_R FILLER_34_365 ();
 DECAPx1_ASAP7_75t_R FILLER_34_379 ();
 DECAPx6_ASAP7_75t_R FILLER_34_418 ();
 DECAPx2_ASAP7_75t_R FILLER_34_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_461 ();
 DECAPx2_ASAP7_75t_R FILLER_34_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_470 ();
 DECAPx1_ASAP7_75t_R FILLER_34_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_497 ();
 FILLER_ASAP7_75t_R FILLER_34_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_537 ();
 DECAPx2_ASAP7_75t_R FILLER_34_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_596 ();
 DECAPx1_ASAP7_75t_R FILLER_34_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_610 ();
 DECAPx4_ASAP7_75t_R FILLER_34_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_624 ();
 DECAPx10_ASAP7_75t_R FILLER_34_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_670 ();
 DECAPx10_ASAP7_75t_R FILLER_34_679 ();
 DECAPx1_ASAP7_75t_R FILLER_34_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_717 ();
 DECAPx2_ASAP7_75t_R FILLER_34_724 ();
 FILLER_ASAP7_75t_R FILLER_34_730 ();
 DECAPx6_ASAP7_75t_R FILLER_34_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_765 ();
 DECAPx6_ASAP7_75t_R FILLER_34_800 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_34_814 ();
 DECAPx4_ASAP7_75t_R FILLER_34_825 ();
 DECAPx4_ASAP7_75t_R FILLER_34_853 ();
 FILLER_ASAP7_75t_R FILLER_34_863 ();
 DECAPx10_ASAP7_75t_R FILLER_34_880 ();
 DECAPx10_ASAP7_75t_R FILLER_34_902 ();
 DECAPx1_ASAP7_75t_R FILLER_34_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_34_928 ();
 DECAPx10_ASAP7_75t_R FILLER_35_2 ();
 DECAPx10_ASAP7_75t_R FILLER_35_24 ();
 DECAPx10_ASAP7_75t_R FILLER_35_46 ();
 DECAPx10_ASAP7_75t_R FILLER_35_68 ();
 DECAPx10_ASAP7_75t_R FILLER_35_90 ();
 DECAPx10_ASAP7_75t_R FILLER_35_112 ();
 DECAPx10_ASAP7_75t_R FILLER_35_134 ();
 DECAPx1_ASAP7_75t_R FILLER_35_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_160 ();
 DECAPx6_ASAP7_75t_R FILLER_35_176 ();
 DECAPx1_ASAP7_75t_R FILLER_35_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_194 ();
 DECAPx10_ASAP7_75t_R FILLER_35_211 ();
 FILLER_ASAP7_75t_R FILLER_35_233 ();
 DECAPx2_ASAP7_75t_R FILLER_35_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_255 ();
 DECAPx2_ASAP7_75t_R FILLER_35_268 ();
 DECAPx2_ASAP7_75t_R FILLER_35_280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_301 ();
 FILLER_ASAP7_75t_R FILLER_35_328 ();
 DECAPx1_ASAP7_75t_R FILLER_35_339 ();
 DECAPx4_ASAP7_75t_R FILLER_35_358 ();
 DECAPx6_ASAP7_75t_R FILLER_35_374 ();
 DECAPx2_ASAP7_75t_R FILLER_35_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_401 ();
 DECAPx1_ASAP7_75t_R FILLER_35_430 ();
 DECAPx1_ASAP7_75t_R FILLER_35_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_524 ();
 FILLER_ASAP7_75t_R FILLER_35_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_544 ();
 DECAPx1_ASAP7_75t_R FILLER_35_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_556 ();
 DECAPx10_ASAP7_75t_R FILLER_35_564 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_586 ();
 DECAPx6_ASAP7_75t_R FILLER_35_601 ();
 DECAPx2_ASAP7_75t_R FILLER_35_615 ();
 DECAPx2_ASAP7_75t_R FILLER_35_636 ();
 FILLER_ASAP7_75t_R FILLER_35_652 ();
 DECAPx10_ASAP7_75t_R FILLER_35_660 ();
 DECAPx2_ASAP7_75t_R FILLER_35_682 ();
 FILLER_ASAP7_75t_R FILLER_35_688 ();
 DECAPx2_ASAP7_75t_R FILLER_35_699 ();
 FILLER_ASAP7_75t_R FILLER_35_705 ();
 DECAPx6_ASAP7_75t_R FILLER_35_727 ();
 FILLER_ASAP7_75t_R FILLER_35_741 ();
 DECAPx6_ASAP7_75t_R FILLER_35_751 ();
 FILLER_ASAP7_75t_R FILLER_35_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_770 ();
 DECAPx6_ASAP7_75t_R FILLER_35_777 ();
 FILLER_ASAP7_75t_R FILLER_35_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_801 ();
 DECAPx4_ASAP7_75t_R FILLER_35_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_35_829 ();
 DECAPx10_ASAP7_75t_R FILLER_35_859 ();
 DECAPx2_ASAP7_75t_R FILLER_35_881 ();
 DECAPx10_ASAP7_75t_R FILLER_35_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_35_922 ();
 FILLER_ASAP7_75t_R FILLER_35_927 ();
 DECAPx10_ASAP7_75t_R FILLER_36_2 ();
 DECAPx10_ASAP7_75t_R FILLER_36_24 ();
 DECAPx10_ASAP7_75t_R FILLER_36_46 ();
 DECAPx10_ASAP7_75t_R FILLER_36_68 ();
 DECAPx6_ASAP7_75t_R FILLER_36_90 ();
 FILLER_ASAP7_75t_R FILLER_36_104 ();
 DECAPx10_ASAP7_75t_R FILLER_36_112 ();
 DECAPx4_ASAP7_75t_R FILLER_36_134 ();
 FILLER_ASAP7_75t_R FILLER_36_144 ();
 DECAPx2_ASAP7_75t_R FILLER_36_184 ();
 FILLER_ASAP7_75t_R FILLER_36_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_198 ();
 DECAPx2_ASAP7_75t_R FILLER_36_211 ();
 FILLER_ASAP7_75t_R FILLER_36_217 ();
 FILLER_ASAP7_75t_R FILLER_36_225 ();
 DECAPx6_ASAP7_75t_R FILLER_36_233 ();
 DECAPx1_ASAP7_75t_R FILLER_36_247 ();
 DECAPx2_ASAP7_75t_R FILLER_36_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_299 ();
 DECAPx1_ASAP7_75t_R FILLER_36_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_314 ();
 FILLER_ASAP7_75t_R FILLER_36_320 ();
 DECAPx4_ASAP7_75t_R FILLER_36_348 ();
 FILLER_ASAP7_75t_R FILLER_36_358 ();
 DECAPx1_ASAP7_75t_R FILLER_36_363 ();
 DECAPx2_ASAP7_75t_R FILLER_36_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_429 ();
 DECAPx1_ASAP7_75t_R FILLER_36_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_461 ();
 DECAPx1_ASAP7_75t_R FILLER_36_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_468 ();
 FILLER_ASAP7_75t_R FILLER_36_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_507 ();
 FILLER_ASAP7_75t_R FILLER_36_514 ();
 FILLER_ASAP7_75t_R FILLER_36_522 ();
 DECAPx10_ASAP7_75t_R FILLER_36_530 ();
 DECAPx6_ASAP7_75t_R FILLER_36_552 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_566 ();
 DECAPx6_ASAP7_75t_R FILLER_36_581 ();
 DECAPx1_ASAP7_75t_R FILLER_36_595 ();
 DECAPx6_ASAP7_75t_R FILLER_36_611 ();
 FILLER_ASAP7_75t_R FILLER_36_625 ();
 DECAPx1_ASAP7_75t_R FILLER_36_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_36_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_708 ();
 DECAPx6_ASAP7_75t_R FILLER_36_719 ();
 DECAPx2_ASAP7_75t_R FILLER_36_733 ();
 DECAPx10_ASAP7_75t_R FILLER_36_765 ();
 DECAPx1_ASAP7_75t_R FILLER_36_787 ();
 DECAPx10_ASAP7_75t_R FILLER_36_811 ();
 DECAPx1_ASAP7_75t_R FILLER_36_833 ();
 DECAPx4_ASAP7_75t_R FILLER_36_855 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_36_865 ();
 DECAPx2_ASAP7_75t_R FILLER_36_873 ();
 FILLER_ASAP7_75t_R FILLER_36_879 ();
 DECAPx2_ASAP7_75t_R FILLER_36_906 ();
 FILLER_ASAP7_75t_R FILLER_36_912 ();
 DECAPx10_ASAP7_75t_R FILLER_37_2 ();
 DECAPx10_ASAP7_75t_R FILLER_37_24 ();
 DECAPx10_ASAP7_75t_R FILLER_37_46 ();
 DECAPx10_ASAP7_75t_R FILLER_37_68 ();
 DECAPx4_ASAP7_75t_R FILLER_37_90 ();
 FILLER_ASAP7_75t_R FILLER_37_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_128 ();
 FILLER_ASAP7_75t_R FILLER_37_138 ();
 DECAPx2_ASAP7_75t_R FILLER_37_143 ();
 FILLER_ASAP7_75t_R FILLER_37_155 ();
 FILLER_ASAP7_75t_R FILLER_37_163 ();
 FILLER_ASAP7_75t_R FILLER_37_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_213 ();
 DECAPx6_ASAP7_75t_R FILLER_37_246 ();
 DECAPx2_ASAP7_75t_R FILLER_37_260 ();
 DECAPx1_ASAP7_75t_R FILLER_37_269 ();
 DECAPx10_ASAP7_75t_R FILLER_37_279 ();
 DECAPx10_ASAP7_75t_R FILLER_37_301 ();
 DECAPx1_ASAP7_75t_R FILLER_37_323 ();
 FILLER_ASAP7_75t_R FILLER_37_333 ();
 DECAPx6_ASAP7_75t_R FILLER_37_344 ();
 DECAPx1_ASAP7_75t_R FILLER_37_358 ();
 DECAPx1_ASAP7_75t_R FILLER_37_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_374 ();
 DECAPx4_ASAP7_75t_R FILLER_37_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_406 ();
 DECAPx6_ASAP7_75t_R FILLER_37_419 ();
 DECAPx2_ASAP7_75t_R FILLER_37_433 ();
 DECAPx6_ASAP7_75t_R FILLER_37_445 ();
 DECAPx1_ASAP7_75t_R FILLER_37_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_463 ();
 DECAPx2_ASAP7_75t_R FILLER_37_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_476 ();
 DECAPx10_ASAP7_75t_R FILLER_37_483 ();
 DECAPx10_ASAP7_75t_R FILLER_37_505 ();
 DECAPx10_ASAP7_75t_R FILLER_37_527 ();
 DECAPx4_ASAP7_75t_R FILLER_37_549 ();
 FILLER_ASAP7_75t_R FILLER_37_559 ();
 DECAPx1_ASAP7_75t_R FILLER_37_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_579 ();
 DECAPx2_ASAP7_75t_R FILLER_37_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_593 ();
 DECAPx4_ASAP7_75t_R FILLER_37_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_678 ();
 DECAPx6_ASAP7_75t_R FILLER_37_704 ();
 DECAPx2_ASAP7_75t_R FILLER_37_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_724 ();
 DECAPx1_ASAP7_75t_R FILLER_37_742 ();
 DECAPx2_ASAP7_75t_R FILLER_37_758 ();
 FILLER_ASAP7_75t_R FILLER_37_764 ();
 DECAPx2_ASAP7_75t_R FILLER_37_774 ();
 FILLER_ASAP7_75t_R FILLER_37_780 ();
 DECAPx6_ASAP7_75t_R FILLER_37_800 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_37_814 ();
 DECAPx10_ASAP7_75t_R FILLER_37_829 ();
 DECAPx1_ASAP7_75t_R FILLER_37_851 ();
 DECAPx1_ASAP7_75t_R FILLER_37_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_37_867 ();
 DECAPx10_ASAP7_75t_R FILLER_37_894 ();
 DECAPx1_ASAP7_75t_R FILLER_37_916 ();
 FILLER_ASAP7_75t_R FILLER_37_927 ();
 DECAPx10_ASAP7_75t_R FILLER_38_2 ();
 DECAPx10_ASAP7_75t_R FILLER_38_24 ();
 DECAPx10_ASAP7_75t_R FILLER_38_46 ();
 DECAPx10_ASAP7_75t_R FILLER_38_68 ();
 DECAPx2_ASAP7_75t_R FILLER_38_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_117 ();
 FILLER_ASAP7_75t_R FILLER_38_170 ();
 DECAPx6_ASAP7_75t_R FILLER_38_180 ();
 DECAPx2_ASAP7_75t_R FILLER_38_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_200 ();
 DECAPx4_ASAP7_75t_R FILLER_38_204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_214 ();
 FILLER_ASAP7_75t_R FILLER_38_232 ();
 DECAPx10_ASAP7_75t_R FILLER_38_248 ();
 DECAPx10_ASAP7_75t_R FILLER_38_270 ();
 DECAPx6_ASAP7_75t_R FILLER_38_292 ();
 FILLER_ASAP7_75t_R FILLER_38_306 ();
 DECAPx6_ASAP7_75t_R FILLER_38_314 ();
 DECAPx2_ASAP7_75t_R FILLER_38_328 ();
 DECAPx4_ASAP7_75t_R FILLER_38_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_356 ();
 DECAPx10_ASAP7_75t_R FILLER_38_360 ();
 DECAPx10_ASAP7_75t_R FILLER_38_382 ();
 DECAPx2_ASAP7_75t_R FILLER_38_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_410 ();
 DECAPx6_ASAP7_75t_R FILLER_38_425 ();
 FILLER_ASAP7_75t_R FILLER_38_445 ();
 DECAPx2_ASAP7_75t_R FILLER_38_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_459 ();
 DECAPx10_ASAP7_75t_R FILLER_38_464 ();
 DECAPx6_ASAP7_75t_R FILLER_38_496 ();
 DECAPx1_ASAP7_75t_R FILLER_38_510 ();
 DECAPx2_ASAP7_75t_R FILLER_38_520 ();
 DECAPx4_ASAP7_75t_R FILLER_38_532 ();
 FILLER_ASAP7_75t_R FILLER_38_542 ();
 DECAPx2_ASAP7_75t_R FILLER_38_556 ();
 FILLER_ASAP7_75t_R FILLER_38_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_608 ();
 DECAPx1_ASAP7_75t_R FILLER_38_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_630 ();
 DECAPx6_ASAP7_75t_R FILLER_38_639 ();
 DECAPx2_ASAP7_75t_R FILLER_38_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_672 ();
 DECAPx10_ASAP7_75t_R FILLER_38_693 ();
 DECAPx2_ASAP7_75t_R FILLER_38_715 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_721 ();
 DECAPx4_ASAP7_75t_R FILLER_38_744 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_754 ();
 FILLER_ASAP7_75t_R FILLER_38_783 ();
 DECAPx10_ASAP7_75t_R FILLER_38_788 ();
 FILLER_ASAP7_75t_R FILLER_38_810 ();
 DECAPx4_ASAP7_75t_R FILLER_38_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_850 ();
 DECAPx1_ASAP7_75t_R FILLER_38_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_38_864 ();
 DECAPx4_ASAP7_75t_R FILLER_38_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_38_895 ();
 DECAPx10_ASAP7_75t_R FILLER_38_905 ();
 FILLER_ASAP7_75t_R FILLER_38_927 ();
 DECAPx10_ASAP7_75t_R FILLER_39_2 ();
 DECAPx10_ASAP7_75t_R FILLER_39_24 ();
 DECAPx10_ASAP7_75t_R FILLER_39_46 ();
 DECAPx10_ASAP7_75t_R FILLER_39_68 ();
 DECAPx4_ASAP7_75t_R FILLER_39_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_100 ();
 FILLER_ASAP7_75t_R FILLER_39_123 ();
 DECAPx10_ASAP7_75t_R FILLER_39_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_156 ();
 DECAPx1_ASAP7_75t_R FILLER_39_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_166 ();
 DECAPx6_ASAP7_75t_R FILLER_39_170 ();
 DECAPx1_ASAP7_75t_R FILLER_39_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_188 ();
 DECAPx1_ASAP7_75t_R FILLER_39_201 ();
 DECAPx1_ASAP7_75t_R FILLER_39_208 ();
 FILLER_ASAP7_75t_R FILLER_39_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_260 ();
 DECAPx1_ASAP7_75t_R FILLER_39_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_283 ();
 DECAPx1_ASAP7_75t_R FILLER_39_306 ();
 DECAPx1_ASAP7_75t_R FILLER_39_316 ();
 DECAPx6_ASAP7_75t_R FILLER_39_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_340 ();
 DECAPx4_ASAP7_75t_R FILLER_39_369 ();
 DECAPx1_ASAP7_75t_R FILLER_39_386 ();
 DECAPx10_ASAP7_75t_R FILLER_39_396 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_418 ();
 DECAPx1_ASAP7_75t_R FILLER_39_427 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_438 ();
 DECAPx1_ASAP7_75t_R FILLER_39_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_453 ();
 DECAPx4_ASAP7_75t_R FILLER_39_468 ();
 FILLER_ASAP7_75t_R FILLER_39_478 ();
 DECAPx2_ASAP7_75t_R FILLER_39_500 ();
 DECAPx1_ASAP7_75t_R FILLER_39_513 ();
 DECAPx1_ASAP7_75t_R FILLER_39_531 ();
 DECAPx1_ASAP7_75t_R FILLER_39_548 ();
 DECAPx10_ASAP7_75t_R FILLER_39_566 ();
 DECAPx10_ASAP7_75t_R FILLER_39_588 ();
 DECAPx2_ASAP7_75t_R FILLER_39_610 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_616 ();
 DECAPx10_ASAP7_75t_R FILLER_39_625 ();
 DECAPx10_ASAP7_75t_R FILLER_39_647 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_674 ();
 DECAPx10_ASAP7_75t_R FILLER_39_680 ();
 DECAPx1_ASAP7_75t_R FILLER_39_702 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_706 ();
 DECAPx1_ASAP7_75t_R FILLER_39_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_719 ();
 DECAPx10_ASAP7_75t_R FILLER_39_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_759 ();
 DECAPx10_ASAP7_75t_R FILLER_39_778 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_39_800 ();
 DECAPx6_ASAP7_75t_R FILLER_39_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_820 ();
 DECAPx1_ASAP7_75t_R FILLER_39_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_877 ();
 FILLER_ASAP7_75t_R FILLER_39_886 ();
 DECAPx4_ASAP7_75t_R FILLER_39_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_39_924 ();
 FILLER_ASAP7_75t_R FILLER_39_927 ();
 DECAPx10_ASAP7_75t_R FILLER_40_2 ();
 DECAPx10_ASAP7_75t_R FILLER_40_24 ();
 DECAPx10_ASAP7_75t_R FILLER_40_46 ();
 DECAPx10_ASAP7_75t_R FILLER_40_68 ();
 DECAPx10_ASAP7_75t_R FILLER_40_90 ();
 DECAPx1_ASAP7_75t_R FILLER_40_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_116 ();
 DECAPx10_ASAP7_75t_R FILLER_40_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_142 ();
 DECAPx10_ASAP7_75t_R FILLER_40_149 ();
 DECAPx4_ASAP7_75t_R FILLER_40_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_181 ();
 DECAPx6_ASAP7_75t_R FILLER_40_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_224 ();
 DECAPx1_ASAP7_75t_R FILLER_40_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_234 ();
 DECAPx6_ASAP7_75t_R FILLER_40_238 ();
 DECAPx2_ASAP7_75t_R FILLER_40_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_328 ();
 DECAPx2_ASAP7_75t_R FILLER_40_339 ();
 FILLER_ASAP7_75t_R FILLER_40_345 ();
 DECAPx10_ASAP7_75t_R FILLER_40_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_395 ();
 DECAPx4_ASAP7_75t_R FILLER_40_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_455 ();
 FILLER_ASAP7_75t_R FILLER_40_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_40_500 ();
 DECAPx1_ASAP7_75t_R FILLER_40_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_522 ();
 DECAPx10_ASAP7_75t_R FILLER_40_557 ();
 DECAPx4_ASAP7_75t_R FILLER_40_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_589 ();
 DECAPx10_ASAP7_75t_R FILLER_40_596 ();
 DECAPx4_ASAP7_75t_R FILLER_40_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_628 ();
 DECAPx6_ASAP7_75t_R FILLER_40_635 ();
 DECAPx1_ASAP7_75t_R FILLER_40_649 ();
 DECAPx6_ASAP7_75t_R FILLER_40_656 ();
 DECAPx6_ASAP7_75t_R FILLER_40_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_693 ();
 DECAPx10_ASAP7_75t_R FILLER_40_723 ();
 DECAPx6_ASAP7_75t_R FILLER_40_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_759 ();
 DECAPx6_ASAP7_75t_R FILLER_40_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_40_777 ();
 DECAPx6_ASAP7_75t_R FILLER_40_784 ();
 FILLER_ASAP7_75t_R FILLER_40_798 ();
 DECAPx4_ASAP7_75t_R FILLER_40_818 ();
 FILLER_ASAP7_75t_R FILLER_40_828 ();
 FILLER_ASAP7_75t_R FILLER_40_850 ();
 DECAPx2_ASAP7_75t_R FILLER_40_858 ();
 DECAPx10_ASAP7_75t_R FILLER_40_872 ();
 FILLER_ASAP7_75t_R FILLER_40_894 ();
 DECAPx10_ASAP7_75t_R FILLER_40_908 ();
 DECAPx1_ASAP7_75t_R FILLER_40_930 ();
 DECAPx10_ASAP7_75t_R FILLER_41_2 ();
 DECAPx10_ASAP7_75t_R FILLER_41_24 ();
 DECAPx10_ASAP7_75t_R FILLER_41_46 ();
 DECAPx10_ASAP7_75t_R FILLER_41_68 ();
 DECAPx6_ASAP7_75t_R FILLER_41_90 ();
 DECAPx2_ASAP7_75t_R FILLER_41_104 ();
 DECAPx6_ASAP7_75t_R FILLER_41_119 ();
 DECAPx10_ASAP7_75t_R FILLER_41_159 ();
 DECAPx6_ASAP7_75t_R FILLER_41_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_195 ();
 DECAPx10_ASAP7_75t_R FILLER_41_201 ();
 DECAPx10_ASAP7_75t_R FILLER_41_223 ();
 DECAPx4_ASAP7_75t_R FILLER_41_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_255 ();
 DECAPx6_ASAP7_75t_R FILLER_41_268 ();
 DECAPx2_ASAP7_75t_R FILLER_41_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_295 ();
 DECAPx1_ASAP7_75t_R FILLER_41_301 ();
 FILLER_ASAP7_75t_R FILLER_41_311 ();
 DECAPx6_ASAP7_75t_R FILLER_41_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_336 ();
 FILLER_ASAP7_75t_R FILLER_41_343 ();
 FILLER_ASAP7_75t_R FILLER_41_351 ();
 DECAPx2_ASAP7_75t_R FILLER_41_373 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_387 ();
 DECAPx10_ASAP7_75t_R FILLER_41_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_445 ();
 DECAPx2_ASAP7_75t_R FILLER_41_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_476 ();
 DECAPx4_ASAP7_75t_R FILLER_41_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_496 ();
 DECAPx10_ASAP7_75t_R FILLER_41_516 ();
 DECAPx10_ASAP7_75t_R FILLER_41_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_560 ();
 FILLER_ASAP7_75t_R FILLER_41_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_579 ();
 DECAPx2_ASAP7_75t_R FILLER_41_586 ();
 FILLER_ASAP7_75t_R FILLER_41_592 ();
 DECAPx4_ASAP7_75t_R FILLER_41_607 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_617 ();
 DECAPx4_ASAP7_75t_R FILLER_41_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_668 ();
 DECAPx1_ASAP7_75t_R FILLER_41_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_693 ();
 FILLER_ASAP7_75t_R FILLER_41_703 ();
 DECAPx6_ASAP7_75t_R FILLER_41_720 ();
 DECAPx2_ASAP7_75t_R FILLER_41_734 ();
 DECAPx6_ASAP7_75t_R FILLER_41_761 ();
 DECAPx2_ASAP7_75t_R FILLER_41_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_781 ();
 DECAPx4_ASAP7_75t_R FILLER_41_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_795 ();
 FILLER_ASAP7_75t_R FILLER_41_805 ();
 DECAPx4_ASAP7_75t_R FILLER_41_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_41_837 ();
 DECAPx2_ASAP7_75t_R FILLER_41_848 ();
 DECAPx10_ASAP7_75t_R FILLER_41_862 ();
 DECAPx10_ASAP7_75t_R FILLER_41_884 ();
 DECAPx6_ASAP7_75t_R FILLER_41_906 ();
 DECAPx1_ASAP7_75t_R FILLER_41_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_41_924 ();
 FILLER_ASAP7_75t_R FILLER_41_927 ();
 DECAPx10_ASAP7_75t_R FILLER_42_2 ();
 DECAPx10_ASAP7_75t_R FILLER_42_24 ();
 DECAPx10_ASAP7_75t_R FILLER_42_46 ();
 DECAPx10_ASAP7_75t_R FILLER_42_68 ();
 DECAPx4_ASAP7_75t_R FILLER_42_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_100 ();
 DECAPx4_ASAP7_75t_R FILLER_42_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_137 ();
 DECAPx1_ASAP7_75t_R FILLER_42_144 ();
 DECAPx6_ASAP7_75t_R FILLER_42_151 ();
 DECAPx1_ASAP7_75t_R FILLER_42_165 ();
 DECAPx2_ASAP7_75t_R FILLER_42_172 ();
 DECAPx2_ASAP7_75t_R FILLER_42_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_190 ();
 DECAPx6_ASAP7_75t_R FILLER_42_199 ();
 DECAPx1_ASAP7_75t_R FILLER_42_213 ();
 DECAPx1_ASAP7_75t_R FILLER_42_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_227 ();
 DECAPx6_ASAP7_75t_R FILLER_42_234 ();
 FILLER_ASAP7_75t_R FILLER_42_248 ();
 DECAPx10_ASAP7_75t_R FILLER_42_276 ();
 DECAPx10_ASAP7_75t_R FILLER_42_298 ();
 DECAPx2_ASAP7_75t_R FILLER_42_320 ();
 FILLER_ASAP7_75t_R FILLER_42_326 ();
 FILLER_ASAP7_75t_R FILLER_42_357 ();
 DECAPx6_ASAP7_75t_R FILLER_42_374 ();
 DECAPx2_ASAP7_75t_R FILLER_42_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_401 ();
 FILLER_ASAP7_75t_R FILLER_42_411 ();
 DECAPx1_ASAP7_75t_R FILLER_42_421 ();
 DECAPx6_ASAP7_75t_R FILLER_42_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_450 ();
 DECAPx1_ASAP7_75t_R FILLER_42_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_464 ();
 DECAPx6_ASAP7_75t_R FILLER_42_471 ();
 DECAPx2_ASAP7_75t_R FILLER_42_485 ();
 DECAPx6_ASAP7_75t_R FILLER_42_497 ();
 DECAPx2_ASAP7_75t_R FILLER_42_511 ();
 DECAPx4_ASAP7_75t_R FILLER_42_529 ();
 FILLER_ASAP7_75t_R FILLER_42_539 ();
 DECAPx2_ASAP7_75t_R FILLER_42_548 ();
 FILLER_ASAP7_75t_R FILLER_42_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_594 ();
 DECAPx1_ASAP7_75t_R FILLER_42_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_604 ();
 DECAPx2_ASAP7_75t_R FILLER_42_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_617 ();
 DECAPx2_ASAP7_75t_R FILLER_42_622 ();
 FILLER_ASAP7_75t_R FILLER_42_628 ();
 DECAPx1_ASAP7_75t_R FILLER_42_651 ();
 DECAPx4_ASAP7_75t_R FILLER_42_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_682 ();
 DECAPx4_ASAP7_75t_R FILLER_42_698 ();
 FILLER_ASAP7_75t_R FILLER_42_708 ();
 DECAPx6_ASAP7_75t_R FILLER_42_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_732 ();
 FILLER_ASAP7_75t_R FILLER_42_741 ();
 DECAPx6_ASAP7_75t_R FILLER_42_746 ();
 DECAPx2_ASAP7_75t_R FILLER_42_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_42_766 ();
 DECAPx1_ASAP7_75t_R FILLER_42_775 ();
 DECAPx1_ASAP7_75t_R FILLER_42_794 ();
 DECAPx2_ASAP7_75t_R FILLER_42_804 ();
 DECAPx6_ASAP7_75t_R FILLER_42_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_42_832 ();
 DECAPx10_ASAP7_75t_R FILLER_42_841 ();
 DECAPx6_ASAP7_75t_R FILLER_42_863 ();
 DECAPx10_ASAP7_75t_R FILLER_42_890 ();
 DECAPx10_ASAP7_75t_R FILLER_42_912 ();
 DECAPx10_ASAP7_75t_R FILLER_43_2 ();
 DECAPx10_ASAP7_75t_R FILLER_43_24 ();
 DECAPx10_ASAP7_75t_R FILLER_43_46 ();
 DECAPx10_ASAP7_75t_R FILLER_43_68 ();
 DECAPx6_ASAP7_75t_R FILLER_43_90 ();
 FILLER_ASAP7_75t_R FILLER_43_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_133 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_157 ();
 FILLER_ASAP7_75t_R FILLER_43_164 ();
 DECAPx1_ASAP7_75t_R FILLER_43_180 ();
 FILLER_ASAP7_75t_R FILLER_43_210 ();
 DECAPx10_ASAP7_75t_R FILLER_43_241 ();
 FILLER_ASAP7_75t_R FILLER_43_263 ();
 DECAPx1_ASAP7_75t_R FILLER_43_268 ();
 DECAPx6_ASAP7_75t_R FILLER_43_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_289 ();
 DECAPx1_ASAP7_75t_R FILLER_43_296 ();
 DECAPx6_ASAP7_75t_R FILLER_43_308 ();
 DECAPx1_ASAP7_75t_R FILLER_43_322 ();
 DECAPx1_ASAP7_75t_R FILLER_43_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_342 ();
 DECAPx10_ASAP7_75t_R FILLER_43_346 ();
 DECAPx2_ASAP7_75t_R FILLER_43_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_374 ();
 DECAPx2_ASAP7_75t_R FILLER_43_383 ();
 DECAPx6_ASAP7_75t_R FILLER_43_392 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_406 ();
 FILLER_ASAP7_75t_R FILLER_43_424 ();
 DECAPx6_ASAP7_75t_R FILLER_43_432 ();
 DECAPx2_ASAP7_75t_R FILLER_43_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_452 ();
 DECAPx1_ASAP7_75t_R FILLER_43_458 ();
 FILLER_ASAP7_75t_R FILLER_43_479 ();
 DECAPx10_ASAP7_75t_R FILLER_43_487 ();
 DECAPx4_ASAP7_75t_R FILLER_43_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_519 ();
 DECAPx2_ASAP7_75t_R FILLER_43_532 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_604 ();
 DECAPx2_ASAP7_75t_R FILLER_43_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_635 ();
 DECAPx1_ASAP7_75t_R FILLER_43_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_648 ();
 DECAPx4_ASAP7_75t_R FILLER_43_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_687 ();
 DECAPx6_ASAP7_75t_R FILLER_43_702 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_716 ();
 DECAPx4_ASAP7_75t_R FILLER_43_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_792 ();
 DECAPx6_ASAP7_75t_R FILLER_43_807 ();
 DECAPx1_ASAP7_75t_R FILLER_43_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_825 ();
 DECAPx10_ASAP7_75t_R FILLER_43_832 ();
 DECAPx6_ASAP7_75t_R FILLER_43_854 ();
 DECAPx2_ASAP7_75t_R FILLER_43_868 ();
 DECAPx10_ASAP7_75t_R FILLER_43_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_43_922 ();
 DECAPx2_ASAP7_75t_R FILLER_43_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_43_933 ();
 DECAPx10_ASAP7_75t_R FILLER_44_2 ();
 DECAPx10_ASAP7_75t_R FILLER_44_24 ();
 DECAPx10_ASAP7_75t_R FILLER_44_46 ();
 DECAPx10_ASAP7_75t_R FILLER_44_68 ();
 DECAPx2_ASAP7_75t_R FILLER_44_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_96 ();
 DECAPx6_ASAP7_75t_R FILLER_44_100 ();
 FILLER_ASAP7_75t_R FILLER_44_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_153 ();
 DECAPx1_ASAP7_75t_R FILLER_44_194 ();
 FILLER_ASAP7_75t_R FILLER_44_201 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_241 ();
 DECAPx10_ASAP7_75t_R FILLER_44_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_284 ();
 DECAPx2_ASAP7_75t_R FILLER_44_314 ();
 DECAPx10_ASAP7_75t_R FILLER_44_346 ();
 DECAPx2_ASAP7_75t_R FILLER_44_368 ();
 DECAPx4_ASAP7_75t_R FILLER_44_403 ();
 DECAPx2_ASAP7_75t_R FILLER_44_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_439 ();
 DECAPx1_ASAP7_75t_R FILLER_44_446 ();
 DECAPx6_ASAP7_75t_R FILLER_44_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_478 ();
 DECAPx10_ASAP7_75t_R FILLER_44_498 ();
 DECAPx4_ASAP7_75t_R FILLER_44_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_530 ();
 DECAPx10_ASAP7_75t_R FILLER_44_551 ();
 DECAPx6_ASAP7_75t_R FILLER_44_573 ();
 FILLER_ASAP7_75t_R FILLER_44_587 ();
 DECAPx1_ASAP7_75t_R FILLER_44_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_599 ();
 DECAPx2_ASAP7_75t_R FILLER_44_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_632 ();
 DECAPx2_ASAP7_75t_R FILLER_44_638 ();
 DECAPx6_ASAP7_75t_R FILLER_44_651 ();
 FILLER_ASAP7_75t_R FILLER_44_665 ();
 DECAPx2_ASAP7_75t_R FILLER_44_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_693 ();
 DECAPx2_ASAP7_75t_R FILLER_44_714 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_768 ();
 DECAPx4_ASAP7_75t_R FILLER_44_784 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_794 ();
 DECAPx1_ASAP7_75t_R FILLER_44_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_44_842 ();
 FILLER_ASAP7_75t_R FILLER_44_851 ();
 DECAPx6_ASAP7_75t_R FILLER_44_864 ();
 DECAPx1_ASAP7_75t_R FILLER_44_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_44_882 ();
 DECAPx2_ASAP7_75t_R FILLER_44_889 ();
 FILLER_ASAP7_75t_R FILLER_44_895 ();
 DECAPx10_ASAP7_75t_R FILLER_44_903 ();
 DECAPx1_ASAP7_75t_R FILLER_44_925 ();
 DECAPx10_ASAP7_75t_R FILLER_45_2 ();
 DECAPx10_ASAP7_75t_R FILLER_45_24 ();
 DECAPx10_ASAP7_75t_R FILLER_45_46 ();
 DECAPx6_ASAP7_75t_R FILLER_45_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_82 ();
 DECAPx6_ASAP7_75t_R FILLER_45_115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_129 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_141 ();
 DECAPx1_ASAP7_75t_R FILLER_45_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_175 ();
 DECAPx2_ASAP7_75t_R FILLER_45_198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_204 ();
 DECAPx4_ASAP7_75t_R FILLER_45_222 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_265 ();
 DECAPx1_ASAP7_75t_R FILLER_45_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_286 ();
 DECAPx1_ASAP7_75t_R FILLER_45_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_297 ();
 FILLER_ASAP7_75t_R FILLER_45_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_332 ();
 DECAPx6_ASAP7_75t_R FILLER_45_338 ();
 DECAPx1_ASAP7_75t_R FILLER_45_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_356 ();
 FILLER_ASAP7_75t_R FILLER_45_373 ();
 DECAPx10_ASAP7_75t_R FILLER_45_381 ();
 DECAPx10_ASAP7_75t_R FILLER_45_403 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_448 ();
 DECAPx2_ASAP7_75t_R FILLER_45_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_463 ();
 DECAPx1_ASAP7_75t_R FILLER_45_486 ();
 DECAPx1_ASAP7_75t_R FILLER_45_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_506 ();
 DECAPx2_ASAP7_75t_R FILLER_45_520 ();
 DECAPx6_ASAP7_75t_R FILLER_45_534 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_548 ();
 DECAPx10_ASAP7_75t_R FILLER_45_557 ();
 DECAPx10_ASAP7_75t_R FILLER_45_579 ();
 DECAPx1_ASAP7_75t_R FILLER_45_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_605 ();
 DECAPx6_ASAP7_75t_R FILLER_45_612 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_626 ();
 DECAPx4_ASAP7_75t_R FILLER_45_643 ();
 FILLER_ASAP7_75t_R FILLER_45_653 ();
 DECAPx1_ASAP7_75t_R FILLER_45_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_666 ();
 DECAPx10_ASAP7_75t_R FILLER_45_674 ();
 DECAPx6_ASAP7_75t_R FILLER_45_696 ();
 DECAPx2_ASAP7_75t_R FILLER_45_710 ();
 DECAPx10_ASAP7_75t_R FILLER_45_742 ();
 DECAPx10_ASAP7_75t_R FILLER_45_764 ();
 DECAPx1_ASAP7_75t_R FILLER_45_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_45_845 ();
 DECAPx6_ASAP7_75t_R FILLER_45_875 ();
 FILLER_ASAP7_75t_R FILLER_45_889 ();
 DECAPx6_ASAP7_75t_R FILLER_45_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_924 ();
 DECAPx2_ASAP7_75t_R FILLER_45_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_45_933 ();
 DECAPx10_ASAP7_75t_R FILLER_46_2 ();
 DECAPx10_ASAP7_75t_R FILLER_46_24 ();
 DECAPx10_ASAP7_75t_R FILLER_46_46 ();
 DECAPx6_ASAP7_75t_R FILLER_46_68 ();
 DECAPx2_ASAP7_75t_R FILLER_46_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_88 ();
 DECAPx10_ASAP7_75t_R FILLER_46_121 ();
 DECAPx10_ASAP7_75t_R FILLER_46_143 ();
 DECAPx10_ASAP7_75t_R FILLER_46_165 ();
 DECAPx10_ASAP7_75t_R FILLER_46_187 ();
 DECAPx10_ASAP7_75t_R FILLER_46_209 ();
 DECAPx2_ASAP7_75t_R FILLER_46_231 ();
 FILLER_ASAP7_75t_R FILLER_46_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_290 ();
 DECAPx4_ASAP7_75t_R FILLER_46_297 ();
 DECAPx10_ASAP7_75t_R FILLER_46_313 ();
 DECAPx2_ASAP7_75t_R FILLER_46_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_341 ();
 DECAPx2_ASAP7_75t_R FILLER_46_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_377 ();
 DECAPx6_ASAP7_75t_R FILLER_46_386 ();
 DECAPx1_ASAP7_75t_R FILLER_46_400 ();
 DECAPx4_ASAP7_75t_R FILLER_46_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_461 ();
 FILLER_ASAP7_75t_R FILLER_46_464 ();
 DECAPx10_ASAP7_75t_R FILLER_46_469 ();
 DECAPx2_ASAP7_75t_R FILLER_46_542 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_548 ();
 DECAPx6_ASAP7_75t_R FILLER_46_578 ();
 DECAPx1_ASAP7_75t_R FILLER_46_592 ();
 FILLER_ASAP7_75t_R FILLER_46_603 ();
 DECAPx1_ASAP7_75t_R FILLER_46_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_615 ();
 FILLER_ASAP7_75t_R FILLER_46_623 ();
 DECAPx10_ASAP7_75t_R FILLER_46_645 ();
 DECAPx2_ASAP7_75t_R FILLER_46_667 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_673 ();
 DECAPx1_ASAP7_75t_R FILLER_46_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_687 ();
 DECAPx10_ASAP7_75t_R FILLER_46_691 ();
 DECAPx10_ASAP7_75t_R FILLER_46_713 ();
 DECAPx10_ASAP7_75t_R FILLER_46_735 ();
 DECAPx10_ASAP7_75t_R FILLER_46_757 ();
 DECAPx10_ASAP7_75t_R FILLER_46_779 ();
 DECAPx2_ASAP7_75t_R FILLER_46_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_807 ();
 DECAPx2_ASAP7_75t_R FILLER_46_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_818 ();
 FILLER_ASAP7_75t_R FILLER_46_831 ();
 DECAPx1_ASAP7_75t_R FILLER_46_846 ();
 DECAPx2_ASAP7_75t_R FILLER_46_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_868 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_46_877 ();
 DECAPx4_ASAP7_75t_R FILLER_46_883 ();
 DECAPx6_ASAP7_75t_R FILLER_46_913 ();
 DECAPx2_ASAP7_75t_R FILLER_46_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_46_933 ();
 DECAPx10_ASAP7_75t_R FILLER_47_2 ();
 DECAPx10_ASAP7_75t_R FILLER_47_24 ();
 DECAPx10_ASAP7_75t_R FILLER_47_46 ();
 DECAPx10_ASAP7_75t_R FILLER_47_68 ();
 DECAPx4_ASAP7_75t_R FILLER_47_122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_132 ();
 DECAPx10_ASAP7_75t_R FILLER_47_141 ();
 DECAPx1_ASAP7_75t_R FILLER_47_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_173 ();
 DECAPx2_ASAP7_75t_R FILLER_47_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_183 ();
 FILLER_ASAP7_75t_R FILLER_47_210 ();
 DECAPx1_ASAP7_75t_R FILLER_47_218 ();
 DECAPx10_ASAP7_75t_R FILLER_47_234 ();
 DECAPx2_ASAP7_75t_R FILLER_47_256 ();
 FILLER_ASAP7_75t_R FILLER_47_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_273 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_280 ();
 FILLER_ASAP7_75t_R FILLER_47_331 ();
 DECAPx2_ASAP7_75t_R FILLER_47_339 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_345 ();
 DECAPx4_ASAP7_75t_R FILLER_47_363 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_373 ();
 FILLER_ASAP7_75t_R FILLER_47_402 ();
 FILLER_ASAP7_75t_R FILLER_47_430 ();
 DECAPx4_ASAP7_75t_R FILLER_47_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_497 ();
 DECAPx2_ASAP7_75t_R FILLER_47_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_516 ();
 DECAPx2_ASAP7_75t_R FILLER_47_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_543 ();
 DECAPx6_ASAP7_75t_R FILLER_47_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_564 ();
 DECAPx2_ASAP7_75t_R FILLER_47_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_593 ();
 DECAPx4_ASAP7_75t_R FILLER_47_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_701 ();
 DECAPx10_ASAP7_75t_R FILLER_47_708 ();
 DECAPx2_ASAP7_75t_R FILLER_47_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_47_736 ();
 DECAPx4_ASAP7_75t_R FILLER_47_744 ();
 DECAPx6_ASAP7_75t_R FILLER_47_768 ();
 DECAPx10_ASAP7_75t_R FILLER_47_796 ();
 DECAPx10_ASAP7_75t_R FILLER_47_818 ();
 DECAPx6_ASAP7_75t_R FILLER_47_840 ();
 DECAPx1_ASAP7_75t_R FILLER_47_854 ();
 DECAPx10_ASAP7_75t_R FILLER_47_890 ();
 DECAPx4_ASAP7_75t_R FILLER_47_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_47_922 ();
 FILLER_ASAP7_75t_R FILLER_47_927 ();
 DECAPx10_ASAP7_75t_R FILLER_48_2 ();
 DECAPx10_ASAP7_75t_R FILLER_48_24 ();
 DECAPx10_ASAP7_75t_R FILLER_48_46 ();
 DECAPx10_ASAP7_75t_R FILLER_48_68 ();
 DECAPx4_ASAP7_75t_R FILLER_48_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_106 ();
 DECAPx1_ASAP7_75t_R FILLER_48_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_122 ();
 FILLER_ASAP7_75t_R FILLER_48_151 ();
 DECAPx10_ASAP7_75t_R FILLER_48_239 ();
 DECAPx10_ASAP7_75t_R FILLER_48_261 ();
 DECAPx1_ASAP7_75t_R FILLER_48_283 ();
 DECAPx1_ASAP7_75t_R FILLER_48_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_297 ();
 DECAPx6_ASAP7_75t_R FILLER_48_301 ();
 DECAPx1_ASAP7_75t_R FILLER_48_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_319 ();
 DECAPx6_ASAP7_75t_R FILLER_48_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_412 ();
 DECAPx1_ASAP7_75t_R FILLER_48_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_427 ();
 DECAPx10_ASAP7_75t_R FILLER_48_431 ();
 DECAPx2_ASAP7_75t_R FILLER_48_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_459 ();
 DECAPx6_ASAP7_75t_R FILLER_48_486 ();
 DECAPx2_ASAP7_75t_R FILLER_48_500 ();
 DECAPx1_ASAP7_75t_R FILLER_48_513 ();
 DECAPx4_ASAP7_75t_R FILLER_48_523 ();
 FILLER_ASAP7_75t_R FILLER_48_533 ();
 DECAPx1_ASAP7_75t_R FILLER_48_542 ();
 DECAPx2_ASAP7_75t_R FILLER_48_573 ();
 DECAPx2_ASAP7_75t_R FILLER_48_613 ();
 FILLER_ASAP7_75t_R FILLER_48_619 ();
 DECAPx4_ASAP7_75t_R FILLER_48_632 ();
 DECAPx10_ASAP7_75t_R FILLER_48_679 ();
 DECAPx2_ASAP7_75t_R FILLER_48_728 ();
 FILLER_ASAP7_75t_R FILLER_48_734 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_48_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_779 ();
 DECAPx2_ASAP7_75t_R FILLER_48_800 ();
 FILLER_ASAP7_75t_R FILLER_48_806 ();
 DECAPx1_ASAP7_75t_R FILLER_48_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_48_820 ();
 DECAPx10_ASAP7_75t_R FILLER_48_827 ();
 DECAPx6_ASAP7_75t_R FILLER_48_849 ();
 DECAPx2_ASAP7_75t_R FILLER_48_863 ();
 DECAPx10_ASAP7_75t_R FILLER_48_876 ();
 DECAPx10_ASAP7_75t_R FILLER_48_898 ();
 DECAPx6_ASAP7_75t_R FILLER_48_920 ();
 DECAPx10_ASAP7_75t_R FILLER_49_2 ();
 DECAPx10_ASAP7_75t_R FILLER_49_24 ();
 DECAPx10_ASAP7_75t_R FILLER_49_46 ();
 DECAPx10_ASAP7_75t_R FILLER_49_68 ();
 DECAPx10_ASAP7_75t_R FILLER_49_90 ();
 DECAPx4_ASAP7_75t_R FILLER_49_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_128 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_137 ();
 DECAPx6_ASAP7_75t_R FILLER_49_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_157 ();
 DECAPx1_ASAP7_75t_R FILLER_49_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_168 ();
 DECAPx4_ASAP7_75t_R FILLER_49_172 ();
 FILLER_ASAP7_75t_R FILLER_49_188 ();
 FILLER_ASAP7_75t_R FILLER_49_198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_206 ();
 DECAPx1_ASAP7_75t_R FILLER_49_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_219 ();
 FILLER_ASAP7_75t_R FILLER_49_223 ();
 DECAPx1_ASAP7_75t_R FILLER_49_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_246 ();
 DECAPx2_ASAP7_75t_R FILLER_49_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_256 ();
 DECAPx10_ASAP7_75t_R FILLER_49_265 ();
 DECAPx10_ASAP7_75t_R FILLER_49_287 ();
 DECAPx2_ASAP7_75t_R FILLER_49_309 ();
 DECAPx10_ASAP7_75t_R FILLER_49_322 ();
 FILLER_ASAP7_75t_R FILLER_49_344 ();
 DECAPx1_ASAP7_75t_R FILLER_49_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_356 ();
 DECAPx1_ASAP7_75t_R FILLER_49_387 ();
 DECAPx10_ASAP7_75t_R FILLER_49_438 ();
 DECAPx6_ASAP7_75t_R FILLER_49_460 ();
 DECAPx1_ASAP7_75t_R FILLER_49_474 ();
 DECAPx10_ASAP7_75t_R FILLER_49_484 ();
 DECAPx10_ASAP7_75t_R FILLER_49_506 ();
 DECAPx6_ASAP7_75t_R FILLER_49_528 ();
 DECAPx1_ASAP7_75t_R FILLER_49_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_546 ();
 DECAPx4_ASAP7_75t_R FILLER_49_553 ();
 DECAPx4_ASAP7_75t_R FILLER_49_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_579 ();
 DECAPx10_ASAP7_75t_R FILLER_49_600 ();
 DECAPx10_ASAP7_75t_R FILLER_49_622 ();
 FILLER_ASAP7_75t_R FILLER_49_644 ();
 DECAPx1_ASAP7_75t_R FILLER_49_652 ();
 DECAPx2_ASAP7_75t_R FILLER_49_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_682 ();
 DECAPx2_ASAP7_75t_R FILLER_49_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_709 ();
 DECAPx6_ASAP7_75t_R FILLER_49_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_732 ();
 DECAPx4_ASAP7_75t_R FILLER_49_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_751 ();
 DECAPx6_ASAP7_75t_R FILLER_49_758 ();
 DECAPx1_ASAP7_75t_R FILLER_49_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_776 ();
 FILLER_ASAP7_75t_R FILLER_49_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_834 ();
 DECAPx10_ASAP7_75t_R FILLER_49_847 ();
 DECAPx2_ASAP7_75t_R FILLER_49_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_875 ();
 DECAPx10_ASAP7_75t_R FILLER_49_886 ();
 DECAPx6_ASAP7_75t_R FILLER_49_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_49_922 ();
 DECAPx2_ASAP7_75t_R FILLER_49_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_49_933 ();
 DECAPx10_ASAP7_75t_R FILLER_50_2 ();
 DECAPx10_ASAP7_75t_R FILLER_50_24 ();
 DECAPx10_ASAP7_75t_R FILLER_50_46 ();
 DECAPx10_ASAP7_75t_R FILLER_50_68 ();
 DECAPx10_ASAP7_75t_R FILLER_50_90 ();
 DECAPx10_ASAP7_75t_R FILLER_50_112 ();
 DECAPx1_ASAP7_75t_R FILLER_50_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_138 ();
 DECAPx4_ASAP7_75t_R FILLER_50_145 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_155 ();
 DECAPx10_ASAP7_75t_R FILLER_50_184 ();
 DECAPx10_ASAP7_75t_R FILLER_50_206 ();
 DECAPx1_ASAP7_75t_R FILLER_50_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_314 ();
 DECAPx2_ASAP7_75t_R FILLER_50_321 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_327 ();
 DECAPx4_ASAP7_75t_R FILLER_50_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_358 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_393 ();
 DECAPx2_ASAP7_75t_R FILLER_50_404 ();
 FILLER_ASAP7_75t_R FILLER_50_410 ();
 DECAPx2_ASAP7_75t_R FILLER_50_421 ();
 DECAPx10_ASAP7_75t_R FILLER_50_430 ();
 DECAPx4_ASAP7_75t_R FILLER_50_452 ();
 DECAPx1_ASAP7_75t_R FILLER_50_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_488 ();
 DECAPx2_ASAP7_75t_R FILLER_50_495 ();
 DECAPx10_ASAP7_75t_R FILLER_50_507 ();
 DECAPx10_ASAP7_75t_R FILLER_50_536 ();
 DECAPx4_ASAP7_75t_R FILLER_50_558 ();
 FILLER_ASAP7_75t_R FILLER_50_568 ();
 DECAPx4_ASAP7_75t_R FILLER_50_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_586 ();
 DECAPx10_ASAP7_75t_R FILLER_50_593 ();
 DECAPx6_ASAP7_75t_R FILLER_50_615 ();
 DECAPx2_ASAP7_75t_R FILLER_50_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_635 ();
 DECAPx10_ASAP7_75t_R FILLER_50_642 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_683 ();
 DECAPx10_ASAP7_75t_R FILLER_50_691 ();
 DECAPx4_ASAP7_75t_R FILLER_50_713 ();
 FILLER_ASAP7_75t_R FILLER_50_723 ();
 FILLER_ASAP7_75t_R FILLER_50_739 ();
 FILLER_ASAP7_75t_R FILLER_50_745 ();
 DECAPx2_ASAP7_75t_R FILLER_50_753 ();
 DECAPx10_ASAP7_75t_R FILLER_50_771 ();
 DECAPx6_ASAP7_75t_R FILLER_50_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_807 ();
 DECAPx4_ASAP7_75t_R FILLER_50_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_50_826 ();
 DECAPx1_ASAP7_75t_R FILLER_50_873 ();
 DECAPx10_ASAP7_75t_R FILLER_50_897 ();
 DECAPx6_ASAP7_75t_R FILLER_50_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_50_933 ();
 DECAPx10_ASAP7_75t_R FILLER_51_2 ();
 DECAPx10_ASAP7_75t_R FILLER_51_24 ();
 DECAPx10_ASAP7_75t_R FILLER_51_46 ();
 DECAPx6_ASAP7_75t_R FILLER_51_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_82 ();
 DECAPx2_ASAP7_75t_R FILLER_51_103 ();
 FILLER_ASAP7_75t_R FILLER_51_109 ();
 DECAPx1_ASAP7_75t_R FILLER_51_117 ();
 DECAPx2_ASAP7_75t_R FILLER_51_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_133 ();
 DECAPx2_ASAP7_75t_R FILLER_51_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_168 ();
 DECAPx10_ASAP7_75t_R FILLER_51_178 ();
 DECAPx10_ASAP7_75t_R FILLER_51_200 ();
 DECAPx6_ASAP7_75t_R FILLER_51_222 ();
 DECAPx6_ASAP7_75t_R FILLER_51_242 ();
 DECAPx2_ASAP7_75t_R FILLER_51_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_262 ();
 DECAPx2_ASAP7_75t_R FILLER_51_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_325 ();
 FILLER_ASAP7_75t_R FILLER_51_340 ();
 FILLER_ASAP7_75t_R FILLER_51_403 ();
 DECAPx6_ASAP7_75t_R FILLER_51_411 ();
 DECAPx1_ASAP7_75t_R FILLER_51_425 ();
 DECAPx2_ASAP7_75t_R FILLER_51_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_449 ();
 DECAPx2_ASAP7_75t_R FILLER_51_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_485 ();
 DECAPx1_ASAP7_75t_R FILLER_51_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_51_521 ();
 DECAPx6_ASAP7_75t_R FILLER_51_547 ();
 DECAPx1_ASAP7_75t_R FILLER_51_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_565 ();
 DECAPx4_ASAP7_75t_R FILLER_51_603 ();
 DECAPx1_ASAP7_75t_R FILLER_51_619 ();
 DECAPx10_ASAP7_75t_R FILLER_51_649 ();
 DECAPx10_ASAP7_75t_R FILLER_51_671 ();
 DECAPx2_ASAP7_75t_R FILLER_51_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_705 ();
 DECAPx4_ASAP7_75t_R FILLER_51_712 ();
 DECAPx6_ASAP7_75t_R FILLER_51_749 ();
 FILLER_ASAP7_75t_R FILLER_51_763 ();
 DECAPx6_ASAP7_75t_R FILLER_51_772 ();
 DECAPx1_ASAP7_75t_R FILLER_51_786 ();
 DECAPx10_ASAP7_75t_R FILLER_51_796 ();
 DECAPx6_ASAP7_75t_R FILLER_51_818 ();
 DECAPx2_ASAP7_75t_R FILLER_51_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_838 ();
 DECAPx1_ASAP7_75t_R FILLER_51_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_854 ();
 DECAPx4_ASAP7_75t_R FILLER_51_865 ();
 DECAPx10_ASAP7_75t_R FILLER_51_881 ();
 DECAPx10_ASAP7_75t_R FILLER_51_903 ();
 DECAPx2_ASAP7_75t_R FILLER_51_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_51_933 ();
 DECAPx10_ASAP7_75t_R FILLER_52_2 ();
 DECAPx10_ASAP7_75t_R FILLER_52_24 ();
 DECAPx10_ASAP7_75t_R FILLER_52_46 ();
 DECAPx4_ASAP7_75t_R FILLER_52_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_78 ();
 DECAPx1_ASAP7_75t_R FILLER_52_111 ();
 DECAPx1_ASAP7_75t_R FILLER_52_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_127 ();
 DECAPx4_ASAP7_75t_R FILLER_52_168 ();
 FILLER_ASAP7_75t_R FILLER_52_178 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_183 ();
 DECAPx1_ASAP7_75t_R FILLER_52_198 ();
 DECAPx10_ASAP7_75t_R FILLER_52_217 ();
 DECAPx2_ASAP7_75t_R FILLER_52_239 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_245 ();
 DECAPx4_ASAP7_75t_R FILLER_52_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_351 ();
 DECAPx4_ASAP7_75t_R FILLER_52_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_396 ();
 DECAPx4_ASAP7_75t_R FILLER_52_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_421 ();
 DECAPx4_ASAP7_75t_R FILLER_52_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_464 ();
 DECAPx1_ASAP7_75t_R FILLER_52_481 ();
 FILLER_ASAP7_75t_R FILLER_52_495 ();
 DECAPx4_ASAP7_75t_R FILLER_52_509 ();
 FILLER_ASAP7_75t_R FILLER_52_519 ();
 DECAPx1_ASAP7_75t_R FILLER_52_531 ();
 DECAPx2_ASAP7_75t_R FILLER_52_553 ();
 FILLER_ASAP7_75t_R FILLER_52_559 ();
 DECAPx2_ASAP7_75t_R FILLER_52_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_582 ();
 DECAPx2_ASAP7_75t_R FILLER_52_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_630 ();
 FILLER_ASAP7_75t_R FILLER_52_660 ();
 DECAPx1_ASAP7_75t_R FILLER_52_668 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_672 ();
 DECAPx2_ASAP7_75t_R FILLER_52_685 ();
 FILLER_ASAP7_75t_R FILLER_52_698 ();
 DECAPx1_ASAP7_75t_R FILLER_52_720 ();
 DECAPx2_ASAP7_75t_R FILLER_52_730 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_736 ();
 DECAPx2_ASAP7_75t_R FILLER_52_763 ();
 FILLER_ASAP7_75t_R FILLER_52_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_775 ();
 DECAPx1_ASAP7_75t_R FILLER_52_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_787 ();
 DECAPx1_ASAP7_75t_R FILLER_52_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_52_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_812 ();
 DECAPx10_ASAP7_75t_R FILLER_52_829 ();
 DECAPx10_ASAP7_75t_R FILLER_52_851 ();
 DECAPx10_ASAP7_75t_R FILLER_52_873 ();
 DECAPx10_ASAP7_75t_R FILLER_52_895 ();
 DECAPx6_ASAP7_75t_R FILLER_52_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_52_931 ();
 DECAPx10_ASAP7_75t_R FILLER_53_2 ();
 DECAPx10_ASAP7_75t_R FILLER_53_24 ();
 DECAPx10_ASAP7_75t_R FILLER_53_46 ();
 DECAPx4_ASAP7_75t_R FILLER_53_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_78 ();
 FILLER_ASAP7_75t_R FILLER_53_110 ();
 DECAPx2_ASAP7_75t_R FILLER_53_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_132 ();
 DECAPx1_ASAP7_75t_R FILLER_53_139 ();
 FILLER_ASAP7_75t_R FILLER_53_146 ();
 DECAPx2_ASAP7_75t_R FILLER_53_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_163 ();
 FILLER_ASAP7_75t_R FILLER_53_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_224 ();
 DECAPx1_ASAP7_75t_R FILLER_53_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_248 ();
 DECAPx2_ASAP7_75t_R FILLER_53_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_299 ();
 DECAPx6_ASAP7_75t_R FILLER_53_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_317 ();
 DECAPx10_ASAP7_75t_R FILLER_53_348 ();
 DECAPx1_ASAP7_75t_R FILLER_53_370 ();
 DECAPx2_ASAP7_75t_R FILLER_53_380 ();
 DECAPx10_ASAP7_75t_R FILLER_53_389 ();
 DECAPx2_ASAP7_75t_R FILLER_53_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_449 ();
 DECAPx4_ASAP7_75t_R FILLER_53_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_474 ();
 DECAPx2_ASAP7_75t_R FILLER_53_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_502 ();
 DECAPx2_ASAP7_75t_R FILLER_53_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_515 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_53_523 ();
 DECAPx2_ASAP7_75t_R FILLER_53_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_538 ();
 DECAPx2_ASAP7_75t_R FILLER_53_546 ();
 FILLER_ASAP7_75t_R FILLER_53_552 ();
 DECAPx1_ASAP7_75t_R FILLER_53_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_690 ();
 DECAPx6_ASAP7_75t_R FILLER_53_732 ();
 DECAPx1_ASAP7_75t_R FILLER_53_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_750 ();
 DECAPx2_ASAP7_75t_R FILLER_53_763 ();
 DECAPx10_ASAP7_75t_R FILLER_53_835 ();
 DECAPx6_ASAP7_75t_R FILLER_53_857 ();
 DECAPx10_ASAP7_75t_R FILLER_53_879 ();
 DECAPx10_ASAP7_75t_R FILLER_53_901 ();
 FILLER_ASAP7_75t_R FILLER_53_923 ();
 DECAPx2_ASAP7_75t_R FILLER_53_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_53_933 ();
 DECAPx10_ASAP7_75t_R FILLER_54_2 ();
 DECAPx10_ASAP7_75t_R FILLER_54_24 ();
 DECAPx10_ASAP7_75t_R FILLER_54_46 ();
 DECAPx10_ASAP7_75t_R FILLER_54_68 ();
 DECAPx2_ASAP7_75t_R FILLER_54_90 ();
 DECAPx2_ASAP7_75t_R FILLER_54_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_108 ();
 DECAPx2_ASAP7_75t_R FILLER_54_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_121 ();
 DECAPx10_ASAP7_75t_R FILLER_54_128 ();
 DECAPx4_ASAP7_75t_R FILLER_54_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_160 ();
 DECAPx4_ASAP7_75t_R FILLER_54_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_239 ();
 DECAPx10_ASAP7_75t_R FILLER_54_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_272 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_289 ();
 DECAPx10_ASAP7_75t_R FILLER_54_298 ();
 DECAPx2_ASAP7_75t_R FILLER_54_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_326 ();
 DECAPx10_ASAP7_75t_R FILLER_54_333 ();
 DECAPx6_ASAP7_75t_R FILLER_54_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_409 ();
 DECAPx2_ASAP7_75t_R FILLER_54_427 ();
 FILLER_ASAP7_75t_R FILLER_54_433 ();
 DECAPx1_ASAP7_75t_R FILLER_54_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_461 ();
 DECAPx10_ASAP7_75t_R FILLER_54_464 ();
 DECAPx6_ASAP7_75t_R FILLER_54_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_500 ();
 DECAPx2_ASAP7_75t_R FILLER_54_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_532 ();
 DECAPx1_ASAP7_75t_R FILLER_54_548 ();
 DECAPx10_ASAP7_75t_R FILLER_54_565 ();
 DECAPx2_ASAP7_75t_R FILLER_54_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_593 ();
 FILLER_ASAP7_75t_R FILLER_54_609 ();
 DECAPx2_ASAP7_75t_R FILLER_54_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_624 ();
 FILLER_ASAP7_75t_R FILLER_54_637 ();
 DECAPx2_ASAP7_75t_R FILLER_54_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_669 ();
 DECAPx2_ASAP7_75t_R FILLER_54_677 ();
 DECAPx1_ASAP7_75t_R FILLER_54_691 ();
 DECAPx6_ASAP7_75t_R FILLER_54_698 ();
 DECAPx10_ASAP7_75t_R FILLER_54_722 ();
 FILLER_ASAP7_75t_R FILLER_54_744 ();
 DECAPx6_ASAP7_75t_R FILLER_54_752 ();
 FILLER_ASAP7_75t_R FILLER_54_766 ();
 DECAPx6_ASAP7_75t_R FILLER_54_774 ();
 DECAPx2_ASAP7_75t_R FILLER_54_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_54_806 ();
 DECAPx2_ASAP7_75t_R FILLER_54_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_820 ();
 FILLER_ASAP7_75t_R FILLER_54_829 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_54_837 ();
 FILLER_ASAP7_75t_R FILLER_54_849 ();
 DECAPx2_ASAP7_75t_R FILLER_54_855 ();
 FILLER_ASAP7_75t_R FILLER_54_861 ();
 DECAPx10_ASAP7_75t_R FILLER_54_889 ();
 DECAPx6_ASAP7_75t_R FILLER_54_911 ();
 DECAPx1_ASAP7_75t_R FILLER_54_925 ();
 DECAPx10_ASAP7_75t_R FILLER_55_2 ();
 DECAPx10_ASAP7_75t_R FILLER_55_24 ();
 DECAPx10_ASAP7_75t_R FILLER_55_46 ();
 DECAPx10_ASAP7_75t_R FILLER_55_68 ();
 DECAPx10_ASAP7_75t_R FILLER_55_90 ();
 DECAPx10_ASAP7_75t_R FILLER_55_112 ();
 DECAPx10_ASAP7_75t_R FILLER_55_134 ();
 DECAPx6_ASAP7_75t_R FILLER_55_156 ();
 DECAPx1_ASAP7_75t_R FILLER_55_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_174 ();
 DECAPx1_ASAP7_75t_R FILLER_55_178 ();
 DECAPx4_ASAP7_75t_R FILLER_55_188 ();
 DECAPx1_ASAP7_75t_R FILLER_55_242 ();
 DECAPx2_ASAP7_75t_R FILLER_55_252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_273 ();
 DECAPx2_ASAP7_75t_R FILLER_55_279 ();
 FILLER_ASAP7_75t_R FILLER_55_285 ();
 DECAPx10_ASAP7_75t_R FILLER_55_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_335 ();
 DECAPx2_ASAP7_75t_R FILLER_55_350 ();
 FILLER_ASAP7_75t_R FILLER_55_356 ();
 DECAPx4_ASAP7_75t_R FILLER_55_364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_380 ();
 DECAPx1_ASAP7_75t_R FILLER_55_400 ();
 DECAPx4_ASAP7_75t_R FILLER_55_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_439 ();
 DECAPx1_ASAP7_75t_R FILLER_55_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_452 ();
 DECAPx10_ASAP7_75t_R FILLER_55_473 ();
 DECAPx10_ASAP7_75t_R FILLER_55_495 ();
 DECAPx10_ASAP7_75t_R FILLER_55_517 ();
 DECAPx4_ASAP7_75t_R FILLER_55_539 ();
 DECAPx10_ASAP7_75t_R FILLER_55_566 ();
 DECAPx10_ASAP7_75t_R FILLER_55_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_610 ();
 DECAPx10_ASAP7_75t_R FILLER_55_631 ();
 DECAPx10_ASAP7_75t_R FILLER_55_653 ();
 DECAPx10_ASAP7_75t_R FILLER_55_675 ();
 DECAPx10_ASAP7_75t_R FILLER_55_697 ();
 DECAPx10_ASAP7_75t_R FILLER_55_719 ();
 DECAPx10_ASAP7_75t_R FILLER_55_741 ();
 DECAPx2_ASAP7_75t_R FILLER_55_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_55_769 ();
 DECAPx10_ASAP7_75t_R FILLER_55_773 ();
 DECAPx10_ASAP7_75t_R FILLER_55_795 ();
 DECAPx1_ASAP7_75t_R FILLER_55_817 ();
 DECAPx10_ASAP7_75t_R FILLER_55_889 ();
 DECAPx2_ASAP7_75t_R FILLER_55_911 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_55_917 ();
 FILLER_ASAP7_75t_R FILLER_55_927 ();
 DECAPx10_ASAP7_75t_R FILLER_56_2 ();
 DECAPx10_ASAP7_75t_R FILLER_56_24 ();
 DECAPx10_ASAP7_75t_R FILLER_56_46 ();
 DECAPx10_ASAP7_75t_R FILLER_56_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_90 ();
 FILLER_ASAP7_75t_R FILLER_56_99 ();
 DECAPx2_ASAP7_75t_R FILLER_56_107 ();
 DECAPx4_ASAP7_75t_R FILLER_56_125 ();
 DECAPx10_ASAP7_75t_R FILLER_56_147 ();
 DECAPx10_ASAP7_75t_R FILLER_56_169 ();
 DECAPx2_ASAP7_75t_R FILLER_56_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_197 ();
 DECAPx4_ASAP7_75t_R FILLER_56_226 ();
 FILLER_ASAP7_75t_R FILLER_56_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_254 ();
 DECAPx6_ASAP7_75t_R FILLER_56_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_295 ();
 DECAPx2_ASAP7_75t_R FILLER_56_307 ();
 FILLER_ASAP7_75t_R FILLER_56_313 ();
 FILLER_ASAP7_75t_R FILLER_56_321 ();
 DECAPx4_ASAP7_75t_R FILLER_56_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_345 ();
 FILLER_ASAP7_75t_R FILLER_56_349 ();
 DECAPx4_ASAP7_75t_R FILLER_56_377 ();
 FILLER_ASAP7_75t_R FILLER_56_387 ();
 DECAPx6_ASAP7_75t_R FILLER_56_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_478 ();
 DECAPx1_ASAP7_75t_R FILLER_56_491 ();
 DECAPx10_ASAP7_75t_R FILLER_56_501 ();
 DECAPx10_ASAP7_75t_R FILLER_56_523 ();
 DECAPx10_ASAP7_75t_R FILLER_56_545 ();
 DECAPx6_ASAP7_75t_R FILLER_56_567 ();
 DECAPx2_ASAP7_75t_R FILLER_56_581 ();
 DECAPx10_ASAP7_75t_R FILLER_56_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_616 ();
 DECAPx6_ASAP7_75t_R FILLER_56_623 ();
 DECAPx2_ASAP7_75t_R FILLER_56_637 ();
 DECAPx4_ASAP7_75t_R FILLER_56_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_656 ();
 DECAPx10_ASAP7_75t_R FILLER_56_683 ();
 DECAPx6_ASAP7_75t_R FILLER_56_705 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_719 ();
 DECAPx1_ASAP7_75t_R FILLER_56_729 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_760 ();
 DECAPx10_ASAP7_75t_R FILLER_56_770 ();
 DECAPx10_ASAP7_75t_R FILLER_56_792 ();
 DECAPx10_ASAP7_75t_R FILLER_56_814 ();
 DECAPx2_ASAP7_75t_R FILLER_56_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_56_873 ();
 DECAPx2_ASAP7_75t_R FILLER_56_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_56_906 ();
 DECAPx10_ASAP7_75t_R FILLER_57_2 ();
 DECAPx10_ASAP7_75t_R FILLER_57_24 ();
 DECAPx10_ASAP7_75t_R FILLER_57_46 ();
 DECAPx6_ASAP7_75t_R FILLER_57_68 ();
 DECAPx1_ASAP7_75t_R FILLER_57_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_86 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_113 ();
 FILLER_ASAP7_75t_R FILLER_57_124 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_155 ();
 DECAPx10_ASAP7_75t_R FILLER_57_170 ();
 DECAPx4_ASAP7_75t_R FILLER_57_192 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_202 ();
 FILLER_ASAP7_75t_R FILLER_57_211 ();
 DECAPx6_ASAP7_75t_R FILLER_57_216 ();
 FILLER_ASAP7_75t_R FILLER_57_230 ();
 DECAPx10_ASAP7_75t_R FILLER_57_258 ();
 FILLER_ASAP7_75t_R FILLER_57_280 ();
 DECAPx6_ASAP7_75t_R FILLER_57_290 ();
 FILLER_ASAP7_75t_R FILLER_57_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_365 ();
 DECAPx6_ASAP7_75t_R FILLER_57_378 ();
 DECAPx2_ASAP7_75t_R FILLER_57_392 ();
 DECAPx2_ASAP7_75t_R FILLER_57_404 ();
 DECAPx2_ASAP7_75t_R FILLER_57_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_462 ();
 FILLER_ASAP7_75t_R FILLER_57_482 ();
 FILLER_ASAP7_75t_R FILLER_57_492 ();
 FILLER_ASAP7_75t_R FILLER_57_502 ();
 DECAPx2_ASAP7_75t_R FILLER_57_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_516 ();
 FILLER_ASAP7_75t_R FILLER_57_523 ();
 FILLER_ASAP7_75t_R FILLER_57_536 ();
 DECAPx6_ASAP7_75t_R FILLER_57_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_558 ();
 DECAPx4_ASAP7_75t_R FILLER_57_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_584 ();
 DECAPx6_ASAP7_75t_R FILLER_57_607 ();
 DECAPx2_ASAP7_75t_R FILLER_57_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_627 ();
 DECAPx4_ASAP7_75t_R FILLER_57_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_664 ();
 DECAPx1_ASAP7_75t_R FILLER_57_680 ();
 DECAPx2_ASAP7_75t_R FILLER_57_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_57_712 ();
 DECAPx4_ASAP7_75t_R FILLER_57_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_751 ();
 FILLER_ASAP7_75t_R FILLER_57_772 ();
 DECAPx6_ASAP7_75t_R FILLER_57_789 ();
 FILLER_ASAP7_75t_R FILLER_57_803 ();
 DECAPx10_ASAP7_75t_R FILLER_57_831 ();
 DECAPx6_ASAP7_75t_R FILLER_57_853 ();
 DECAPx2_ASAP7_75t_R FILLER_57_867 ();
 DECAPx6_ASAP7_75t_R FILLER_57_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_57_900 ();
 FILLER_ASAP7_75t_R FILLER_57_927 ();
 DECAPx10_ASAP7_75t_R FILLER_58_2 ();
 DECAPx10_ASAP7_75t_R FILLER_58_24 ();
 DECAPx10_ASAP7_75t_R FILLER_58_46 ();
 DECAPx6_ASAP7_75t_R FILLER_58_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_82 ();
 FILLER_ASAP7_75t_R FILLER_58_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_122 ();
 DECAPx4_ASAP7_75t_R FILLER_58_131 ();
 DECAPx2_ASAP7_75t_R FILLER_58_144 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_150 ();
 DECAPx6_ASAP7_75t_R FILLER_58_193 ();
 DECAPx1_ASAP7_75t_R FILLER_58_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_211 ();
 DECAPx10_ASAP7_75t_R FILLER_58_218 ();
 DECAPx2_ASAP7_75t_R FILLER_58_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_246 ();
 DECAPx4_ASAP7_75t_R FILLER_58_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_260 ();
 DECAPx6_ASAP7_75t_R FILLER_58_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_283 ();
 DECAPx1_ASAP7_75t_R FILLER_58_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_314 ();
 DECAPx6_ASAP7_75t_R FILLER_58_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_345 ();
 DECAPx10_ASAP7_75t_R FILLER_58_355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_387 ();
 DECAPx10_ASAP7_75t_R FILLER_58_393 ();
 DECAPx4_ASAP7_75t_R FILLER_58_415 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_425 ();
 DECAPx1_ASAP7_75t_R FILLER_58_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_461 ();
 DECAPx2_ASAP7_75t_R FILLER_58_484 ();
 FILLER_ASAP7_75t_R FILLER_58_490 ();
 DECAPx2_ASAP7_75t_R FILLER_58_498 ();
 FILLER_ASAP7_75t_R FILLER_58_504 ();
 DECAPx4_ASAP7_75t_R FILLER_58_536 ();
 FILLER_ASAP7_75t_R FILLER_58_546 ();
 DECAPx2_ASAP7_75t_R FILLER_58_554 ();
 FILLER_ASAP7_75t_R FILLER_58_560 ();
 DECAPx1_ASAP7_75t_R FILLER_58_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_598 ();
 DECAPx6_ASAP7_75t_R FILLER_58_607 ();
 FILLER_ASAP7_75t_R FILLER_58_621 ();
 DECAPx2_ASAP7_75t_R FILLER_58_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_676 ();
 FILLER_ASAP7_75t_R FILLER_58_694 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_737 ();
 DECAPx2_ASAP7_75t_R FILLER_58_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_763 ();
 DECAPx2_ASAP7_75t_R FILLER_58_770 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_58_776 ();
 DECAPx10_ASAP7_75t_R FILLER_58_826 ();
 DECAPx10_ASAP7_75t_R FILLER_58_848 ();
 DECAPx10_ASAP7_75t_R FILLER_58_870 ();
 DECAPx2_ASAP7_75t_R FILLER_58_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_58_898 ();
 DECAPx1_ASAP7_75t_R FILLER_58_930 ();
 DECAPx10_ASAP7_75t_R FILLER_59_2 ();
 DECAPx10_ASAP7_75t_R FILLER_59_24 ();
 DECAPx10_ASAP7_75t_R FILLER_59_46 ();
 DECAPx6_ASAP7_75t_R FILLER_59_68 ();
 DECAPx2_ASAP7_75t_R FILLER_59_82 ();
 FILLER_ASAP7_75t_R FILLER_59_100 ();
 DECAPx1_ASAP7_75t_R FILLER_59_108 ();
 DECAPx10_ASAP7_75t_R FILLER_59_118 ();
 DECAPx4_ASAP7_75t_R FILLER_59_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_150 ();
 DECAPx1_ASAP7_75t_R FILLER_59_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_208 ();
 FILLER_ASAP7_75t_R FILLER_59_235 ();
 DECAPx2_ASAP7_75t_R FILLER_59_245 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_251 ();
 DECAPx2_ASAP7_75t_R FILLER_59_290 ();
 DECAPx1_ASAP7_75t_R FILLER_59_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_327 ();
 DECAPx10_ASAP7_75t_R FILLER_59_346 ();
 DECAPx4_ASAP7_75t_R FILLER_59_368 ();
 DECAPx1_ASAP7_75t_R FILLER_59_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_414 ();
 DECAPx6_ASAP7_75t_R FILLER_59_422 ();
 DECAPx2_ASAP7_75t_R FILLER_59_436 ();
 DECAPx10_ASAP7_75t_R FILLER_59_472 ();
 DECAPx6_ASAP7_75t_R FILLER_59_494 ();
 DECAPx2_ASAP7_75t_R FILLER_59_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_514 ();
 DECAPx4_ASAP7_75t_R FILLER_59_521 ();
 DECAPx2_ASAP7_75t_R FILLER_59_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_592 ();
 DECAPx1_ASAP7_75t_R FILLER_59_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_640 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_654 ();
 DECAPx4_ASAP7_75t_R FILLER_59_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_697 ();
 DECAPx1_ASAP7_75t_R FILLER_59_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_730 ();
 DECAPx6_ASAP7_75t_R FILLER_59_734 ();
 FILLER_ASAP7_75t_R FILLER_59_748 ();
 DECAPx6_ASAP7_75t_R FILLER_59_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_774 ();
 DECAPx1_ASAP7_75t_R FILLER_59_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_809 ();
 DECAPx2_ASAP7_75t_R FILLER_59_817 ();
 FILLER_ASAP7_75t_R FILLER_59_823 ();
 DECAPx10_ASAP7_75t_R FILLER_59_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_59_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_858 ();
 DECAPx10_ASAP7_75t_R FILLER_59_864 ();
 DECAPx6_ASAP7_75t_R FILLER_59_886 ();
 DECAPx1_ASAP7_75t_R FILLER_59_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_59_914 ();
 FILLER_ASAP7_75t_R FILLER_59_932 ();
 DECAPx10_ASAP7_75t_R FILLER_60_2 ();
 DECAPx10_ASAP7_75t_R FILLER_60_24 ();
 DECAPx10_ASAP7_75t_R FILLER_60_46 ();
 DECAPx10_ASAP7_75t_R FILLER_60_68 ();
 DECAPx10_ASAP7_75t_R FILLER_60_90 ();
 DECAPx6_ASAP7_75t_R FILLER_60_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_147 ();
 DECAPx4_ASAP7_75t_R FILLER_60_157 ();
 DECAPx1_ASAP7_75t_R FILLER_60_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_192 ();
 FILLER_ASAP7_75t_R FILLER_60_209 ();
 DECAPx2_ASAP7_75t_R FILLER_60_217 ();
 DECAPx1_ASAP7_75t_R FILLER_60_254 ();
 FILLER_ASAP7_75t_R FILLER_60_264 ();
 DECAPx1_ASAP7_75t_R FILLER_60_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_289 ();
 DECAPx2_ASAP7_75t_R FILLER_60_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_305 ();
 DECAPx1_ASAP7_75t_R FILLER_60_318 ();
 DECAPx2_ASAP7_75t_R FILLER_60_329 ();
 DECAPx6_ASAP7_75t_R FILLER_60_349 ();
 DECAPx2_ASAP7_75t_R FILLER_60_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_376 ();
 FILLER_ASAP7_75t_R FILLER_60_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_461 ();
 DECAPx2_ASAP7_75t_R FILLER_60_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_470 ();
 DECAPx2_ASAP7_75t_R FILLER_60_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_487 ();
 DECAPx10_ASAP7_75t_R FILLER_60_511 ();
 DECAPx2_ASAP7_75t_R FILLER_60_533 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_565 ();
 DECAPx1_ASAP7_75t_R FILLER_60_572 ();
 DECAPx2_ASAP7_75t_R FILLER_60_582 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_588 ();
 DECAPx1_ASAP7_75t_R FILLER_60_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_601 ();
 FILLER_ASAP7_75t_R FILLER_60_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_656 ();
 FILLER_ASAP7_75t_R FILLER_60_678 ();
 DECAPx6_ASAP7_75t_R FILLER_60_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_702 ();
 DECAPx10_ASAP7_75t_R FILLER_60_709 ();
 DECAPx10_ASAP7_75t_R FILLER_60_731 ();
 DECAPx2_ASAP7_75t_R FILLER_60_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_765 ();
 DECAPx2_ASAP7_75t_R FILLER_60_769 ();
 DECAPx2_ASAP7_75t_R FILLER_60_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_798 ();
 DECAPx1_ASAP7_75t_R FILLER_60_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_819 ();
 DECAPx1_ASAP7_75t_R FILLER_60_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_60_850 ();
 DECAPx10_ASAP7_75t_R FILLER_60_881 ();
 DECAPx2_ASAP7_75t_R FILLER_60_903 ();
 FILLER_ASAP7_75t_R FILLER_60_909 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_60_931 ();
 DECAPx10_ASAP7_75t_R FILLER_61_2 ();
 DECAPx10_ASAP7_75t_R FILLER_61_24 ();
 DECAPx10_ASAP7_75t_R FILLER_61_46 ();
 DECAPx10_ASAP7_75t_R FILLER_61_68 ();
 DECAPx6_ASAP7_75t_R FILLER_61_90 ();
 DECAPx2_ASAP7_75t_R FILLER_61_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_110 ();
 DECAPx4_ASAP7_75t_R FILLER_61_118 ();
 DECAPx2_ASAP7_75t_R FILLER_61_154 ();
 DECAPx6_ASAP7_75t_R FILLER_61_166 ();
 DECAPx2_ASAP7_75t_R FILLER_61_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_190 ();
 FILLER_ASAP7_75t_R FILLER_61_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_228 ();
 FILLER_ASAP7_75t_R FILLER_61_239 ();
 DECAPx1_ASAP7_75t_R FILLER_61_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_267 ();
 DECAPx4_ASAP7_75t_R FILLER_61_271 ();
 FILLER_ASAP7_75t_R FILLER_61_281 ();
 DECAPx10_ASAP7_75t_R FILLER_61_309 ();
 DECAPx10_ASAP7_75t_R FILLER_61_331 ();
 DECAPx1_ASAP7_75t_R FILLER_61_353 ();
 DECAPx1_ASAP7_75t_R FILLER_61_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_443 ();
 DECAPx4_ASAP7_75t_R FILLER_61_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_491 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_499 ();
 DECAPx6_ASAP7_75t_R FILLER_61_512 ();
 DECAPx1_ASAP7_75t_R FILLER_61_526 ();
 DECAPx10_ASAP7_75t_R FILLER_61_540 ();
 DECAPx10_ASAP7_75t_R FILLER_61_562 ();
 DECAPx10_ASAP7_75t_R FILLER_61_584 ();
 DECAPx1_ASAP7_75t_R FILLER_61_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_610 ();
 DECAPx6_ASAP7_75t_R FILLER_61_617 ();
 DECAPx2_ASAP7_75t_R FILLER_61_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_637 ();
 DECAPx4_ASAP7_75t_R FILLER_61_644 ();
 FILLER_ASAP7_75t_R FILLER_61_654 ();
 DECAPx10_ASAP7_75t_R FILLER_61_665 ();
 DECAPx10_ASAP7_75t_R FILLER_61_687 ();
 DECAPx10_ASAP7_75t_R FILLER_61_709 ();
 FILLER_ASAP7_75t_R FILLER_61_731 ();
 DECAPx6_ASAP7_75t_R FILLER_61_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_750 ();
 DECAPx4_ASAP7_75t_R FILLER_61_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_778 ();
 DECAPx4_ASAP7_75t_R FILLER_61_785 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_61_795 ();
 DECAPx2_ASAP7_75t_R FILLER_61_804 ();
 FILLER_ASAP7_75t_R FILLER_61_810 ();
 FILLER_ASAP7_75t_R FILLER_61_818 ();
 FILLER_ASAP7_75t_R FILLER_61_838 ();
 DECAPx6_ASAP7_75t_R FILLER_61_885 ();
 DECAPx1_ASAP7_75t_R FILLER_61_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_61_924 ();
 FILLER_ASAP7_75t_R FILLER_61_932 ();
 DECAPx10_ASAP7_75t_R FILLER_62_2 ();
 DECAPx10_ASAP7_75t_R FILLER_62_24 ();
 DECAPx10_ASAP7_75t_R FILLER_62_46 ();
 DECAPx10_ASAP7_75t_R FILLER_62_68 ();
 DECAPx2_ASAP7_75t_R FILLER_62_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_96 ();
 DECAPx2_ASAP7_75t_R FILLER_62_125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_131 ();
 FILLER_ASAP7_75t_R FILLER_62_140 ();
 DECAPx1_ASAP7_75t_R FILLER_62_151 ();
 DECAPx10_ASAP7_75t_R FILLER_62_172 ();
 DECAPx4_ASAP7_75t_R FILLER_62_194 ();
 FILLER_ASAP7_75t_R FILLER_62_204 ();
 DECAPx1_ASAP7_75t_R FILLER_62_212 ();
 DECAPx2_ASAP7_75t_R FILLER_62_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_225 ();
 FILLER_ASAP7_75t_R FILLER_62_246 ();
 DECAPx10_ASAP7_75t_R FILLER_62_255 ();
 DECAPx4_ASAP7_75t_R FILLER_62_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_294 ();
 DECAPx10_ASAP7_75t_R FILLER_62_304 ();
 DECAPx6_ASAP7_75t_R FILLER_62_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_347 ();
 DECAPx2_ASAP7_75t_R FILLER_62_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_386 ();
 DECAPx2_ASAP7_75t_R FILLER_62_415 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_421 ();
 FILLER_ASAP7_75t_R FILLER_62_427 ();
 FILLER_ASAP7_75t_R FILLER_62_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_464 ();
 FILLER_ASAP7_75t_R FILLER_62_483 ();
 DECAPx1_ASAP7_75t_R FILLER_62_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_506 ();
 DECAPx4_ASAP7_75t_R FILLER_62_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_537 ();
 DECAPx10_ASAP7_75t_R FILLER_62_547 ();
 DECAPx4_ASAP7_75t_R FILLER_62_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_579 ();
 DECAPx10_ASAP7_75t_R FILLER_62_587 ();
 DECAPx2_ASAP7_75t_R FILLER_62_609 ();
 FILLER_ASAP7_75t_R FILLER_62_615 ();
 DECAPx2_ASAP7_75t_R FILLER_62_623 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_629 ();
 DECAPx2_ASAP7_75t_R FILLER_62_638 ();
 FILLER_ASAP7_75t_R FILLER_62_644 ();
 DECAPx10_ASAP7_75t_R FILLER_62_649 ();
 DECAPx10_ASAP7_75t_R FILLER_62_671 ();
 DECAPx6_ASAP7_75t_R FILLER_62_693 ();
 DECAPx1_ASAP7_75t_R FILLER_62_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_711 ();
 FILLER_ASAP7_75t_R FILLER_62_744 ();
 DECAPx1_ASAP7_75t_R FILLER_62_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_756 ();
 DECAPx10_ASAP7_75t_R FILLER_62_763 ();
 DECAPx10_ASAP7_75t_R FILLER_62_785 ();
 DECAPx10_ASAP7_75t_R FILLER_62_807 ();
 DECAPx2_ASAP7_75t_R FILLER_62_829 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_835 ();
 DECAPx2_ASAP7_75t_R FILLER_62_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_874 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_62_898 ();
 DECAPx2_ASAP7_75t_R FILLER_62_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_62_933 ();
 DECAPx10_ASAP7_75t_R FILLER_63_2 ();
 DECAPx10_ASAP7_75t_R FILLER_63_24 ();
 DECAPx10_ASAP7_75t_R FILLER_63_46 ();
 DECAPx10_ASAP7_75t_R FILLER_63_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_90 ();
 DECAPx2_ASAP7_75t_R FILLER_63_138 ();
 FILLER_ASAP7_75t_R FILLER_63_144 ();
 DECAPx10_ASAP7_75t_R FILLER_63_152 ();
 DECAPx10_ASAP7_75t_R FILLER_63_174 ();
 DECAPx4_ASAP7_75t_R FILLER_63_196 ();
 DECAPx4_ASAP7_75t_R FILLER_63_212 ();
 FILLER_ASAP7_75t_R FILLER_63_222 ();
 DECAPx10_ASAP7_75t_R FILLER_63_236 ();
 DECAPx2_ASAP7_75t_R FILLER_63_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_270 ();
 DECAPx2_ASAP7_75t_R FILLER_63_279 ();
 DECAPx10_ASAP7_75t_R FILLER_63_290 ();
 DECAPx10_ASAP7_75t_R FILLER_63_312 ();
 DECAPx1_ASAP7_75t_R FILLER_63_360 ();
 DECAPx10_ASAP7_75t_R FILLER_63_376 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_398 ();
 DECAPx4_ASAP7_75t_R FILLER_63_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_417 ();
 DECAPx4_ASAP7_75t_R FILLER_63_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_434 ();
 DECAPx4_ASAP7_75t_R FILLER_63_440 ();
 FILLER_ASAP7_75t_R FILLER_63_450 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_473 ();
 DECAPx4_ASAP7_75t_R FILLER_63_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_504 ();
 FILLER_ASAP7_75t_R FILLER_63_532 ();
 FILLER_ASAP7_75t_R FILLER_63_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_550 ();
 DECAPx1_ASAP7_75t_R FILLER_63_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_565 ();
 DECAPx2_ASAP7_75t_R FILLER_63_572 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_578 ();
 DECAPx1_ASAP7_75t_R FILLER_63_607 ();
 FILLER_ASAP7_75t_R FILLER_63_617 ();
 DECAPx2_ASAP7_75t_R FILLER_63_626 ();
 FILLER_ASAP7_75t_R FILLER_63_632 ();
 DECAPx2_ASAP7_75t_R FILLER_63_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_665 ();
 DECAPx1_ASAP7_75t_R FILLER_63_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_673 ();
 DECAPx6_ASAP7_75t_R FILLER_63_710 ();
 DECAPx10_ASAP7_75t_R FILLER_63_730 ();
 DECAPx4_ASAP7_75t_R FILLER_63_752 ();
 FILLER_ASAP7_75t_R FILLER_63_762 ();
 DECAPx6_ASAP7_75t_R FILLER_63_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_791 ();
 DECAPx6_ASAP7_75t_R FILLER_63_801 ();
 DECAPx2_ASAP7_75t_R FILLER_63_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_821 ();
 DECAPx10_ASAP7_75t_R FILLER_63_848 ();
 FILLER_ASAP7_75t_R FILLER_63_870 ();
 DECAPx10_ASAP7_75t_R FILLER_63_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_63_907 ();
 DECAPx1_ASAP7_75t_R FILLER_63_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_924 ();
 DECAPx2_ASAP7_75t_R FILLER_63_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_63_933 ();
 DECAPx10_ASAP7_75t_R FILLER_64_2 ();
 DECAPx10_ASAP7_75t_R FILLER_64_24 ();
 DECAPx10_ASAP7_75t_R FILLER_64_46 ();
 DECAPx6_ASAP7_75t_R FILLER_64_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_108 ();
 FILLER_ASAP7_75t_R FILLER_64_125 ();
 FILLER_ASAP7_75t_R FILLER_64_142 ();
 DECAPx1_ASAP7_75t_R FILLER_64_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_151 ();
 FILLER_ASAP7_75t_R FILLER_64_158 ();
 DECAPx1_ASAP7_75t_R FILLER_64_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_176 ();
 DECAPx1_ASAP7_75t_R FILLER_64_189 ();
 DECAPx10_ASAP7_75t_R FILLER_64_199 ();
 DECAPx2_ASAP7_75t_R FILLER_64_233 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_248 ();
 DECAPx4_ASAP7_75t_R FILLER_64_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_297 ();
 DECAPx4_ASAP7_75t_R FILLER_64_304 ();
 FILLER_ASAP7_75t_R FILLER_64_314 ();
 DECAPx2_ASAP7_75t_R FILLER_64_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_336 ();
 DECAPx1_ASAP7_75t_R FILLER_64_343 ();
 DECAPx10_ASAP7_75t_R FILLER_64_356 ();
 DECAPx10_ASAP7_75t_R FILLER_64_378 ();
 DECAPx6_ASAP7_75t_R FILLER_64_400 ();
 FILLER_ASAP7_75t_R FILLER_64_414 ();
 DECAPx4_ASAP7_75t_R FILLER_64_452 ();
 FILLER_ASAP7_75t_R FILLER_64_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_473 ();
 DECAPx10_ASAP7_75t_R FILLER_64_480 ();
 DECAPx1_ASAP7_75t_R FILLER_64_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_506 ();
 DECAPx10_ASAP7_75t_R FILLER_64_513 ();
 DECAPx6_ASAP7_75t_R FILLER_64_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_64_549 ();
 DECAPx1_ASAP7_75t_R FILLER_64_590 ();
 DECAPx1_ASAP7_75t_R FILLER_64_614 ();
 DECAPx6_ASAP7_75t_R FILLER_64_638 ();
 DECAPx1_ASAP7_75t_R FILLER_64_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_760 ();
 DECAPx6_ASAP7_75t_R FILLER_64_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_64_836 ();
 FILLER_ASAP7_75t_R FILLER_64_840 ();
 DECAPx10_ASAP7_75t_R FILLER_64_850 ();
 DECAPx10_ASAP7_75t_R FILLER_64_872 ();
 DECAPx10_ASAP7_75t_R FILLER_64_894 ();
 DECAPx6_ASAP7_75t_R FILLER_64_916 ();
 DECAPx1_ASAP7_75t_R FILLER_64_930 ();
 DECAPx10_ASAP7_75t_R FILLER_65_2 ();
 DECAPx10_ASAP7_75t_R FILLER_65_24 ();
 DECAPx10_ASAP7_75t_R FILLER_65_46 ();
 DECAPx10_ASAP7_75t_R FILLER_65_68 ();
 DECAPx2_ASAP7_75t_R FILLER_65_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_96 ();
 FILLER_ASAP7_75t_R FILLER_65_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_118 ();
 DECAPx6_ASAP7_75t_R FILLER_65_217 ();
 DECAPx2_ASAP7_75t_R FILLER_65_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_270 ();
 DECAPx1_ASAP7_75t_R FILLER_65_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_319 ();
 DECAPx2_ASAP7_75t_R FILLER_65_356 ();
 FILLER_ASAP7_75t_R FILLER_65_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_371 ();
 DECAPx10_ASAP7_75t_R FILLER_65_386 ();
 DECAPx10_ASAP7_75t_R FILLER_65_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_457 ();
 DECAPx10_ASAP7_75t_R FILLER_65_473 ();
 DECAPx10_ASAP7_75t_R FILLER_65_495 ();
 DECAPx10_ASAP7_75t_R FILLER_65_517 ();
 DECAPx6_ASAP7_75t_R FILLER_65_539 ();
 DECAPx2_ASAP7_75t_R FILLER_65_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_567 ();
 DECAPx1_ASAP7_75t_R FILLER_65_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_578 ();
 DECAPx2_ASAP7_75t_R FILLER_65_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_590 ();
 DECAPx2_ASAP7_75t_R FILLER_65_602 ();
 FILLER_ASAP7_75t_R FILLER_65_608 ();
 DECAPx2_ASAP7_75t_R FILLER_65_616 ();
 FILLER_ASAP7_75t_R FILLER_65_622 ();
 DECAPx4_ASAP7_75t_R FILLER_65_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_656 ();
 DECAPx6_ASAP7_75t_R FILLER_65_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_65_685 ();
 DECAPx4_ASAP7_75t_R FILLER_65_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_704 ();
 DECAPx2_ASAP7_75t_R FILLER_65_713 ();
 FILLER_ASAP7_75t_R FILLER_65_727 ();
 DECAPx1_ASAP7_75t_R FILLER_65_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_741 ();
 DECAPx6_ASAP7_75t_R FILLER_65_750 ();
 FILLER_ASAP7_75t_R FILLER_65_773 ();
 DECAPx1_ASAP7_75t_R FILLER_65_778 ();
 DECAPx2_ASAP7_75t_R FILLER_65_785 ();
 FILLER_ASAP7_75t_R FILLER_65_791 ();
 DECAPx1_ASAP7_75t_R FILLER_65_858 ();
 DECAPx2_ASAP7_75t_R FILLER_65_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_882 ();
 DECAPx10_ASAP7_75t_R FILLER_65_889 ();
 DECAPx6_ASAP7_75t_R FILLER_65_911 ();
 DECAPx2_ASAP7_75t_R FILLER_65_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_65_933 ();
 DECAPx10_ASAP7_75t_R FILLER_66_2 ();
 DECAPx10_ASAP7_75t_R FILLER_66_24 ();
 DECAPx10_ASAP7_75t_R FILLER_66_46 ();
 DECAPx10_ASAP7_75t_R FILLER_66_68 ();
 DECAPx4_ASAP7_75t_R FILLER_66_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_100 ();
 DECAPx2_ASAP7_75t_R FILLER_66_106 ();
 DECAPx10_ASAP7_75t_R FILLER_66_118 ();
 DECAPx6_ASAP7_75t_R FILLER_66_140 ();
 FILLER_ASAP7_75t_R FILLER_66_154 ();
 DECAPx2_ASAP7_75t_R FILLER_66_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_184 ();
 DECAPx1_ASAP7_75t_R FILLER_66_188 ();
 DECAPx1_ASAP7_75t_R FILLER_66_195 ();
 DECAPx2_ASAP7_75t_R FILLER_66_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_244 ();
 FILLER_ASAP7_75t_R FILLER_66_268 ();
 DECAPx2_ASAP7_75t_R FILLER_66_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_293 ();
 FILLER_ASAP7_75t_R FILLER_66_300 ();
 FILLER_ASAP7_75t_R FILLER_66_319 ();
 DECAPx1_ASAP7_75t_R FILLER_66_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_332 ();
 DECAPx2_ASAP7_75t_R FILLER_66_339 ();
 DECAPx6_ASAP7_75t_R FILLER_66_348 ();
 DECAPx1_ASAP7_75t_R FILLER_66_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_429 ();
 DECAPx1_ASAP7_75t_R FILLER_66_458 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_493 ();
 DECAPx10_ASAP7_75t_R FILLER_66_502 ();
 DECAPx6_ASAP7_75t_R FILLER_66_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_538 ();
 DECAPx1_ASAP7_75t_R FILLER_66_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_550 ();
 DECAPx6_ASAP7_75t_R FILLER_66_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_571 ();
 DECAPx2_ASAP7_75t_R FILLER_66_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_605 ();
 DECAPx10_ASAP7_75t_R FILLER_66_612 ();
 DECAPx6_ASAP7_75t_R FILLER_66_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_648 ();
 DECAPx10_ASAP7_75t_R FILLER_66_659 ();
 DECAPx4_ASAP7_75t_R FILLER_66_681 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_691 ();
 DECAPx10_ASAP7_75t_R FILLER_66_701 ();
 DECAPx2_ASAP7_75t_R FILLER_66_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_729 ();
 FILLER_ASAP7_75t_R FILLER_66_736 ();
 DECAPx2_ASAP7_75t_R FILLER_66_744 ();
 FILLER_ASAP7_75t_R FILLER_66_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_66_764 ();
 DECAPx4_ASAP7_75t_R FILLER_66_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_66_803 ();
 FILLER_ASAP7_75t_R FILLER_66_807 ();
 FILLER_ASAP7_75t_R FILLER_66_822 ();
 DECAPx1_ASAP7_75t_R FILLER_66_836 ();
 DECAPx6_ASAP7_75t_R FILLER_66_852 ();
 FILLER_ASAP7_75t_R FILLER_66_866 ();
 DECAPx10_ASAP7_75t_R FILLER_66_896 ();
 DECAPx6_ASAP7_75t_R FILLER_66_918 ();
 FILLER_ASAP7_75t_R FILLER_66_932 ();
 DECAPx10_ASAP7_75t_R FILLER_67_2 ();
 DECAPx10_ASAP7_75t_R FILLER_67_24 ();
 DECAPx10_ASAP7_75t_R FILLER_67_46 ();
 DECAPx10_ASAP7_75t_R FILLER_67_68 ();
 DECAPx10_ASAP7_75t_R FILLER_67_90 ();
 DECAPx6_ASAP7_75t_R FILLER_67_112 ();
 DECAPx2_ASAP7_75t_R FILLER_67_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_132 ();
 DECAPx10_ASAP7_75t_R FILLER_67_139 ();
 DECAPx6_ASAP7_75t_R FILLER_67_161 ();
 DECAPx2_ASAP7_75t_R FILLER_67_175 ();
 DECAPx10_ASAP7_75t_R FILLER_67_187 ();
 DECAPx1_ASAP7_75t_R FILLER_67_209 ();
 DECAPx4_ASAP7_75t_R FILLER_67_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_226 ();
 DECAPx6_ASAP7_75t_R FILLER_67_253 ();
 DECAPx2_ASAP7_75t_R FILLER_67_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_273 ();
 DECAPx2_ASAP7_75t_R FILLER_67_310 ();
 FILLER_ASAP7_75t_R FILLER_67_316 ();
 DECAPx10_ASAP7_75t_R FILLER_67_324 ();
 FILLER_ASAP7_75t_R FILLER_67_346 ();
 DECAPx1_ASAP7_75t_R FILLER_67_360 ();
 DECAPx1_ASAP7_75t_R FILLER_67_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_417 ();
 DECAPx6_ASAP7_75t_R FILLER_67_457 ();
 FILLER_ASAP7_75t_R FILLER_67_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_513 ();
 DECAPx1_ASAP7_75t_R FILLER_67_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_528 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_537 ();
 DECAPx10_ASAP7_75t_R FILLER_67_574 ();
 DECAPx10_ASAP7_75t_R FILLER_67_596 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_67_618 ();
 FILLER_ASAP7_75t_R FILLER_67_634 ();
 DECAPx10_ASAP7_75t_R FILLER_67_642 ();
 DECAPx6_ASAP7_75t_R FILLER_67_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_678 ();
 DECAPx1_ASAP7_75t_R FILLER_67_682 ();
 DECAPx6_ASAP7_75t_R FILLER_67_696 ();
 DECAPx10_ASAP7_75t_R FILLER_67_719 ();
 DECAPx10_ASAP7_75t_R FILLER_67_741 ();
 DECAPx2_ASAP7_75t_R FILLER_67_763 ();
 DECAPx10_ASAP7_75t_R FILLER_67_782 ();
 DECAPx6_ASAP7_75t_R FILLER_67_804 ();
 FILLER_ASAP7_75t_R FILLER_67_818 ();
 DECAPx10_ASAP7_75t_R FILLER_67_823 ();
 DECAPx4_ASAP7_75t_R FILLER_67_845 ();
 DECAPx10_ASAP7_75t_R FILLER_67_861 ();
 DECAPx6_ASAP7_75t_R FILLER_67_883 ();
 DECAPx2_ASAP7_75t_R FILLER_67_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_67_903 ();
 DECAPx6_ASAP7_75t_R FILLER_67_907 ();
 DECAPx1_ASAP7_75t_R FILLER_67_921 ();
 FILLER_ASAP7_75t_R FILLER_67_927 ();
 DECAPx10_ASAP7_75t_R FILLER_68_2 ();
 DECAPx10_ASAP7_75t_R FILLER_68_24 ();
 DECAPx10_ASAP7_75t_R FILLER_68_46 ();
 DECAPx10_ASAP7_75t_R FILLER_68_68 ();
 DECAPx10_ASAP7_75t_R FILLER_68_90 ();
 DECAPx2_ASAP7_75t_R FILLER_68_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_118 ();
 DECAPx10_ASAP7_75t_R FILLER_68_143 ();
 DECAPx2_ASAP7_75t_R FILLER_68_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_171 ();
 DECAPx4_ASAP7_75t_R FILLER_68_200 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_210 ();
 DECAPx10_ASAP7_75t_R FILLER_68_219 ();
 DECAPx10_ASAP7_75t_R FILLER_68_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_266 ();
 DECAPx1_ASAP7_75t_R FILLER_68_275 ();
 DECAPx2_ASAP7_75t_R FILLER_68_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_308 ();
 DECAPx2_ASAP7_75t_R FILLER_68_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_321 ();
 DECAPx2_ASAP7_75t_R FILLER_68_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_335 ();
 DECAPx1_ASAP7_75t_R FILLER_68_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_367 ();
 DECAPx2_ASAP7_75t_R FILLER_68_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_379 ();
 DECAPx6_ASAP7_75t_R FILLER_68_386 ();
 DECAPx2_ASAP7_75t_R FILLER_68_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_406 ();
 DECAPx6_ASAP7_75t_R FILLER_68_419 ();
 DECAPx2_ASAP7_75t_R FILLER_68_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_439 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_448 ();
 DECAPx2_ASAP7_75t_R FILLER_68_456 ();
 DECAPx2_ASAP7_75t_R FILLER_68_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_496 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_549 ();
 DECAPx2_ASAP7_75t_R FILLER_68_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_575 ();
 DECAPx4_ASAP7_75t_R FILLER_68_584 ();
 DECAPx2_ASAP7_75t_R FILLER_68_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_620 ();
 DECAPx2_ASAP7_75t_R FILLER_68_647 ();
 DECAPx4_ASAP7_75t_R FILLER_68_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_692 ();
 FILLER_ASAP7_75t_R FILLER_68_704 ();
 DECAPx2_ASAP7_75t_R FILLER_68_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_745 ();
 DECAPx6_ASAP7_75t_R FILLER_68_752 ();
 FILLER_ASAP7_75t_R FILLER_68_766 ();
 DECAPx2_ASAP7_75t_R FILLER_68_774 ();
 FILLER_ASAP7_75t_R FILLER_68_780 ();
 DECAPx1_ASAP7_75t_R FILLER_68_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_793 ();
 DECAPx2_ASAP7_75t_R FILLER_68_801 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_68_807 ();
 DECAPx10_ASAP7_75t_R FILLER_68_813 ();
 DECAPx6_ASAP7_75t_R FILLER_68_835 ();
 DECAPx1_ASAP7_75t_R FILLER_68_849 ();
 DECAPx6_ASAP7_75t_R FILLER_68_870 ();
 DECAPx2_ASAP7_75t_R FILLER_68_884 ();
 DECAPx6_ASAP7_75t_R FILLER_68_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_68_933 ();
 DECAPx10_ASAP7_75t_R FILLER_69_2 ();
 DECAPx10_ASAP7_75t_R FILLER_69_24 ();
 DECAPx10_ASAP7_75t_R FILLER_69_46 ();
 DECAPx10_ASAP7_75t_R FILLER_69_68 ();
 DECAPx2_ASAP7_75t_R FILLER_69_90 ();
 FILLER_ASAP7_75t_R FILLER_69_96 ();
 FILLER_ASAP7_75t_R FILLER_69_104 ();
 FILLER_ASAP7_75t_R FILLER_69_112 ();
 DECAPx6_ASAP7_75t_R FILLER_69_122 ();
 DECAPx2_ASAP7_75t_R FILLER_69_136 ();
 DECAPx2_ASAP7_75t_R FILLER_69_148 ();
 DECAPx2_ASAP7_75t_R FILLER_69_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_176 ();
 DECAPx2_ASAP7_75t_R FILLER_69_183 ();
 DECAPx4_ASAP7_75t_R FILLER_69_192 ();
 DECAPx6_ASAP7_75t_R FILLER_69_228 ();
 DECAPx1_ASAP7_75t_R FILLER_69_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_246 ();
 FILLER_ASAP7_75t_R FILLER_69_256 ();
 DECAPx2_ASAP7_75t_R FILLER_69_284 ();
 FILLER_ASAP7_75t_R FILLER_69_290 ();
 DECAPx2_ASAP7_75t_R FILLER_69_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_320 ();
 DECAPx1_ASAP7_75t_R FILLER_69_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_333 ();
 DECAPx2_ASAP7_75t_R FILLER_69_385 ();
 DECAPx10_ASAP7_75t_R FILLER_69_407 ();
 DECAPx1_ASAP7_75t_R FILLER_69_429 ();
 DECAPx4_ASAP7_75t_R FILLER_69_441 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_457 ();
 DECAPx2_ASAP7_75t_R FILLER_69_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_504 ();
 FILLER_ASAP7_75t_R FILLER_69_516 ();
 DECAPx10_ASAP7_75t_R FILLER_69_532 ();
 DECAPx6_ASAP7_75t_R FILLER_69_554 ();
 FILLER_ASAP7_75t_R FILLER_69_568 ();
 DECAPx1_ASAP7_75t_R FILLER_69_590 ();
 DECAPx1_ASAP7_75t_R FILLER_69_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_667 ();
 DECAPx2_ASAP7_75t_R FILLER_69_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_730 ();
 DECAPx10_ASAP7_75t_R FILLER_69_757 ();
 DECAPx2_ASAP7_75t_R FILLER_69_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_837 ();
 FILLER_ASAP7_75t_R FILLER_69_880 ();
 DECAPx2_ASAP7_75t_R FILLER_69_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_69_891 ();
 DECAPx6_ASAP7_75t_R FILLER_69_907 ();
 DECAPx1_ASAP7_75t_R FILLER_69_921 ();
 DECAPx2_ASAP7_75t_R FILLER_69_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_69_933 ();
 DECAPx10_ASAP7_75t_R FILLER_70_2 ();
 DECAPx10_ASAP7_75t_R FILLER_70_24 ();
 DECAPx10_ASAP7_75t_R FILLER_70_46 ();
 DECAPx10_ASAP7_75t_R FILLER_70_68 ();
 FILLER_ASAP7_75t_R FILLER_70_127 ();
 DECAPx2_ASAP7_75t_R FILLER_70_135 ();
 DECAPx2_ASAP7_75t_R FILLER_70_155 ();
 DECAPx10_ASAP7_75t_R FILLER_70_173 ();
 DECAPx4_ASAP7_75t_R FILLER_70_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_205 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_214 ();
 DECAPx2_ASAP7_75t_R FILLER_70_220 ();
 DECAPx6_ASAP7_75t_R FILLER_70_229 ();
 DECAPx1_ASAP7_75t_R FILLER_70_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_275 ();
 DECAPx4_ASAP7_75t_R FILLER_70_302 ();
 DECAPx6_ASAP7_75t_R FILLER_70_318 ();
 FILLER_ASAP7_75t_R FILLER_70_332 ();
 DECAPx4_ASAP7_75t_R FILLER_70_348 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_358 ();
 DECAPx1_ASAP7_75t_R FILLER_70_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_371 ();
 DECAPx2_ASAP7_75t_R FILLER_70_378 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_384 ();
 DECAPx6_ASAP7_75t_R FILLER_70_395 ();
 DECAPx1_ASAP7_75t_R FILLER_70_409 ();
 DECAPx2_ASAP7_75t_R FILLER_70_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_482 ();
 DECAPx10_ASAP7_75t_R FILLER_70_488 ();
 DECAPx10_ASAP7_75t_R FILLER_70_510 ();
 DECAPx10_ASAP7_75t_R FILLER_70_532 ();
 DECAPx4_ASAP7_75t_R FILLER_70_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_564 ();
 DECAPx6_ASAP7_75t_R FILLER_70_574 ();
 DECAPx2_ASAP7_75t_R FILLER_70_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_608 ();
 DECAPx4_ASAP7_75t_R FILLER_70_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_705 ();
 FILLER_ASAP7_75t_R FILLER_70_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_754 ();
 DECAPx6_ASAP7_75t_R FILLER_70_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_781 ();
 DECAPx2_ASAP7_75t_R FILLER_70_806 ();
 FILLER_ASAP7_75t_R FILLER_70_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_824 ();
 DECAPx1_ASAP7_75t_R FILLER_70_834 ();
 DECAPx6_ASAP7_75t_R FILLER_70_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_859 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_70_875 ();
 DECAPx10_ASAP7_75t_R FILLER_70_893 ();
 DECAPx6_ASAP7_75t_R FILLER_70_915 ();
 DECAPx1_ASAP7_75t_R FILLER_70_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_70_933 ();
 DECAPx10_ASAP7_75t_R FILLER_71_2 ();
 DECAPx10_ASAP7_75t_R FILLER_71_24 ();
 DECAPx10_ASAP7_75t_R FILLER_71_46 ();
 DECAPx10_ASAP7_75t_R FILLER_71_68 ();
 DECAPx4_ASAP7_75t_R FILLER_71_90 ();
 FILLER_ASAP7_75t_R FILLER_71_100 ();
 FILLER_ASAP7_75t_R FILLER_71_108 ();
 DECAPx2_ASAP7_75t_R FILLER_71_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_128 ();
 DECAPx1_ASAP7_75t_R FILLER_71_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_145 ();
 DECAPx10_ASAP7_75t_R FILLER_71_200 ();
 DECAPx2_ASAP7_75t_R FILLER_71_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_228 ();
 DECAPx4_ASAP7_75t_R FILLER_71_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_249 ();
 DECAPx4_ASAP7_75t_R FILLER_71_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_272 ();
 DECAPx2_ASAP7_75t_R FILLER_71_276 ();
 DECAPx1_ASAP7_75t_R FILLER_71_297 ();
 FILLER_ASAP7_75t_R FILLER_71_310 ();
 DECAPx1_ASAP7_75t_R FILLER_71_326 ();
 DECAPx10_ASAP7_75t_R FILLER_71_342 ();
 FILLER_ASAP7_75t_R FILLER_71_364 ();
 DECAPx1_ASAP7_75t_R FILLER_71_376 ();
 FILLER_ASAP7_75t_R FILLER_71_408 ();
 FILLER_ASAP7_75t_R FILLER_71_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_445 ();
 DECAPx1_ASAP7_75t_R FILLER_71_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_493 ();
 DECAPx10_ASAP7_75t_R FILLER_71_506 ();
 DECAPx4_ASAP7_75t_R FILLER_71_528 ();
 DECAPx2_ASAP7_75t_R FILLER_71_561 ();
 FILLER_ASAP7_75t_R FILLER_71_567 ();
 DECAPx10_ASAP7_75t_R FILLER_71_595 ();
 DECAPx6_ASAP7_75t_R FILLER_71_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_631 ();
 DECAPx10_ASAP7_75t_R FILLER_71_638 ();
 DECAPx10_ASAP7_75t_R FILLER_71_660 ();
 DECAPx10_ASAP7_75t_R FILLER_71_682 ();
 DECAPx1_ASAP7_75t_R FILLER_71_704 ();
 FILLER_ASAP7_75t_R FILLER_71_714 ();
 DECAPx4_ASAP7_75t_R FILLER_71_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_748 ();
 DECAPx1_ASAP7_75t_R FILLER_71_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_786 ();
 DECAPx6_ASAP7_75t_R FILLER_71_798 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_812 ();
 DECAPx10_ASAP7_75t_R FILLER_71_847 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_71_898 ();
 DECAPx1_ASAP7_75t_R FILLER_71_908 ();
 DECAPx4_ASAP7_75t_R FILLER_71_915 ();
 DECAPx2_ASAP7_75t_R FILLER_71_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_71_933 ();
 DECAPx10_ASAP7_75t_R FILLER_72_2 ();
 DECAPx10_ASAP7_75t_R FILLER_72_24 ();
 DECAPx10_ASAP7_75t_R FILLER_72_46 ();
 DECAPx10_ASAP7_75t_R FILLER_72_68 ();
 DECAPx10_ASAP7_75t_R FILLER_72_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_163 ();
 DECAPx2_ASAP7_75t_R FILLER_72_169 ();
 FILLER_ASAP7_75t_R FILLER_72_175 ();
 DECAPx10_ASAP7_75t_R FILLER_72_249 ();
 DECAPx6_ASAP7_75t_R FILLER_72_271 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_285 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_294 ();
 FILLER_ASAP7_75t_R FILLER_72_311 ();
 DECAPx1_ASAP7_75t_R FILLER_72_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_323 ();
 DECAPx10_ASAP7_75t_R FILLER_72_353 ();
 DECAPx10_ASAP7_75t_R FILLER_72_375 ();
 FILLER_ASAP7_75t_R FILLER_72_397 ();
 DECAPx2_ASAP7_75t_R FILLER_72_454 ();
 FILLER_ASAP7_75t_R FILLER_72_460 ();
 DECAPx1_ASAP7_75t_R FILLER_72_497 ();
 DECAPx6_ASAP7_75t_R FILLER_72_507 ();
 DECAPx2_ASAP7_75t_R FILLER_72_521 ();
 FILLER_ASAP7_75t_R FILLER_72_535 ();
 DECAPx4_ASAP7_75t_R FILLER_72_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_554 ();
 DECAPx2_ASAP7_75t_R FILLER_72_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_581 ();
 DECAPx10_ASAP7_75t_R FILLER_72_627 ();
 DECAPx2_ASAP7_75t_R FILLER_72_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_661 ();
 DECAPx10_ASAP7_75t_R FILLER_72_670 ();
 DECAPx10_ASAP7_75t_R FILLER_72_692 ();
 DECAPx10_ASAP7_75t_R FILLER_72_714 ();
 DECAPx4_ASAP7_75t_R FILLER_72_736 ();
 FILLER_ASAP7_75t_R FILLER_72_761 ();
 FILLER_ASAP7_75t_R FILLER_72_769 ();
 DECAPx6_ASAP7_75t_R FILLER_72_777 ();
 DECAPx2_ASAP7_75t_R FILLER_72_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_813 ();
 DECAPx4_ASAP7_75t_R FILLER_72_817 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_72_827 ();
 DECAPx10_ASAP7_75t_R FILLER_72_833 ();
 DECAPx10_ASAP7_75t_R FILLER_72_855 ();
 DECAPx6_ASAP7_75t_R FILLER_72_883 ();
 DECAPx4_ASAP7_75t_R FILLER_72_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_72_933 ();
 DECAPx10_ASAP7_75t_R FILLER_73_2 ();
 DECAPx10_ASAP7_75t_R FILLER_73_24 ();
 DECAPx10_ASAP7_75t_R FILLER_73_46 ();
 DECAPx10_ASAP7_75t_R FILLER_73_68 ();
 DECAPx10_ASAP7_75t_R FILLER_73_90 ();
 DECAPx4_ASAP7_75t_R FILLER_73_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_122 ();
 DECAPx1_ASAP7_75t_R FILLER_73_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_135 ();
 DECAPx4_ASAP7_75t_R FILLER_73_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_149 ();
 DECAPx2_ASAP7_75t_R FILLER_73_158 ();
 DECAPx6_ASAP7_75t_R FILLER_73_171 ();
 DECAPx1_ASAP7_75t_R FILLER_73_185 ();
 FILLER_ASAP7_75t_R FILLER_73_192 ();
 FILLER_ASAP7_75t_R FILLER_73_206 ();
 FILLER_ASAP7_75t_R FILLER_73_230 ();
 DECAPx2_ASAP7_75t_R FILLER_73_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_250 ();
 DECAPx2_ASAP7_75t_R FILLER_73_257 ();
 DECAPx2_ASAP7_75t_R FILLER_73_266 ();
 FILLER_ASAP7_75t_R FILLER_73_272 ();
 DECAPx4_ASAP7_75t_R FILLER_73_306 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_316 ();
 DECAPx4_ASAP7_75t_R FILLER_73_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_368 ();
 DECAPx2_ASAP7_75t_R FILLER_73_374 ();
 FILLER_ASAP7_75t_R FILLER_73_380 ();
 DECAPx1_ASAP7_75t_R FILLER_73_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_394 ();
 DECAPx4_ASAP7_75t_R FILLER_73_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_408 ();
 DECAPx6_ASAP7_75t_R FILLER_73_415 ();
 FILLER_ASAP7_75t_R FILLER_73_429 ();
 DECAPx1_ASAP7_75t_R FILLER_73_439 ();
 FILLER_ASAP7_75t_R FILLER_73_491 ();
 DECAPx2_ASAP7_75t_R FILLER_73_499 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_505 ();
 DECAPx1_ASAP7_75t_R FILLER_73_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_533 ();
 FILLER_ASAP7_75t_R FILLER_73_544 ();
 DECAPx6_ASAP7_75t_R FILLER_73_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_584 ();
 DECAPx10_ASAP7_75t_R FILLER_73_593 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_615 ();
 DECAPx10_ASAP7_75t_R FILLER_73_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_73_683 ();
 DECAPx2_ASAP7_75t_R FILLER_73_693 ();
 DECAPx10_ASAP7_75t_R FILLER_73_706 ();
 DECAPx10_ASAP7_75t_R FILLER_73_728 ();
 DECAPx10_ASAP7_75t_R FILLER_73_750 ();
 DECAPx10_ASAP7_75t_R FILLER_73_772 ();
 DECAPx1_ASAP7_75t_R FILLER_73_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_798 ();
 DECAPx6_ASAP7_75t_R FILLER_73_825 ();
 DECAPx2_ASAP7_75t_R FILLER_73_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_73_845 ();
 DECAPx6_ASAP7_75t_R FILLER_73_860 ();
 DECAPx4_ASAP7_75t_R FILLER_73_880 ();
 FILLER_ASAP7_75t_R FILLER_73_890 ();
 DECAPx4_ASAP7_75t_R FILLER_73_913 ();
 FILLER_ASAP7_75t_R FILLER_73_923 ();
 FILLER_ASAP7_75t_R FILLER_73_927 ();
 DECAPx10_ASAP7_75t_R FILLER_74_2 ();
 DECAPx10_ASAP7_75t_R FILLER_74_24 ();
 DECAPx10_ASAP7_75t_R FILLER_74_46 ();
 DECAPx10_ASAP7_75t_R FILLER_74_68 ();
 DECAPx6_ASAP7_75t_R FILLER_74_90 ();
 DECAPx10_ASAP7_75t_R FILLER_74_113 ();
 DECAPx10_ASAP7_75t_R FILLER_74_135 ();
 DECAPx10_ASAP7_75t_R FILLER_74_157 ();
 DECAPx6_ASAP7_75t_R FILLER_74_179 ();
 DECAPx2_ASAP7_75t_R FILLER_74_199 ();
 DECAPx10_ASAP7_75t_R FILLER_74_208 ();
 DECAPx1_ASAP7_75t_R FILLER_74_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_287 ();
 DECAPx10_ASAP7_75t_R FILLER_74_291 ();
 DECAPx1_ASAP7_75t_R FILLER_74_313 ();
 DECAPx6_ASAP7_75t_R FILLER_74_323 ();
 FILLER_ASAP7_75t_R FILLER_74_337 ();
 DECAPx2_ASAP7_75t_R FILLER_74_342 ();
 FILLER_ASAP7_75t_R FILLER_74_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_356 ();
 DECAPx6_ASAP7_75t_R FILLER_74_409 ();
 FILLER_ASAP7_75t_R FILLER_74_423 ();
 FILLER_ASAP7_75t_R FILLER_74_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_464 ();
 FILLER_ASAP7_75t_R FILLER_74_471 ();
 DECAPx1_ASAP7_75t_R FILLER_74_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_501 ();
 DECAPx1_ASAP7_75t_R FILLER_74_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_520 ();
 DECAPx10_ASAP7_75t_R FILLER_74_578 ();
 DECAPx2_ASAP7_75t_R FILLER_74_600 ();
 DECAPx1_ASAP7_75t_R FILLER_74_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_616 ();
 DECAPx1_ASAP7_75t_R FILLER_74_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_679 ();
 DECAPx1_ASAP7_75t_R FILLER_74_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_74_718 ();
 DECAPx1_ASAP7_75t_R FILLER_74_746 ();
 DECAPx4_ASAP7_75t_R FILLER_74_756 ();
 FILLER_ASAP7_75t_R FILLER_74_766 ();
 DECAPx10_ASAP7_75t_R FILLER_74_774 ();
 DECAPx6_ASAP7_75t_R FILLER_74_796 ();
 DECAPx1_ASAP7_75t_R FILLER_74_810 ();
 DECAPx6_ASAP7_75t_R FILLER_74_817 ();
 DECAPx2_ASAP7_75t_R FILLER_74_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_837 ();
 FILLER_ASAP7_75t_R FILLER_74_864 ();
 FILLER_ASAP7_75t_R FILLER_74_874 ();
 FILLERxp5_ASAP7_75t_R FILLER_74_883 ();
 DECAPx10_ASAP7_75t_R FILLER_74_892 ();
 DECAPx6_ASAP7_75t_R FILLER_74_914 ();
 DECAPx2_ASAP7_75t_R FILLER_74_928 ();
 DECAPx10_ASAP7_75t_R FILLER_75_2 ();
 DECAPx10_ASAP7_75t_R FILLER_75_24 ();
 DECAPx10_ASAP7_75t_R FILLER_75_46 ();
 DECAPx10_ASAP7_75t_R FILLER_75_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_90 ();
 FILLER_ASAP7_75t_R FILLER_75_120 ();
 DECAPx10_ASAP7_75t_R FILLER_75_128 ();
 FILLER_ASAP7_75t_R FILLER_75_150 ();
 DECAPx1_ASAP7_75t_R FILLER_75_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_163 ();
 FILLER_ASAP7_75t_R FILLER_75_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_175 ();
 DECAPx1_ASAP7_75t_R FILLER_75_183 ();
 FILLER_ASAP7_75t_R FILLER_75_199 ();
 DECAPx10_ASAP7_75t_R FILLER_75_209 ();
 DECAPx2_ASAP7_75t_R FILLER_75_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_237 ();
 FILLER_ASAP7_75t_R FILLER_75_246 ();
 DECAPx1_ASAP7_75t_R FILLER_75_254 ();
 DECAPx2_ASAP7_75t_R FILLER_75_261 ();
 FILLER_ASAP7_75t_R FILLER_75_267 ();
 DECAPx10_ASAP7_75t_R FILLER_75_279 ();
 DECAPx2_ASAP7_75t_R FILLER_75_301 ();
 FILLER_ASAP7_75t_R FILLER_75_307 ();
 DECAPx10_ASAP7_75t_R FILLER_75_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_334 ();
 DECAPx6_ASAP7_75t_R FILLER_75_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_366 ();
 DECAPx10_ASAP7_75t_R FILLER_75_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_473 ();
 DECAPx6_ASAP7_75t_R FILLER_75_482 ();
 DECAPx1_ASAP7_75t_R FILLER_75_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_500 ();
 DECAPx2_ASAP7_75t_R FILLER_75_513 ();
 DECAPx10_ASAP7_75t_R FILLER_75_526 ();
 DECAPx2_ASAP7_75t_R FILLER_75_548 ();
 FILLER_ASAP7_75t_R FILLER_75_554 ();
 DECAPx4_ASAP7_75t_R FILLER_75_588 ();
 DECAPx2_ASAP7_75t_R FILLER_75_628 ();
 DECAPx4_ASAP7_75t_R FILLER_75_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_650 ();
 DECAPx2_ASAP7_75t_R FILLER_75_654 ();
 FILLER_ASAP7_75t_R FILLER_75_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_692 ();
 DECAPx1_ASAP7_75t_R FILLER_75_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_761 ();
 DECAPx10_ASAP7_75t_R FILLER_75_798 ();
 DECAPx4_ASAP7_75t_R FILLER_75_820 ();
 FILLER_ASAP7_75t_R FILLER_75_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_75_854 ();
 DECAPx2_ASAP7_75t_R FILLER_75_858 ();
 DECAPx10_ASAP7_75t_R FILLER_75_890 ();
 DECAPx4_ASAP7_75t_R FILLER_75_912 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_75_922 ();
 FILLER_ASAP7_75t_R FILLER_75_927 ();
 DECAPx10_ASAP7_75t_R FILLER_76_2 ();
 DECAPx10_ASAP7_75t_R FILLER_76_24 ();
 DECAPx10_ASAP7_75t_R FILLER_76_46 ();
 DECAPx10_ASAP7_75t_R FILLER_76_68 ();
 DECAPx2_ASAP7_75t_R FILLER_76_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_96 ();
 FILLER_ASAP7_75t_R FILLER_76_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_179 ();
 DECAPx10_ASAP7_75t_R FILLER_76_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_219 ();
 DECAPx10_ASAP7_75t_R FILLER_76_229 ();
 DECAPx2_ASAP7_75t_R FILLER_76_251 ();
 DECAPx2_ASAP7_75t_R FILLER_76_285 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_291 ();
 DECAPx2_ASAP7_75t_R FILLER_76_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_326 ();
 DECAPx6_ASAP7_75t_R FILLER_76_353 ();
 DECAPx2_ASAP7_75t_R FILLER_76_367 ();
 DECAPx2_ASAP7_75t_R FILLER_76_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_76_385 ();
 DECAPx10_ASAP7_75t_R FILLER_76_391 ();
 DECAPx4_ASAP7_75t_R FILLER_76_413 ();
 DECAPx10_ASAP7_75t_R FILLER_76_429 ();
 DECAPx4_ASAP7_75t_R FILLER_76_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_461 ();
 DECAPx10_ASAP7_75t_R FILLER_76_467 ();
 DECAPx10_ASAP7_75t_R FILLER_76_489 ();
 DECAPx6_ASAP7_75t_R FILLER_76_511 ();
 DECAPx2_ASAP7_75t_R FILLER_76_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_531 ();
 DECAPx6_ASAP7_75t_R FILLER_76_540 ();
 DECAPx2_ASAP7_75t_R FILLER_76_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_560 ();
 DECAPx1_ASAP7_75t_R FILLER_76_574 ();
 DECAPx2_ASAP7_75t_R FILLER_76_584 ();
 FILLER_ASAP7_75t_R FILLER_76_590 ();
 DECAPx1_ASAP7_75t_R FILLER_76_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_602 ();
 DECAPx6_ASAP7_75t_R FILLER_76_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_632 ();
 FILLER_ASAP7_75t_R FILLER_76_645 ();
 FILLER_ASAP7_75t_R FILLER_76_657 ();
 DECAPx2_ASAP7_75t_R FILLER_76_671 ();
 DECAPx1_ASAP7_75t_R FILLER_76_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_712 ();
 DECAPx2_ASAP7_75t_R FILLER_76_724 ();
 FILLER_ASAP7_75t_R FILLER_76_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_746 ();
 FILLER_ASAP7_75t_R FILLER_76_802 ();
 FILLER_ASAP7_75t_R FILLER_76_815 ();
 DECAPx1_ASAP7_75t_R FILLER_76_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_76_829 ();
 DECAPx10_ASAP7_75t_R FILLER_76_846 ();
 DECAPx10_ASAP7_75t_R FILLER_76_868 ();
 DECAPx6_ASAP7_75t_R FILLER_76_890 ();
 DECAPx1_ASAP7_75t_R FILLER_76_904 ();
 DECAPx10_ASAP7_75t_R FILLER_77_2 ();
 DECAPx10_ASAP7_75t_R FILLER_77_24 ();
 DECAPx10_ASAP7_75t_R FILLER_77_46 ();
 DECAPx10_ASAP7_75t_R FILLER_77_68 ();
 DECAPx10_ASAP7_75t_R FILLER_77_90 ();
 FILLER_ASAP7_75t_R FILLER_77_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_120 ();
 DECAPx6_ASAP7_75t_R FILLER_77_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_202 ();
 DECAPx2_ASAP7_75t_R FILLER_77_240 ();
 FILLER_ASAP7_75t_R FILLER_77_246 ();
 FILLER_ASAP7_75t_R FILLER_77_258 ();
 DECAPx1_ASAP7_75t_R FILLER_77_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_269 ();
 FILLER_ASAP7_75t_R FILLER_77_296 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_310 ();
 DECAPx10_ASAP7_75t_R FILLER_77_346 ();
 DECAPx10_ASAP7_75t_R FILLER_77_368 ();
 DECAPx6_ASAP7_75t_R FILLER_77_390 ();
 FILLER_ASAP7_75t_R FILLER_77_404 ();
 DECAPx2_ASAP7_75t_R FILLER_77_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_431 ();
 DECAPx1_ASAP7_75t_R FILLER_77_435 ();
 DECAPx10_ASAP7_75t_R FILLER_77_442 ();
 DECAPx10_ASAP7_75t_R FILLER_77_464 ();
 DECAPx4_ASAP7_75t_R FILLER_77_486 ();
 FILLER_ASAP7_75t_R FILLER_77_496 ();
 DECAPx1_ASAP7_75t_R FILLER_77_504 ();
 DECAPx6_ASAP7_75t_R FILLER_77_514 ();
 DECAPx2_ASAP7_75t_R FILLER_77_528 ();
 DECAPx2_ASAP7_75t_R FILLER_77_544 ();
 FILLER_ASAP7_75t_R FILLER_77_550 ();
 DECAPx10_ASAP7_75t_R FILLER_77_560 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_582 ();
 DECAPx10_ASAP7_75t_R FILLER_77_605 ();
 DECAPx10_ASAP7_75t_R FILLER_77_633 ();
 DECAPx10_ASAP7_75t_R FILLER_77_655 ();
 DECAPx10_ASAP7_75t_R FILLER_77_677 ();
 DECAPx10_ASAP7_75t_R FILLER_77_699 ();
 DECAPx10_ASAP7_75t_R FILLER_77_721 ();
 DECAPx2_ASAP7_75t_R FILLER_77_743 ();
 FILLER_ASAP7_75t_R FILLER_77_749 ();
 DECAPx2_ASAP7_75t_R FILLER_77_767 ();
 FILLER_ASAP7_75t_R FILLER_77_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_798 ();
 DECAPx2_ASAP7_75t_R FILLER_77_847 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_859 ();
 DECAPx4_ASAP7_75t_R FILLER_77_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_878 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_77_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_77_905 ();
 FILLER_ASAP7_75t_R FILLER_77_909 ();
 DECAPx1_ASAP7_75t_R FILLER_77_918 ();
 FILLER_ASAP7_75t_R FILLER_77_927 ();
 DECAPx10_ASAP7_75t_R FILLER_78_2 ();
 DECAPx10_ASAP7_75t_R FILLER_78_24 ();
 DECAPx10_ASAP7_75t_R FILLER_78_46 ();
 DECAPx10_ASAP7_75t_R FILLER_78_68 ();
 DECAPx10_ASAP7_75t_R FILLER_78_90 ();
 DECAPx10_ASAP7_75t_R FILLER_78_112 ();
 DECAPx2_ASAP7_75t_R FILLER_78_134 ();
 FILLER_ASAP7_75t_R FILLER_78_140 ();
 DECAPx6_ASAP7_75t_R FILLER_78_148 ();
 DECAPx1_ASAP7_75t_R FILLER_78_162 ();
 DECAPx1_ASAP7_75t_R FILLER_78_172 ();
 FILLER_ASAP7_75t_R FILLER_78_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_215 ();
 DECAPx1_ASAP7_75t_R FILLER_78_222 ();
 DECAPx6_ASAP7_75t_R FILLER_78_242 ();
 DECAPx2_ASAP7_75t_R FILLER_78_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_262 ();
 DECAPx2_ASAP7_75t_R FILLER_78_269 ();
 FILLER_ASAP7_75t_R FILLER_78_275 ();
 DECAPx6_ASAP7_75t_R FILLER_78_292 ();
 FILLER_ASAP7_75t_R FILLER_78_306 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_322 ();
 DECAPx2_ASAP7_75t_R FILLER_78_351 ();
 DECAPx1_ASAP7_75t_R FILLER_78_383 ();
 DECAPx1_ASAP7_75t_R FILLER_78_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_402 ();
 DECAPx4_ASAP7_75t_R FILLER_78_452 ();
 FILLER_ASAP7_75t_R FILLER_78_470 ();
 DECAPx2_ASAP7_75t_R FILLER_78_475 ();
 FILLER_ASAP7_75t_R FILLER_78_481 ();
 FILLER_ASAP7_75t_R FILLER_78_489 ();
 DECAPx2_ASAP7_75t_R FILLER_78_509 ();
 FILLER_ASAP7_75t_R FILLER_78_515 ();
 DECAPx2_ASAP7_75t_R FILLER_78_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_533 ();
 FILLER_ASAP7_75t_R FILLER_78_541 ();
 DECAPx6_ASAP7_75t_R FILLER_78_571 ();
 DECAPx1_ASAP7_75t_R FILLER_78_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_589 ();
 DECAPx10_ASAP7_75t_R FILLER_78_608 ();
 DECAPx4_ASAP7_75t_R FILLER_78_630 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_649 ();
 DECAPx6_ASAP7_75t_R FILLER_78_659 ();
 DECAPx4_ASAP7_75t_R FILLER_78_683 ();
 DECAPx10_ASAP7_75t_R FILLER_78_705 ();
 DECAPx10_ASAP7_75t_R FILLER_78_727 ();
 DECAPx10_ASAP7_75t_R FILLER_78_749 ();
 DECAPx10_ASAP7_75t_R FILLER_78_771 ();
 DECAPx2_ASAP7_75t_R FILLER_78_793 ();
 FILLER_ASAP7_75t_R FILLER_78_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_807 ();
 DECAPx4_ASAP7_75t_R FILLER_78_839 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_860 ();
 FILLER_ASAP7_75t_R FILLER_78_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_78_923 ();
 DECAPx1_ASAP7_75t_R FILLER_78_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_78_933 ();
 DECAPx10_ASAP7_75t_R FILLER_79_2 ();
 DECAPx10_ASAP7_75t_R FILLER_79_24 ();
 DECAPx10_ASAP7_75t_R FILLER_79_46 ();
 DECAPx6_ASAP7_75t_R FILLER_79_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_100 ();
 DECAPx2_ASAP7_75t_R FILLER_79_104 ();
 FILLER_ASAP7_75t_R FILLER_79_110 ();
 DECAPx4_ASAP7_75t_R FILLER_79_118 ();
 FILLER_ASAP7_75t_R FILLER_79_134 ();
 DECAPx2_ASAP7_75t_R FILLER_79_142 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_148 ();
 DECAPx6_ASAP7_75t_R FILLER_79_164 ();
 DECAPx1_ASAP7_75t_R FILLER_79_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_182 ();
 DECAPx6_ASAP7_75t_R FILLER_79_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_203 ();
 DECAPx2_ASAP7_75t_R FILLER_79_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_223 ();
 DECAPx1_ASAP7_75t_R FILLER_79_232 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_248 ();
 FILLER_ASAP7_75t_R FILLER_79_277 ();
 DECAPx6_ASAP7_75t_R FILLER_79_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_299 ();
 FILLER_ASAP7_75t_R FILLER_79_329 ();
 FILLER_ASAP7_75t_R FILLER_79_337 ();
 FILLER_ASAP7_75t_R FILLER_79_342 ();
 DECAPx2_ASAP7_75t_R FILLER_79_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_400 ();
 DECAPx1_ASAP7_75t_R FILLER_79_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_431 ();
 DECAPx2_ASAP7_75t_R FILLER_79_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_484 ();
 DECAPx1_ASAP7_75t_R FILLER_79_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_509 ();
 DECAPx2_ASAP7_75t_R FILLER_79_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_534 ();
 DECAPx10_ASAP7_75t_R FILLER_79_541 ();
 DECAPx2_ASAP7_75t_R FILLER_79_563 ();
 FILLER_ASAP7_75t_R FILLER_79_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_584 ();
 DECAPx10_ASAP7_75t_R FILLER_79_593 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_615 ();
 DECAPx4_ASAP7_75t_R FILLER_79_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_665 ();
 DECAPx2_ASAP7_75t_R FILLER_79_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_684 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_695 ();
 DECAPx4_ASAP7_75t_R FILLER_79_732 ();
 DECAPx1_ASAP7_75t_R FILLER_79_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_757 ();
 DECAPx6_ASAP7_75t_R FILLER_79_766 ();
 DECAPx6_ASAP7_75t_R FILLER_79_794 ();
 DECAPx2_ASAP7_75t_R FILLER_79_808 ();
 FILLER_ASAP7_75t_R FILLER_79_820 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_79_825 ();
 DECAPx6_ASAP7_75t_R FILLER_79_831 ();
 DECAPx2_ASAP7_75t_R FILLER_79_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_887 ();
 FILLER_ASAP7_75t_R FILLER_79_894 ();
 FILLER_ASAP7_75t_R FILLER_79_899 ();
 DECAPx6_ASAP7_75t_R FILLER_79_907 ();
 DECAPx1_ASAP7_75t_R FILLER_79_921 ();
 DECAPx2_ASAP7_75t_R FILLER_79_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_79_933 ();
 DECAPx10_ASAP7_75t_R FILLER_80_2 ();
 DECAPx10_ASAP7_75t_R FILLER_80_24 ();
 DECAPx10_ASAP7_75t_R FILLER_80_46 ();
 DECAPx4_ASAP7_75t_R FILLER_80_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_113 ();
 FILLER_ASAP7_75t_R FILLER_80_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_172 ();
 DECAPx2_ASAP7_75t_R FILLER_80_179 ();
 FILLER_ASAP7_75t_R FILLER_80_185 ();
 DECAPx10_ASAP7_75t_R FILLER_80_201 ();
 DECAPx6_ASAP7_75t_R FILLER_80_223 ();
 DECAPx2_ASAP7_75t_R FILLER_80_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_265 ();
 DECAPx1_ASAP7_75t_R FILLER_80_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_314 ();
 DECAPx2_ASAP7_75t_R FILLER_80_318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_324 ();
 DECAPx4_ASAP7_75t_R FILLER_80_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_357 ();
 FILLER_ASAP7_75t_R FILLER_80_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_382 ();
 DECAPx2_ASAP7_75t_R FILLER_80_395 ();
 DECAPx2_ASAP7_75t_R FILLER_80_407 ();
 FILLER_ASAP7_75t_R FILLER_80_413 ();
 DECAPx4_ASAP7_75t_R FILLER_80_418 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_428 ();
 DECAPx1_ASAP7_75t_R FILLER_80_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_453 ();
 DECAPx10_ASAP7_75t_R FILLER_80_490 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_512 ();
 FILLER_ASAP7_75t_R FILLER_80_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_531 ();
 DECAPx10_ASAP7_75t_R FILLER_80_541 ();
 DECAPx2_ASAP7_75t_R FILLER_80_563 ();
 FILLER_ASAP7_75t_R FILLER_80_569 ();
 DECAPx1_ASAP7_75t_R FILLER_80_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_601 ();
 DECAPx1_ASAP7_75t_R FILLER_80_614 ();
 DECAPx6_ASAP7_75t_R FILLER_80_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_676 ();
 DECAPx2_ASAP7_75t_R FILLER_80_684 ();
 FILLER_ASAP7_75t_R FILLER_80_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_704 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_80_762 ();
 DECAPx10_ASAP7_75t_R FILLER_80_805 ();
 DECAPx10_ASAP7_75t_R FILLER_80_827 ();
 DECAPx10_ASAP7_75t_R FILLER_80_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_80_871 ();
 DECAPx10_ASAP7_75t_R FILLER_80_878 ();
 DECAPx10_ASAP7_75t_R FILLER_80_900 ();
 DECAPx4_ASAP7_75t_R FILLER_80_922 ();
 FILLER_ASAP7_75t_R FILLER_80_932 ();
 DECAPx10_ASAP7_75t_R FILLER_81_2 ();
 DECAPx10_ASAP7_75t_R FILLER_81_24 ();
 DECAPx10_ASAP7_75t_R FILLER_81_46 ();
 DECAPx10_ASAP7_75t_R FILLER_81_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_90 ();
 DECAPx6_ASAP7_75t_R FILLER_81_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_157 ();
 DECAPx10_ASAP7_75t_R FILLER_81_187 ();
 DECAPx4_ASAP7_75t_R FILLER_81_209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_219 ();
 DECAPx10_ASAP7_75t_R FILLER_81_231 ();
 DECAPx10_ASAP7_75t_R FILLER_81_253 ();
 DECAPx2_ASAP7_75t_R FILLER_81_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_287 ();
 DECAPx10_ASAP7_75t_R FILLER_81_297 ();
 DECAPx4_ASAP7_75t_R FILLER_81_319 ();
 FILLER_ASAP7_75t_R FILLER_81_329 ();
 DECAPx2_ASAP7_75t_R FILLER_81_363 ();
 FILLER_ASAP7_75t_R FILLER_81_369 ();
 DECAPx6_ASAP7_75t_R FILLER_81_374 ();
 FILLER_ASAP7_75t_R FILLER_81_388 ();
 DECAPx6_ASAP7_75t_R FILLER_81_395 ();
 DECAPx1_ASAP7_75t_R FILLER_81_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_413 ();
 DECAPx6_ASAP7_75t_R FILLER_81_422 ();
 DECAPx1_ASAP7_75t_R FILLER_81_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_440 ();
 FILLER_ASAP7_75t_R FILLER_81_469 ();
 DECAPx10_ASAP7_75t_R FILLER_81_488 ();
 DECAPx10_ASAP7_75t_R FILLER_81_510 ();
 DECAPx2_ASAP7_75t_R FILLER_81_532 ();
 FILLER_ASAP7_75t_R FILLER_81_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_570 ();
 DECAPx6_ASAP7_75t_R FILLER_81_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_607 ();
 DECAPx6_ASAP7_75t_R FILLER_81_648 ();
 DECAPx1_ASAP7_75t_R FILLER_81_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_666 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_707 ();
 DECAPx2_ASAP7_75t_R FILLER_81_716 ();
 FILLER_ASAP7_75t_R FILLER_81_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_727 ();
 DECAPx2_ASAP7_75t_R FILLER_81_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_737 ();
 DECAPx1_ASAP7_75t_R FILLER_81_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_748 ();
 DECAPx1_ASAP7_75t_R FILLER_81_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_756 ();
 DECAPx2_ASAP7_75t_R FILLER_81_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_789 ();
 DECAPx2_ASAP7_75t_R FILLER_81_793 ();
 FILLER_ASAP7_75t_R FILLER_81_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_804 ();
 DECAPx6_ASAP7_75t_R FILLER_81_817 ();
 FILLER_ASAP7_75t_R FILLER_81_831 ();
 DECAPx1_ASAP7_75t_R FILLER_81_840 ();
 DECAPx10_ASAP7_75t_R FILLER_81_851 ();
 DECAPx10_ASAP7_75t_R FILLER_81_873 ();
 DECAPx2_ASAP7_75t_R FILLER_81_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_81_901 ();
 DECAPx1_ASAP7_75t_R FILLER_81_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_924 ();
 DECAPx2_ASAP7_75t_R FILLER_81_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_81_933 ();
 DECAPx10_ASAP7_75t_R FILLER_82_2 ();
 DECAPx10_ASAP7_75t_R FILLER_82_24 ();
 DECAPx10_ASAP7_75t_R FILLER_82_46 ();
 DECAPx4_ASAP7_75t_R FILLER_82_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_78 ();
 DECAPx1_ASAP7_75t_R FILLER_82_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_111 ();
 FILLER_ASAP7_75t_R FILLER_82_118 ();
 DECAPx6_ASAP7_75t_R FILLER_82_129 ();
 DECAPx2_ASAP7_75t_R FILLER_82_143 ();
 DECAPx4_ASAP7_75t_R FILLER_82_155 ();
 FILLER_ASAP7_75t_R FILLER_82_165 ();
 FILLER_ASAP7_75t_R FILLER_82_173 ();
 DECAPx6_ASAP7_75t_R FILLER_82_192 ();
 DECAPx2_ASAP7_75t_R FILLER_82_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_212 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_239 ();
 DECAPx6_ASAP7_75t_R FILLER_82_268 ();
 DECAPx1_ASAP7_75t_R FILLER_82_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_286 ();
 DECAPx6_ASAP7_75t_R FILLER_82_301 ();
 FILLER_ASAP7_75t_R FILLER_82_315 ();
 DECAPx2_ASAP7_75t_R FILLER_82_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_329 ();
 DECAPx2_ASAP7_75t_R FILLER_82_340 ();
 DECAPx6_ASAP7_75t_R FILLER_82_354 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_368 ();
 DECAPx6_ASAP7_75t_R FILLER_82_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_395 ();
 DECAPx2_ASAP7_75t_R FILLER_82_404 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_422 ();
 DECAPx2_ASAP7_75t_R FILLER_82_439 ();
 DECAPx2_ASAP7_75t_R FILLER_82_456 ();
 DECAPx2_ASAP7_75t_R FILLER_82_464 ();
 FILLER_ASAP7_75t_R FILLER_82_470 ();
 DECAPx4_ASAP7_75t_R FILLER_82_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_488 ();
 DECAPx1_ASAP7_75t_R FILLER_82_495 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_499 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_513 ();
 DECAPx6_ASAP7_75t_R FILLER_82_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_548 ();
 DECAPx2_ASAP7_75t_R FILLER_82_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_608 ();
 DECAPx1_ASAP7_75t_R FILLER_82_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_625 ();
 DECAPx10_ASAP7_75t_R FILLER_82_652 ();
 DECAPx1_ASAP7_75t_R FILLER_82_674 ();
 DECAPx2_ASAP7_75t_R FILLER_82_684 ();
 DECAPx6_ASAP7_75t_R FILLER_82_696 ();
 DECAPx1_ASAP7_75t_R FILLER_82_715 ();
 DECAPx10_ASAP7_75t_R FILLER_82_726 ();
 DECAPx4_ASAP7_75t_R FILLER_82_748 ();
 FILLER_ASAP7_75t_R FILLER_82_758 ();
 DECAPx2_ASAP7_75t_R FILLER_82_766 ();
 DECAPx6_ASAP7_75t_R FILLER_82_775 ();
 DECAPx2_ASAP7_75t_R FILLER_82_789 ();
 DECAPx1_ASAP7_75t_R FILLER_82_830 ();
 DECAPx2_ASAP7_75t_R FILLER_82_866 ();
 FILLER_ASAP7_75t_R FILLER_82_878 ();
 DECAPx2_ASAP7_75t_R FILLER_82_894 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_82_900 ();
 DECAPx1_ASAP7_75t_R FILLER_82_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_82_933 ();
 DECAPx10_ASAP7_75t_R FILLER_83_2 ();
 DECAPx10_ASAP7_75t_R FILLER_83_24 ();
 DECAPx10_ASAP7_75t_R FILLER_83_46 ();
 DECAPx6_ASAP7_75t_R FILLER_83_68 ();
 DECAPx1_ASAP7_75t_R FILLER_83_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_86 ();
 DECAPx10_ASAP7_75t_R FILLER_83_102 ();
 DECAPx6_ASAP7_75t_R FILLER_83_124 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_138 ();
 DECAPx6_ASAP7_75t_R FILLER_83_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_181 ();
 DECAPx2_ASAP7_75t_R FILLER_83_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_206 ();
 DECAPx1_ASAP7_75t_R FILLER_83_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_234 ();
 DECAPx2_ASAP7_75t_R FILLER_83_243 ();
 FILLER_ASAP7_75t_R FILLER_83_261 ();
 DECAPx2_ASAP7_75t_R FILLER_83_283 ();
 FILLER_ASAP7_75t_R FILLER_83_289 ();
 DECAPx2_ASAP7_75t_R FILLER_83_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_304 ();
 DECAPx6_ASAP7_75t_R FILLER_83_335 ();
 FILLER_ASAP7_75t_R FILLER_83_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_360 ();
 FILLER_ASAP7_75t_R FILLER_83_393 ();
 DECAPx10_ASAP7_75t_R FILLER_83_445 ();
 DECAPx6_ASAP7_75t_R FILLER_83_467 ();
 DECAPx1_ASAP7_75t_R FILLER_83_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_485 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_499 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_512 ();
 DECAPx10_ASAP7_75t_R FILLER_83_523 ();
 DECAPx10_ASAP7_75t_R FILLER_83_565 ();
 DECAPx10_ASAP7_75t_R FILLER_83_587 ();
 DECAPx10_ASAP7_75t_R FILLER_83_609 ();
 FILLER_ASAP7_75t_R FILLER_83_631 ();
 DECAPx10_ASAP7_75t_R FILLER_83_659 ();
 DECAPx6_ASAP7_75t_R FILLER_83_681 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_695 ();
 DECAPx2_ASAP7_75t_R FILLER_83_731 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_737 ();
 DECAPx10_ASAP7_75t_R FILLER_83_766 ();
 DECAPx2_ASAP7_75t_R FILLER_83_788 ();
 DECAPx1_ASAP7_75t_R FILLER_83_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_804 ();
 DECAPx6_ASAP7_75t_R FILLER_83_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_83_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_83_841 ();
 FILLER_ASAP7_75t_R FILLER_83_864 ();
 DECAPx6_ASAP7_75t_R FILLER_83_905 ();
 DECAPx2_ASAP7_75t_R FILLER_83_919 ();
 FILLER_ASAP7_75t_R FILLER_83_927 ();
 DECAPx10_ASAP7_75t_R FILLER_84_2 ();
 DECAPx10_ASAP7_75t_R FILLER_84_24 ();
 DECAPx10_ASAP7_75t_R FILLER_84_46 ();
 DECAPx10_ASAP7_75t_R FILLER_84_68 ();
 DECAPx10_ASAP7_75t_R FILLER_84_90 ();
 DECAPx2_ASAP7_75t_R FILLER_84_112 ();
 FILLER_ASAP7_75t_R FILLER_84_118 ();
 DECAPx6_ASAP7_75t_R FILLER_84_126 ();
 DECAPx1_ASAP7_75t_R FILLER_84_140 ();
 DECAPx2_ASAP7_75t_R FILLER_84_150 ();
 DECAPx6_ASAP7_75t_R FILLER_84_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_197 ();
 DECAPx2_ASAP7_75t_R FILLER_84_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_256 ();
 DECAPx1_ASAP7_75t_R FILLER_84_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_267 ();
 DECAPx6_ASAP7_75t_R FILLER_84_290 ();
 FILLER_ASAP7_75t_R FILLER_84_304 ();
 DECAPx6_ASAP7_75t_R FILLER_84_318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_332 ();
 DECAPx1_ASAP7_75t_R FILLER_84_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_351 ();
 FILLER_ASAP7_75t_R FILLER_84_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_419 ();
 FILLER_ASAP7_75t_R FILLER_84_460 ();
 DECAPx4_ASAP7_75t_R FILLER_84_470 ();
 DECAPx2_ASAP7_75t_R FILLER_84_494 ();
 FILLER_ASAP7_75t_R FILLER_84_500 ();
 DECAPx6_ASAP7_75t_R FILLER_84_508 ();
 DECAPx2_ASAP7_75t_R FILLER_84_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_528 ();
 DECAPx2_ASAP7_75t_R FILLER_84_536 ();
 FILLER_ASAP7_75t_R FILLER_84_542 ();
 DECAPx10_ASAP7_75t_R FILLER_84_551 ();
 DECAPx1_ASAP7_75t_R FILLER_84_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_577 ();
 DECAPx2_ASAP7_75t_R FILLER_84_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_600 ();
 DECAPx10_ASAP7_75t_R FILLER_84_610 ();
 DECAPx2_ASAP7_75t_R FILLER_84_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_645 ();
 DECAPx1_ASAP7_75t_R FILLER_84_661 ();
 FILLER_ASAP7_75t_R FILLER_84_675 ();
 DECAPx1_ASAP7_75t_R FILLER_84_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_688 ();
 DECAPx6_ASAP7_75t_R FILLER_84_695 ();
 FILLER_ASAP7_75t_R FILLER_84_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_718 ();
 FILLER_ASAP7_75t_R FILLER_84_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_84_746 ();
 DECAPx6_ASAP7_75t_R FILLER_84_765 ();
 DECAPx2_ASAP7_75t_R FILLER_84_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_785 ();
 DECAPx10_ASAP7_75t_R FILLER_84_789 ();
 DECAPx2_ASAP7_75t_R FILLER_84_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_817 ();
 DECAPx10_ASAP7_75t_R FILLER_84_825 ();
 DECAPx4_ASAP7_75t_R FILLER_84_847 ();
 FILLER_ASAP7_75t_R FILLER_84_857 ();
 DECAPx4_ASAP7_75t_R FILLER_84_866 ();
 FILLER_ASAP7_75t_R FILLER_84_876 ();
 DECAPx10_ASAP7_75t_R FILLER_84_907 ();
 DECAPx1_ASAP7_75t_R FILLER_84_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_84_933 ();
 DECAPx10_ASAP7_75t_R FILLER_85_2 ();
 DECAPx10_ASAP7_75t_R FILLER_85_24 ();
 DECAPx10_ASAP7_75t_R FILLER_85_46 ();
 DECAPx10_ASAP7_75t_R FILLER_85_68 ();
 DECAPx10_ASAP7_75t_R FILLER_85_90 ();
 DECAPx6_ASAP7_75t_R FILLER_85_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_155 ();
 DECAPx2_ASAP7_75t_R FILLER_85_159 ();
 DECAPx4_ASAP7_75t_R FILLER_85_191 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_201 ();
 DECAPx6_ASAP7_75t_R FILLER_85_219 ();
 DECAPx1_ASAP7_75t_R FILLER_85_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_237 ();
 DECAPx10_ASAP7_75t_R FILLER_85_241 ();
 DECAPx1_ASAP7_75t_R FILLER_85_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_267 ();
 DECAPx2_ASAP7_75t_R FILLER_85_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_282 ();
 DECAPx2_ASAP7_75t_R FILLER_85_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_297 ();
 DECAPx6_ASAP7_75t_R FILLER_85_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_462 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_487 ();
 DECAPx10_ASAP7_75t_R FILLER_85_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_516 ();
 DECAPx1_ASAP7_75t_R FILLER_85_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_529 ();
 DECAPx10_ASAP7_75t_R FILLER_85_550 ();
 DECAPx1_ASAP7_75t_R FILLER_85_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_613 ();
 DECAPx10_ASAP7_75t_R FILLER_85_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_646 ();
 DECAPx1_ASAP7_75t_R FILLER_85_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_698 ();
 FILLER_ASAP7_75t_R FILLER_85_731 ();
 FILLER_ASAP7_75t_R FILLER_85_738 ();
 DECAPx6_ASAP7_75t_R FILLER_85_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_85_779 ();
 FILLER_ASAP7_75t_R FILLER_85_797 ();
 DECAPx6_ASAP7_75t_R FILLER_85_803 ();
 FILLER_ASAP7_75t_R FILLER_85_817 ();
 DECAPx10_ASAP7_75t_R FILLER_85_839 ();
 FILLER_ASAP7_75t_R FILLER_85_861 ();
 DECAPx6_ASAP7_75t_R FILLER_85_876 ();
 FILLER_ASAP7_75t_R FILLER_85_890 ();
 DECAPx10_ASAP7_75t_R FILLER_85_898 ();
 DECAPx1_ASAP7_75t_R FILLER_85_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_924 ();
 DECAPx2_ASAP7_75t_R FILLER_85_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_85_933 ();
 DECAPx10_ASAP7_75t_R FILLER_86_2 ();
 DECAPx10_ASAP7_75t_R FILLER_86_24 ();
 DECAPx10_ASAP7_75t_R FILLER_86_46 ();
 DECAPx10_ASAP7_75t_R FILLER_86_68 ();
 DECAPx1_ASAP7_75t_R FILLER_86_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_94 ();
 DECAPx6_ASAP7_75t_R FILLER_86_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_115 ();
 DECAPx1_ASAP7_75t_R FILLER_86_122 ();
 DECAPx10_ASAP7_75t_R FILLER_86_129 ();
 DECAPx2_ASAP7_75t_R FILLER_86_151 ();
 DECAPx2_ASAP7_75t_R FILLER_86_163 ();
 DECAPx1_ASAP7_75t_R FILLER_86_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_179 ();
 DECAPx10_ASAP7_75t_R FILLER_86_183 ();
 DECAPx10_ASAP7_75t_R FILLER_86_205 ();
 DECAPx6_ASAP7_75t_R FILLER_86_227 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_241 ();
 DECAPx1_ASAP7_75t_R FILLER_86_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_254 ();
 DECAPx2_ASAP7_75t_R FILLER_86_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_274 ();
 FILLER_ASAP7_75t_R FILLER_86_301 ();
 DECAPx10_ASAP7_75t_R FILLER_86_312 ();
 DECAPx4_ASAP7_75t_R FILLER_86_334 ();
 FILLER_ASAP7_75t_R FILLER_86_344 ();
 DECAPx4_ASAP7_75t_R FILLER_86_349 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_359 ();
 DECAPx1_ASAP7_75t_R FILLER_86_374 ();
 FILLER_ASAP7_75t_R FILLER_86_409 ();
 FILLER_ASAP7_75t_R FILLER_86_423 ();
 DECAPx2_ASAP7_75t_R FILLER_86_464 ();
 DECAPx2_ASAP7_75t_R FILLER_86_476 ();
 DECAPx10_ASAP7_75t_R FILLER_86_485 ();
 FILLER_ASAP7_75t_R FILLER_86_514 ();
 DECAPx2_ASAP7_75t_R FILLER_86_536 ();
 FILLER_ASAP7_75t_R FILLER_86_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_588 ();
 DECAPx1_ASAP7_75t_R FILLER_86_612 ();
 DECAPx10_ASAP7_75t_R FILLER_86_631 ();
 DECAPx2_ASAP7_75t_R FILLER_86_653 ();
 FILLER_ASAP7_75t_R FILLER_86_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_682 ();
 FILLER_ASAP7_75t_R FILLER_86_712 ();
 DECAPx6_ASAP7_75t_R FILLER_86_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_779 ();
 DECAPx4_ASAP7_75t_R FILLER_86_800 ();
 DECAPx4_ASAP7_75t_R FILLER_86_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_86_826 ();
 DECAPx2_ASAP7_75t_R FILLER_86_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_86_842 ();
 DECAPx10_ASAP7_75t_R FILLER_86_856 ();
 DECAPx10_ASAP7_75t_R FILLER_86_878 ();
 DECAPx2_ASAP7_75t_R FILLER_86_900 ();
 FILLER_ASAP7_75t_R FILLER_86_906 ();
 DECAPx10_ASAP7_75t_R FILLER_87_2 ();
 DECAPx10_ASAP7_75t_R FILLER_87_24 ();
 DECAPx10_ASAP7_75t_R FILLER_87_46 ();
 DECAPx6_ASAP7_75t_R FILLER_87_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_82 ();
 DECAPx10_ASAP7_75t_R FILLER_87_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_139 ();
 DECAPx4_ASAP7_75t_R FILLER_87_143 ();
 FILLER_ASAP7_75t_R FILLER_87_153 ();
 DECAPx2_ASAP7_75t_R FILLER_87_169 ();
 DECAPx2_ASAP7_75t_R FILLER_87_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_187 ();
 DECAPx10_ASAP7_75t_R FILLER_87_191 ();
 DECAPx1_ASAP7_75t_R FILLER_87_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_217 ();
 DECAPx2_ASAP7_75t_R FILLER_87_227 ();
 DECAPx1_ASAP7_75t_R FILLER_87_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_287 ();
 DECAPx2_ASAP7_75t_R FILLER_87_293 ();
 DECAPx6_ASAP7_75t_R FILLER_87_305 ();
 FILLER_ASAP7_75t_R FILLER_87_319 ();
 DECAPx6_ASAP7_75t_R FILLER_87_329 ();
 DECAPx2_ASAP7_75t_R FILLER_87_343 ();
 DECAPx10_ASAP7_75t_R FILLER_87_355 ();
 DECAPx1_ASAP7_75t_R FILLER_87_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_381 ();
 DECAPx10_ASAP7_75t_R FILLER_87_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_445 ();
 DECAPx4_ASAP7_75t_R FILLER_87_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_487 ();
 DECAPx2_ASAP7_75t_R FILLER_87_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_506 ();
 DECAPx6_ASAP7_75t_R FILLER_87_527 ();
 FILLER_ASAP7_75t_R FILLER_87_541 ();
 DECAPx6_ASAP7_75t_R FILLER_87_550 ();
 DECAPx1_ASAP7_75t_R FILLER_87_564 ();
 DECAPx4_ASAP7_75t_R FILLER_87_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_590 ();
 DECAPx2_ASAP7_75t_R FILLER_87_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_603 ();
 DECAPx4_ASAP7_75t_R FILLER_87_610 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_620 ();
 FILLER_ASAP7_75t_R FILLER_87_629 ();
 DECAPx10_ASAP7_75t_R FILLER_87_647 ();
 DECAPx6_ASAP7_75t_R FILLER_87_669 ();
 DECAPx1_ASAP7_75t_R FILLER_87_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_693 ();
 DECAPx2_ASAP7_75t_R FILLER_87_708 ();
 DECAPx1_ASAP7_75t_R FILLER_87_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_721 ();
 FILLER_ASAP7_75t_R FILLER_87_754 ();
 DECAPx2_ASAP7_75t_R FILLER_87_762 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_768 ();
 DECAPx4_ASAP7_75t_R FILLER_87_777 ();
 DECAPx1_ASAP7_75t_R FILLER_87_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_811 ();
 DECAPx1_ASAP7_75t_R FILLER_87_817 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_87_827 ();
 FILLER_ASAP7_75t_R FILLER_87_850 ();
 DECAPx2_ASAP7_75t_R FILLER_87_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_865 ();
 DECAPx10_ASAP7_75t_R FILLER_87_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_898 ();
 DECAPx2_ASAP7_75t_R FILLER_87_905 ();
 DECAPx2_ASAP7_75t_R FILLER_87_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_87_924 ();
 DECAPx1_ASAP7_75t_R FILLER_87_930 ();
 DECAPx10_ASAP7_75t_R FILLER_88_2 ();
 DECAPx10_ASAP7_75t_R FILLER_88_24 ();
 DECAPx10_ASAP7_75t_R FILLER_88_46 ();
 DECAPx10_ASAP7_75t_R FILLER_88_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_192 ();
 DECAPx2_ASAP7_75t_R FILLER_88_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_205 ();
 DECAPx10_ASAP7_75t_R FILLER_88_270 ();
 DECAPx6_ASAP7_75t_R FILLER_88_292 ();
 DECAPx1_ASAP7_75t_R FILLER_88_306 ();
 DECAPx6_ASAP7_75t_R FILLER_88_364 ();
 DECAPx10_ASAP7_75t_R FILLER_88_386 ();
 DECAPx10_ASAP7_75t_R FILLER_88_418 ();
 DECAPx4_ASAP7_75t_R FILLER_88_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_450 ();
 DECAPx1_ASAP7_75t_R FILLER_88_464 ();
 DECAPx2_ASAP7_75t_R FILLER_88_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_477 ();
 DECAPx6_ASAP7_75t_R FILLER_88_504 ();
 DECAPx1_ASAP7_75t_R FILLER_88_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_522 ();
 DECAPx10_ASAP7_75t_R FILLER_88_529 ();
 DECAPx4_ASAP7_75t_R FILLER_88_551 ();
 FILLER_ASAP7_75t_R FILLER_88_561 ();
 DECAPx10_ASAP7_75t_R FILLER_88_573 ();
 DECAPx4_ASAP7_75t_R FILLER_88_595 ();
 FILLER_ASAP7_75t_R FILLER_88_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_619 ();
 DECAPx10_ASAP7_75t_R FILLER_88_656 ();
 DECAPx10_ASAP7_75t_R FILLER_88_678 ();
 DECAPx10_ASAP7_75t_R FILLER_88_700 ();
 DECAPx6_ASAP7_75t_R FILLER_88_722 ();
 DECAPx2_ASAP7_75t_R FILLER_88_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_742 ();
 DECAPx10_ASAP7_75t_R FILLER_88_772 ();
 DECAPx4_ASAP7_75t_R FILLER_88_794 ();
 DECAPx10_ASAP7_75t_R FILLER_88_810 ();
 DECAPx6_ASAP7_75t_R FILLER_88_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_88_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_88_876 ();
 DECAPx2_ASAP7_75t_R FILLER_88_888 ();
 FILLER_ASAP7_75t_R FILLER_88_922 ();
 DECAPx10_ASAP7_75t_R FILLER_89_2 ();
 DECAPx10_ASAP7_75t_R FILLER_89_24 ();
 DECAPx10_ASAP7_75t_R FILLER_89_46 ();
 DECAPx10_ASAP7_75t_R FILLER_89_68 ();
 DECAPx4_ASAP7_75t_R FILLER_89_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_100 ();
 DECAPx4_ASAP7_75t_R FILLER_89_109 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_170 ();
 FILLER_ASAP7_75t_R FILLER_89_177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_211 ();
 DECAPx1_ASAP7_75t_R FILLER_89_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_230 ();
 DECAPx1_ASAP7_75t_R FILLER_89_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_243 ();
 DECAPx10_ASAP7_75t_R FILLER_89_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_292 ();
 DECAPx2_ASAP7_75t_R FILLER_89_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_350 ();
 DECAPx2_ASAP7_75t_R FILLER_89_356 ();
 FILLER_ASAP7_75t_R FILLER_89_362 ();
 FILLER_ASAP7_75t_R FILLER_89_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_419 ();
 DECAPx2_ASAP7_75t_R FILLER_89_446 ();
 FILLER_ASAP7_75t_R FILLER_89_463 ();
 DECAPx2_ASAP7_75t_R FILLER_89_471 ();
 FILLER_ASAP7_75t_R FILLER_89_477 ();
 FILLER_ASAP7_75t_R FILLER_89_489 ();
 DECAPx1_ASAP7_75t_R FILLER_89_519 ();
 DECAPx1_ASAP7_75t_R FILLER_89_530 ();
 DECAPx6_ASAP7_75t_R FILLER_89_561 ();
 DECAPx1_ASAP7_75t_R FILLER_89_575 ();
 DECAPx2_ASAP7_75t_R FILLER_89_585 ();
 FILLER_ASAP7_75t_R FILLER_89_591 ();
 DECAPx4_ASAP7_75t_R FILLER_89_605 ();
 DECAPx1_ASAP7_75t_R FILLER_89_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_630 ();
 DECAPx4_ASAP7_75t_R FILLER_89_669 ();
 FILLER_ASAP7_75t_R FILLER_89_679 ();
 DECAPx2_ASAP7_75t_R FILLER_89_687 ();
 DECAPx10_ASAP7_75t_R FILLER_89_696 ();
 DECAPx6_ASAP7_75t_R FILLER_89_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_732 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_743 ();
 DECAPx4_ASAP7_75t_R FILLER_89_762 ();
 FILLER_ASAP7_75t_R FILLER_89_772 ();
 DECAPx6_ASAP7_75t_R FILLER_89_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_89_800 ();
 DECAPx4_ASAP7_75t_R FILLER_89_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_89_829 ();
 DECAPx6_ASAP7_75t_R FILLER_89_836 ();
 FILLER_ASAP7_75t_R FILLER_89_850 ();
 DECAPx1_ASAP7_75t_R FILLER_89_866 ();
 DECAPx1_ASAP7_75t_R FILLER_89_930 ();
 DECAPx10_ASAP7_75t_R FILLER_90_2 ();
 DECAPx10_ASAP7_75t_R FILLER_90_24 ();
 DECAPx10_ASAP7_75t_R FILLER_90_46 ();
 DECAPx10_ASAP7_75t_R FILLER_90_68 ();
 DECAPx10_ASAP7_75t_R FILLER_90_90 ();
 FILLER_ASAP7_75t_R FILLER_90_112 ();
 FILLER_ASAP7_75t_R FILLER_90_140 ();
 FILLER_ASAP7_75t_R FILLER_90_150 ();
 DECAPx10_ASAP7_75t_R FILLER_90_158 ();
 DECAPx2_ASAP7_75t_R FILLER_90_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_193 ();
 DECAPx1_ASAP7_75t_R FILLER_90_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_229 ();
 DECAPx6_ASAP7_75t_R FILLER_90_238 ();
 DECAPx1_ASAP7_75t_R FILLER_90_252 ();
 FILLER_ASAP7_75t_R FILLER_90_262 ();
 FILLER_ASAP7_75t_R FILLER_90_267 ();
 DECAPx1_ASAP7_75t_R FILLER_90_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_307 ();
 DECAPx6_ASAP7_75t_R FILLER_90_340 ();
 DECAPx2_ASAP7_75t_R FILLER_90_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_385 ();
 FILLER_ASAP7_75t_R FILLER_90_412 ();
 DECAPx10_ASAP7_75t_R FILLER_90_471 ();
 DECAPx10_ASAP7_75t_R FILLER_90_493 ();
 DECAPx2_ASAP7_75t_R FILLER_90_515 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_521 ();
 DECAPx2_ASAP7_75t_R FILLER_90_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_550 ();
 FILLER_ASAP7_75t_R FILLER_90_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_589 ();
 DECAPx10_ASAP7_75t_R FILLER_90_616 ();
 FILLER_ASAP7_75t_R FILLER_90_638 ();
 DECAPx1_ASAP7_75t_R FILLER_90_653 ();
 DECAPx4_ASAP7_75t_R FILLER_90_665 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_675 ();
 DECAPx2_ASAP7_75t_R FILLER_90_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_716 ();
 FILLER_ASAP7_75t_R FILLER_90_733 ();
 DECAPx4_ASAP7_75t_R FILLER_90_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_755 ();
 DECAPx1_ASAP7_75t_R FILLER_90_763 ();
 FILLER_ASAP7_75t_R FILLER_90_770 ();
 FILLER_ASAP7_75t_R FILLER_90_784 ();
 DECAPx6_ASAP7_75t_R FILLER_90_798 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_812 ();
 DECAPx2_ASAP7_75t_R FILLER_90_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_90_847 ();
 DECAPx6_ASAP7_75t_R FILLER_90_854 ();
 FILLER_ASAP7_75t_R FILLER_90_868 ();
 FILLER_ASAP7_75t_R FILLER_90_896 ();
 DECAPx4_ASAP7_75t_R FILLER_90_904 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_90_914 ();
 DECAPx6_ASAP7_75t_R FILLER_90_920 ();
 DECAPx10_ASAP7_75t_R FILLER_91_2 ();
 DECAPx10_ASAP7_75t_R FILLER_91_24 ();
 DECAPx10_ASAP7_75t_R FILLER_91_46 ();
 DECAPx10_ASAP7_75t_R FILLER_91_68 ();
 DECAPx10_ASAP7_75t_R FILLER_91_90 ();
 DECAPx2_ASAP7_75t_R FILLER_91_112 ();
 DECAPx1_ASAP7_75t_R FILLER_91_124 ();
 DECAPx2_ASAP7_75t_R FILLER_91_131 ();
 DECAPx10_ASAP7_75t_R FILLER_91_140 ();
 DECAPx10_ASAP7_75t_R FILLER_91_162 ();
 DECAPx10_ASAP7_75t_R FILLER_91_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_206 ();
 DECAPx1_ASAP7_75t_R FILLER_91_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_217 ();
 DECAPx2_ASAP7_75t_R FILLER_91_221 ();
 DECAPx2_ASAP7_75t_R FILLER_91_239 ();
 DECAPx4_ASAP7_75t_R FILLER_91_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_295 ();
 DECAPx10_ASAP7_75t_R FILLER_91_299 ();
 FILLER_ASAP7_75t_R FILLER_91_321 ();
 DECAPx6_ASAP7_75t_R FILLER_91_326 ();
 DECAPx1_ASAP7_75t_R FILLER_91_340 ();
 FILLER_ASAP7_75t_R FILLER_91_350 ();
 FILLER_ASAP7_75t_R FILLER_91_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_422 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_433 ();
 DECAPx1_ASAP7_75t_R FILLER_91_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_449 ();
 DECAPx4_ASAP7_75t_R FILLER_91_456 ();
 DECAPx2_ASAP7_75t_R FILLER_91_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_481 ();
 FILLER_ASAP7_75t_R FILLER_91_485 ();
 DECAPx1_ASAP7_75t_R FILLER_91_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_496 ();
 FILLER_ASAP7_75t_R FILLER_91_502 ();
 FILLER_ASAP7_75t_R FILLER_91_514 ();
 DECAPx4_ASAP7_75t_R FILLER_91_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_533 ();
 DECAPx1_ASAP7_75t_R FILLER_91_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_565 ();
 DECAPx6_ASAP7_75t_R FILLER_91_603 ();
 DECAPx2_ASAP7_75t_R FILLER_91_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_623 ();
 DECAPx2_ASAP7_75t_R FILLER_91_636 ();
 DECAPx1_ASAP7_75t_R FILLER_91_680 ();
 FILLER_ASAP7_75t_R FILLER_91_694 ();
 DECAPx2_ASAP7_75t_R FILLER_91_728 ();
 DECAPx4_ASAP7_75t_R FILLER_91_740 ();
 FILLER_ASAP7_75t_R FILLER_91_750 ();
 DECAPx2_ASAP7_75t_R FILLER_91_778 ();
 DECAPx2_ASAP7_75t_R FILLER_91_790 ();
 DECAPx6_ASAP7_75t_R FILLER_91_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_816 ();
 DECAPx4_ASAP7_75t_R FILLER_91_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_91_833 ();
 DECAPx6_ASAP7_75t_R FILLER_91_863 ();
 DECAPx2_ASAP7_75t_R FILLER_91_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_883 ();
 DECAPx6_ASAP7_75t_R FILLER_91_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_91_924 ();
 FILLER_ASAP7_75t_R FILLER_91_927 ();
 DECAPx10_ASAP7_75t_R FILLER_92_2 ();
 DECAPx10_ASAP7_75t_R FILLER_92_24 ();
 DECAPx10_ASAP7_75t_R FILLER_92_46 ();
 DECAPx10_ASAP7_75t_R FILLER_92_68 ();
 DECAPx2_ASAP7_75t_R FILLER_92_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_105 ();
 DECAPx1_ASAP7_75t_R FILLER_92_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_115 ();
 DECAPx10_ASAP7_75t_R FILLER_92_122 ();
 FILLER_ASAP7_75t_R FILLER_92_144 ();
 DECAPx1_ASAP7_75t_R FILLER_92_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_156 ();
 DECAPx4_ASAP7_75t_R FILLER_92_169 ();
 FILLER_ASAP7_75t_R FILLER_92_179 ();
 DECAPx10_ASAP7_75t_R FILLER_92_184 ();
 DECAPx10_ASAP7_75t_R FILLER_92_206 ();
 DECAPx10_ASAP7_75t_R FILLER_92_228 ();
 FILLER_ASAP7_75t_R FILLER_92_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_258 ();
 DECAPx1_ASAP7_75t_R FILLER_92_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_266 ();
 DECAPx1_ASAP7_75t_R FILLER_92_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_283 ();
 DECAPx1_ASAP7_75t_R FILLER_92_296 ();
 DECAPx10_ASAP7_75t_R FILLER_92_303 ();
 DECAPx2_ASAP7_75t_R FILLER_92_325 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_331 ();
 DECAPx2_ASAP7_75t_R FILLER_92_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_374 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_396 ();
 FILLER_ASAP7_75t_R FILLER_92_407 ();
 DECAPx2_ASAP7_75t_R FILLER_92_428 ();
 FILLER_ASAP7_75t_R FILLER_92_434 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_461 ();
 DECAPx1_ASAP7_75t_R FILLER_92_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_468 ();
 FILLER_ASAP7_75t_R FILLER_92_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_514 ();
 DECAPx10_ASAP7_75t_R FILLER_92_535 ();
 FILLER_ASAP7_75t_R FILLER_92_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_567 ();
 FILLER_ASAP7_75t_R FILLER_92_623 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_641 ();
 DECAPx2_ASAP7_75t_R FILLER_92_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_656 ();
 FILLER_ASAP7_75t_R FILLER_92_660 ();
 DECAPx10_ASAP7_75t_R FILLER_92_708 ();
 DECAPx6_ASAP7_75t_R FILLER_92_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_744 ();
 DECAPx4_ASAP7_75t_R FILLER_92_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_761 ();
 DECAPx10_ASAP7_75t_R FILLER_92_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_789 ();
 DECAPx1_ASAP7_75t_R FILLER_92_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_800 ();
 FILLER_ASAP7_75t_R FILLER_92_810 ();
 DECAPx2_ASAP7_75t_R FILLER_92_818 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_92_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_92_830 ();
 DECAPx10_ASAP7_75t_R FILLER_92_844 ();
 DECAPx10_ASAP7_75t_R FILLER_92_866 ();
 DECAPx10_ASAP7_75t_R FILLER_92_888 ();
 DECAPx10_ASAP7_75t_R FILLER_92_910 ();
 FILLER_ASAP7_75t_R FILLER_92_932 ();
 DECAPx10_ASAP7_75t_R FILLER_93_2 ();
 DECAPx10_ASAP7_75t_R FILLER_93_24 ();
 DECAPx10_ASAP7_75t_R FILLER_93_46 ();
 DECAPx6_ASAP7_75t_R FILLER_93_68 ();
 FILLER_ASAP7_75t_R FILLER_93_82 ();
 DECAPx2_ASAP7_75t_R FILLER_93_139 ();
 DECAPx1_ASAP7_75t_R FILLER_93_192 ();
 DECAPx10_ASAP7_75t_R FILLER_93_210 ();
 DECAPx2_ASAP7_75t_R FILLER_93_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_238 ();
 DECAPx6_ASAP7_75t_R FILLER_93_257 ();
 DECAPx2_ASAP7_75t_R FILLER_93_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_328 ();
 DECAPx2_ASAP7_75t_R FILLER_93_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_338 ();
 DECAPx1_ASAP7_75t_R FILLER_93_345 ();
 FILLER_ASAP7_75t_R FILLER_93_352 ();
 DECAPx10_ASAP7_75t_R FILLER_93_360 ();
 DECAPx2_ASAP7_75t_R FILLER_93_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_388 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_421 ();
 FILLER_ASAP7_75t_R FILLER_93_460 ();
 FILLER_ASAP7_75t_R FILLER_93_493 ();
 DECAPx4_ASAP7_75t_R FILLER_93_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_543 ();
 DECAPx2_ASAP7_75t_R FILLER_93_547 ();
 FILLER_ASAP7_75t_R FILLER_93_553 ();
 DECAPx1_ASAP7_75t_R FILLER_93_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_565 ();
 DECAPx6_ASAP7_75t_R FILLER_93_576 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_618 ();
 DECAPx10_ASAP7_75t_R FILLER_93_639 ();
 DECAPx4_ASAP7_75t_R FILLER_93_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_671 ();
 FILLER_ASAP7_75t_R FILLER_93_684 ();
 DECAPx10_ASAP7_75t_R FILLER_93_695 ();
 DECAPx1_ASAP7_75t_R FILLER_93_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_721 ();
 DECAPx6_ASAP7_75t_R FILLER_93_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_742 ();
 DECAPx10_ASAP7_75t_R FILLER_93_756 ();
 DECAPx1_ASAP7_75t_R FILLER_93_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_782 ();
 DECAPx1_ASAP7_75t_R FILLER_93_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_802 ();
 DECAPx10_ASAP7_75t_R FILLER_93_822 ();
 DECAPx6_ASAP7_75t_R FILLER_93_844 ();
 DECAPx2_ASAP7_75t_R FILLER_93_858 ();
 DECAPx10_ASAP7_75t_R FILLER_93_872 ();
 DECAPx6_ASAP7_75t_R FILLER_93_894 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_93_908 ();
 DECAPx2_ASAP7_75t_R FILLER_93_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_93_924 ();
 FILLER_ASAP7_75t_R FILLER_93_927 ();
 DECAPx10_ASAP7_75t_R FILLER_94_2 ();
 DECAPx10_ASAP7_75t_R FILLER_94_24 ();
 DECAPx10_ASAP7_75t_R FILLER_94_46 ();
 DECAPx10_ASAP7_75t_R FILLER_94_68 ();
 DECAPx1_ASAP7_75t_R FILLER_94_90 ();
 FILLER_ASAP7_75t_R FILLER_94_100 ();
 DECAPx4_ASAP7_75t_R FILLER_94_105 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_115 ();
 DECAPx1_ASAP7_75t_R FILLER_94_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_157 ();
 FILLER_ASAP7_75t_R FILLER_94_196 ();
 DECAPx1_ASAP7_75t_R FILLER_94_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_217 ();
 DECAPx4_ASAP7_75t_R FILLER_94_221 ();
 FILLER_ASAP7_75t_R FILLER_94_231 ();
 DECAPx10_ASAP7_75t_R FILLER_94_259 ();
 DECAPx4_ASAP7_75t_R FILLER_94_281 ();
 FILLER_ASAP7_75t_R FILLER_94_291 ();
 FILLER_ASAP7_75t_R FILLER_94_296 ();
 DECAPx1_ASAP7_75t_R FILLER_94_310 ();
 DECAPx2_ASAP7_75t_R FILLER_94_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_346 ();
 DECAPx6_ASAP7_75t_R FILLER_94_356 ();
 DECAPx1_ASAP7_75t_R FILLER_94_370 ();
 FILLER_ASAP7_75t_R FILLER_94_445 ();
 FILLER_ASAP7_75t_R FILLER_94_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_464 ();
 DECAPx4_ASAP7_75t_R FILLER_94_500 ();
 DECAPx6_ASAP7_75t_R FILLER_94_513 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_527 ();
 FILLER_ASAP7_75t_R FILLER_94_556 ();
 DECAPx6_ASAP7_75t_R FILLER_94_565 ();
 DECAPx10_ASAP7_75t_R FILLER_94_584 ();
 DECAPx2_ASAP7_75t_R FILLER_94_606 ();
 FILLER_ASAP7_75t_R FILLER_94_612 ();
 DECAPx4_ASAP7_75t_R FILLER_94_630 ();
 DECAPx2_ASAP7_75t_R FILLER_94_649 ();
 FILLER_ASAP7_75t_R FILLER_94_655 ();
 DECAPx10_ASAP7_75t_R FILLER_94_667 ();
 DECAPx10_ASAP7_75t_R FILLER_94_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_742 ();
 DECAPx1_ASAP7_75t_R FILLER_94_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_776 ();
 FILLER_ASAP7_75t_R FILLER_94_785 ();
 DECAPx6_ASAP7_75t_R FILLER_94_790 ();
 FILLER_ASAP7_75t_R FILLER_94_804 ();
 DECAPx2_ASAP7_75t_R FILLER_94_824 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_830 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_94_847 ();
 DECAPx2_ASAP7_75t_R FILLER_94_891 ();
 DECAPx1_ASAP7_75t_R FILLER_94_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_94_907 ();
 DECAPx10_ASAP7_75t_R FILLER_95_2 ();
 DECAPx10_ASAP7_75t_R FILLER_95_24 ();
 DECAPx10_ASAP7_75t_R FILLER_95_46 ();
 DECAPx10_ASAP7_75t_R FILLER_95_68 ();
 DECAPx10_ASAP7_75t_R FILLER_95_90 ();
 DECAPx6_ASAP7_75t_R FILLER_95_112 ();
 DECAPx6_ASAP7_75t_R FILLER_95_154 ();
 DECAPx1_ASAP7_75t_R FILLER_95_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_179 ();
 DECAPx1_ASAP7_75t_R FILLER_95_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_202 ();
 FILLER_ASAP7_75t_R FILLER_95_232 ();
 DECAPx10_ASAP7_75t_R FILLER_95_256 ();
 DECAPx10_ASAP7_75t_R FILLER_95_278 ();
 DECAPx6_ASAP7_75t_R FILLER_95_300 ();
 DECAPx1_ASAP7_75t_R FILLER_95_314 ();
 DECAPx1_ASAP7_75t_R FILLER_95_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_341 ();
 FILLER_ASAP7_75t_R FILLER_95_363 ();
 FILLER_ASAP7_75t_R FILLER_95_387 ();
 DECAPx2_ASAP7_75t_R FILLER_95_411 ();
 FILLER_ASAP7_75t_R FILLER_95_417 ();
 DECAPx4_ASAP7_75t_R FILLER_95_462 ();
 FILLER_ASAP7_75t_R FILLER_95_472 ();
 DECAPx10_ASAP7_75t_R FILLER_95_479 ();
 DECAPx4_ASAP7_75t_R FILLER_95_501 ();
 DECAPx2_ASAP7_75t_R FILLER_95_516 ();
 DECAPx4_ASAP7_75t_R FILLER_95_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_537 ();
 DECAPx10_ASAP7_75t_R FILLER_95_549 ();
 DECAPx1_ASAP7_75t_R FILLER_95_571 ();
 DECAPx6_ASAP7_75t_R FILLER_95_591 ();
 FILLER_ASAP7_75t_R FILLER_95_605 ();
 DECAPx6_ASAP7_75t_R FILLER_95_613 ();
 DECAPx2_ASAP7_75t_R FILLER_95_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_650 ();
 DECAPx4_ASAP7_75t_R FILLER_95_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_691 ();
 DECAPx6_ASAP7_75t_R FILLER_95_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_755 ();
 DECAPx6_ASAP7_75t_R FILLER_95_799 ();
 DECAPx1_ASAP7_75t_R FILLER_95_813 ();
 DECAPx1_ASAP7_75t_R FILLER_95_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_95_849 ();
 DECAPx1_ASAP7_75t_R FILLER_95_868 ();
 DECAPx1_ASAP7_75t_R FILLER_95_888 ();
 DECAPx1_ASAP7_75t_R FILLER_95_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_95_933 ();
 DECAPx10_ASAP7_75t_R FILLER_96_2 ();
 DECAPx10_ASAP7_75t_R FILLER_96_24 ();
 DECAPx10_ASAP7_75t_R FILLER_96_46 ();
 DECAPx10_ASAP7_75t_R FILLER_96_68 ();
 DECAPx6_ASAP7_75t_R FILLER_96_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_104 ();
 DECAPx10_ASAP7_75t_R FILLER_96_167 ();
 DECAPx6_ASAP7_75t_R FILLER_96_189 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_203 ();
 DECAPx1_ASAP7_75t_R FILLER_96_244 ();
 FILLER_ASAP7_75t_R FILLER_96_260 ();
 DECAPx1_ASAP7_75t_R FILLER_96_276 ();
 FILLER_ASAP7_75t_R FILLER_96_286 ();
 DECAPx10_ASAP7_75t_R FILLER_96_297 ();
 DECAPx6_ASAP7_75t_R FILLER_96_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_369 ();
 FILLER_ASAP7_75t_R FILLER_96_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_459 ();
 DECAPx10_ASAP7_75t_R FILLER_96_474 ();
 FILLER_ASAP7_75t_R FILLER_96_496 ();
 DECAPx1_ASAP7_75t_R FILLER_96_509 ();
 DECAPx6_ASAP7_75t_R FILLER_96_525 ();
 DECAPx1_ASAP7_75t_R FILLER_96_539 ();
 DECAPx1_ASAP7_75t_R FILLER_96_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_553 ();
 FILLER_ASAP7_75t_R FILLER_96_561 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_598 ();
 DECAPx6_ASAP7_75t_R FILLER_96_621 ();
 DECAPx1_ASAP7_75t_R FILLER_96_635 ();
 DECAPx6_ASAP7_75t_R FILLER_96_645 ();
 DECAPx1_ASAP7_75t_R FILLER_96_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_663 ();
 DECAPx4_ASAP7_75t_R FILLER_96_667 ();
 DECAPx6_ASAP7_75t_R FILLER_96_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_96_717 ();
 DECAPx4_ASAP7_75t_R FILLER_96_726 ();
 FILLER_ASAP7_75t_R FILLER_96_736 ();
 DECAPx6_ASAP7_75t_R FILLER_96_741 ();
 FILLER_ASAP7_75t_R FILLER_96_755 ();
 DECAPx1_ASAP7_75t_R FILLER_96_783 ();
 DECAPx10_ASAP7_75t_R FILLER_96_790 ();
 DECAPx4_ASAP7_75t_R FILLER_96_812 ();
 FILLER_ASAP7_75t_R FILLER_96_822 ();
 DECAPx2_ASAP7_75t_R FILLER_96_844 ();
 DECAPx1_ASAP7_75t_R FILLER_96_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_874 ();
 DECAPx2_ASAP7_75t_R FILLER_96_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_96_933 ();
 DECAPx10_ASAP7_75t_R FILLER_97_2 ();
 DECAPx10_ASAP7_75t_R FILLER_97_24 ();
 DECAPx10_ASAP7_75t_R FILLER_97_46 ();
 DECAPx10_ASAP7_75t_R FILLER_97_68 ();
 DECAPx6_ASAP7_75t_R FILLER_97_90 ();
 FILLER_ASAP7_75t_R FILLER_97_104 ();
 DECAPx2_ASAP7_75t_R FILLER_97_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_144 ();
 FILLER_ASAP7_75t_R FILLER_97_153 ();
 DECAPx10_ASAP7_75t_R FILLER_97_161 ();
 DECAPx10_ASAP7_75t_R FILLER_97_183 ();
 DECAPx2_ASAP7_75t_R FILLER_97_205 ();
 FILLER_ASAP7_75t_R FILLER_97_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_240 ();
 DECAPx2_ASAP7_75t_R FILLER_97_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_315 ();
 FILLER_ASAP7_75t_R FILLER_97_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_397 ();
 FILLER_ASAP7_75t_R FILLER_97_429 ();
 FILLER_ASAP7_75t_R FILLER_97_446 ();
 DECAPx2_ASAP7_75t_R FILLER_97_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_480 ();
 DECAPx6_ASAP7_75t_R FILLER_97_533 ();
 DECAPx1_ASAP7_75t_R FILLER_97_580 ();
 FILLER_ASAP7_75t_R FILLER_97_624 ();
 DECAPx6_ASAP7_75t_R FILLER_97_636 ();
 DECAPx1_ASAP7_75t_R FILLER_97_682 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_699 ();
 FILLER_ASAP7_75t_R FILLER_97_716 ();
 DECAPx6_ASAP7_75t_R FILLER_97_738 ();
 DECAPx1_ASAP7_75t_R FILLER_97_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_756 ();
 DECAPx2_ASAP7_75t_R FILLER_97_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_97_769 ();
 DECAPx10_ASAP7_75t_R FILLER_97_778 ();
 DECAPx6_ASAP7_75t_R FILLER_97_800 ();
 DECAPx1_ASAP7_75t_R FILLER_97_814 ();
 DECAPx4_ASAP7_75t_R FILLER_97_831 ();
 DECAPx4_ASAP7_75t_R FILLER_97_857 ();
 FILLER_ASAP7_75t_R FILLER_97_867 ();
 DECAPx4_ASAP7_75t_R FILLER_97_875 ();
 DECAPx6_ASAP7_75t_R FILLER_97_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_913 ();
 DECAPx2_ASAP7_75t_R FILLER_97_917 ();
 FILLER_ASAP7_75t_R FILLER_97_923 ();
 DECAPx2_ASAP7_75t_R FILLER_97_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_97_933 ();
 DECAPx10_ASAP7_75t_R FILLER_98_2 ();
 DECAPx10_ASAP7_75t_R FILLER_98_24 ();
 DECAPx10_ASAP7_75t_R FILLER_98_46 ();
 DECAPx10_ASAP7_75t_R FILLER_98_68 ();
 DECAPx10_ASAP7_75t_R FILLER_98_90 ();
 DECAPx1_ASAP7_75t_R FILLER_98_112 ();
 FILLER_ASAP7_75t_R FILLER_98_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_142 ();
 DECAPx1_ASAP7_75t_R FILLER_98_161 ();
 DECAPx10_ASAP7_75t_R FILLER_98_200 ();
 DECAPx1_ASAP7_75t_R FILLER_98_222 ();
 DECAPx1_ASAP7_75t_R FILLER_98_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_233 ();
 DECAPx4_ASAP7_75t_R FILLER_98_242 ();
 FILLER_ASAP7_75t_R FILLER_98_252 ();
 FILLER_ASAP7_75t_R FILLER_98_263 ();
 DECAPx1_ASAP7_75t_R FILLER_98_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_297 ();
 FILLER_ASAP7_75t_R FILLER_98_301 ();
 DECAPx2_ASAP7_75t_R FILLER_98_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_327 ();
 FILLER_ASAP7_75t_R FILLER_98_336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_354 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_368 ();
 DECAPx1_ASAP7_75t_R FILLER_98_381 ();
 DECAPx2_ASAP7_75t_R FILLER_98_391 ();
 DECAPx6_ASAP7_75t_R FILLER_98_407 ();
 DECAPx2_ASAP7_75t_R FILLER_98_421 ();
 DECAPx2_ASAP7_75t_R FILLER_98_430 ();
 FILLER_ASAP7_75t_R FILLER_98_436 ();
 DECAPx2_ASAP7_75t_R FILLER_98_445 ();
 DECAPx1_ASAP7_75t_R FILLER_98_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_461 ();
 FILLER_ASAP7_75t_R FILLER_98_470 ();
 FILLER_ASAP7_75t_R FILLER_98_478 ();
 FILLER_ASAP7_75t_R FILLER_98_550 ();
 DECAPx2_ASAP7_75t_R FILLER_98_572 ();
 FILLER_ASAP7_75t_R FILLER_98_578 ();
 DECAPx4_ASAP7_75t_R FILLER_98_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_596 ();
 DECAPx4_ASAP7_75t_R FILLER_98_611 ();
 DECAPx10_ASAP7_75t_R FILLER_98_649 ();
 DECAPx2_ASAP7_75t_R FILLER_98_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_677 ();
 DECAPx6_ASAP7_75t_R FILLER_98_686 ();
 DECAPx2_ASAP7_75t_R FILLER_98_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_706 ();
 DECAPx2_ASAP7_75t_R FILLER_98_719 ();
 FILLER_ASAP7_75t_R FILLER_98_725 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_732 ();
 DECAPx10_ASAP7_75t_R FILLER_98_745 ();
 DECAPx10_ASAP7_75t_R FILLER_98_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_98_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_798 ();
 DECAPx1_ASAP7_75t_R FILLER_98_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_817 ();
 DECAPx10_ASAP7_75t_R FILLER_98_821 ();
 DECAPx10_ASAP7_75t_R FILLER_98_843 ();
 DECAPx10_ASAP7_75t_R FILLER_98_865 ();
 DECAPx6_ASAP7_75t_R FILLER_98_887 ();
 DECAPx2_ASAP7_75t_R FILLER_98_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_98_907 ();
 DECAPx10_ASAP7_75t_R FILLER_99_2 ();
 DECAPx10_ASAP7_75t_R FILLER_99_24 ();
 DECAPx10_ASAP7_75t_R FILLER_99_46 ();
 DECAPx6_ASAP7_75t_R FILLER_99_68 ();
 FILLER_ASAP7_75t_R FILLER_99_82 ();
 DECAPx2_ASAP7_75t_R FILLER_99_110 ();
 DECAPx1_ASAP7_75t_R FILLER_99_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_172 ();
 FILLER_ASAP7_75t_R FILLER_99_179 ();
 DECAPx10_ASAP7_75t_R FILLER_99_207 ();
 DECAPx6_ASAP7_75t_R FILLER_99_229 ();
 DECAPx6_ASAP7_75t_R FILLER_99_272 ();
 DECAPx2_ASAP7_75t_R FILLER_99_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_292 ();
 DECAPx10_ASAP7_75t_R FILLER_99_327 ();
 FILLER_ASAP7_75t_R FILLER_99_349 ();
 DECAPx10_ASAP7_75t_R FILLER_99_357 ();
 DECAPx2_ASAP7_75t_R FILLER_99_407 ();
 DECAPx6_ASAP7_75t_R FILLER_99_439 ();
 DECAPx1_ASAP7_75t_R FILLER_99_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_457 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_492 ();
 DECAPx4_ASAP7_75t_R FILLER_99_506 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_524 ();
 FILLER_ASAP7_75t_R FILLER_99_533 ();
 DECAPx2_ASAP7_75t_R FILLER_99_538 ();
 DECAPx2_ASAP7_75t_R FILLER_99_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_576 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_99_585 ();
 DECAPx6_ASAP7_75t_R FILLER_99_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_610 ();
 DECAPx1_ASAP7_75t_R FILLER_99_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_641 ();
 DECAPx10_ASAP7_75t_R FILLER_99_674 ();
 DECAPx10_ASAP7_75t_R FILLER_99_696 ();
 DECAPx2_ASAP7_75t_R FILLER_99_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_724 ();
 DECAPx4_ASAP7_75t_R FILLER_99_733 ();
 DECAPx1_ASAP7_75t_R FILLER_99_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_760 ();
 DECAPx2_ASAP7_75t_R FILLER_99_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_778 ();
 FILLER_ASAP7_75t_R FILLER_99_787 ();
 DECAPx10_ASAP7_75t_R FILLER_99_821 ();
 DECAPx6_ASAP7_75t_R FILLER_99_843 ();
 DECAPx1_ASAP7_75t_R FILLER_99_857 ();
 DECAPx10_ASAP7_75t_R FILLER_99_867 ();
 DECAPx10_ASAP7_75t_R FILLER_99_889 ();
 DECAPx6_ASAP7_75t_R FILLER_99_911 ();
 DECAPx2_ASAP7_75t_R FILLER_99_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_99_933 ();
 DECAPx10_ASAP7_75t_R FILLER_100_2 ();
 DECAPx10_ASAP7_75t_R FILLER_100_24 ();
 DECAPx10_ASAP7_75t_R FILLER_100_46 ();
 DECAPx10_ASAP7_75t_R FILLER_100_68 ();
 DECAPx2_ASAP7_75t_R FILLER_100_90 ();
 FILLER_ASAP7_75t_R FILLER_100_96 ();
 DECAPx1_ASAP7_75t_R FILLER_100_101 ();
 DECAPx10_ASAP7_75t_R FILLER_100_108 ();
 DECAPx4_ASAP7_75t_R FILLER_100_133 ();
 FILLER_ASAP7_75t_R FILLER_100_143 ();
 DECAPx2_ASAP7_75t_R FILLER_100_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_166 ();
 DECAPx2_ASAP7_75t_R FILLER_100_173 ();
 FILLER_ASAP7_75t_R FILLER_100_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_193 ();
 FILLER_ASAP7_75t_R FILLER_100_214 ();
 DECAPx2_ASAP7_75t_R FILLER_100_222 ();
 DECAPx6_ASAP7_75t_R FILLER_100_231 ();
 DECAPx1_ASAP7_75t_R FILLER_100_245 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_255 ();
 DECAPx10_ASAP7_75t_R FILLER_100_261 ();
 DECAPx6_ASAP7_75t_R FILLER_100_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_297 ();
 DECAPx1_ASAP7_75t_R FILLER_100_304 ();
 DECAPx4_ASAP7_75t_R FILLER_100_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_330 ();
 DECAPx10_ASAP7_75t_R FILLER_100_342 ();
 DECAPx4_ASAP7_75t_R FILLER_100_364 ();
 DECAPx1_ASAP7_75t_R FILLER_100_410 ();
 DECAPx6_ASAP7_75t_R FILLER_100_448 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_470 ();
 FILLER_ASAP7_75t_R FILLER_100_476 ();
 DECAPx2_ASAP7_75t_R FILLER_100_481 ();
 FILLER_ASAP7_75t_R FILLER_100_487 ();
 DECAPx10_ASAP7_75t_R FILLER_100_495 ();
 DECAPx6_ASAP7_75t_R FILLER_100_517 ();
 FILLER_ASAP7_75t_R FILLER_100_531 ();
 DECAPx6_ASAP7_75t_R FILLER_100_539 ();
 DECAPx1_ASAP7_75t_R FILLER_100_560 ();
 DECAPx4_ASAP7_75t_R FILLER_100_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_577 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_586 ();
 DECAPx2_ASAP7_75t_R FILLER_100_609 ();
 FILLER_ASAP7_75t_R FILLER_100_624 ();
 DECAPx2_ASAP7_75t_R FILLER_100_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_638 ();
 DECAPx1_ASAP7_75t_R FILLER_100_648 ();
 DECAPx1_ASAP7_75t_R FILLER_100_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_662 ();
 DECAPx4_ASAP7_75t_R FILLER_100_675 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_685 ();
 DECAPx2_ASAP7_75t_R FILLER_100_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_725 ();
 DECAPx2_ASAP7_75t_R FILLER_100_733 ();
 DECAPx1_ASAP7_75t_R FILLER_100_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_100_793 ();
 FILLER_ASAP7_75t_R FILLER_100_803 ();
 DECAPx2_ASAP7_75t_R FILLER_100_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_820 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_830 ();
 DECAPx2_ASAP7_75t_R FILLER_100_845 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_851 ();
 FILLER_ASAP7_75t_R FILLER_100_893 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_100_910 ();
 FILLER_ASAP7_75t_R FILLER_100_932 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_2 ();
 DECAPx10_ASAP7_75t_R FILLER_101_13 ();
 DECAPx10_ASAP7_75t_R FILLER_101_35 ();
 DECAPx10_ASAP7_75t_R FILLER_101_57 ();
 DECAPx10_ASAP7_75t_R FILLER_101_79 ();
 DECAPx10_ASAP7_75t_R FILLER_101_101 ();
 DECAPx10_ASAP7_75t_R FILLER_101_123 ();
 DECAPx6_ASAP7_75t_R FILLER_101_145 ();
 DECAPx1_ASAP7_75t_R FILLER_101_159 ();
 DECAPx6_ASAP7_75t_R FILLER_101_178 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_192 ();
 DECAPx1_ASAP7_75t_R FILLER_101_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_213 ();
 DECAPx10_ASAP7_75t_R FILLER_101_243 ();
 DECAPx2_ASAP7_75t_R FILLER_101_265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_271 ();
 DECAPx6_ASAP7_75t_R FILLER_101_282 ();
 DECAPx2_ASAP7_75t_R FILLER_101_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_372 ();
 DECAPx1_ASAP7_75t_R FILLER_101_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_446 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_455 ();
 DECAPx10_ASAP7_75t_R FILLER_101_466 ();
 DECAPx6_ASAP7_75t_R FILLER_101_494 ();
 FILLER_ASAP7_75t_R FILLER_101_508 ();
 DECAPx6_ASAP7_75t_R FILLER_101_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_532 ();
 DECAPx1_ASAP7_75t_R FILLER_101_541 ();
 DECAPx1_ASAP7_75t_R FILLER_101_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_556 ();
 DECAPx4_ASAP7_75t_R FILLER_101_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_572 ();
 DECAPx2_ASAP7_75t_R FILLER_101_599 ();
 FILLER_ASAP7_75t_R FILLER_101_605 ();
 DECAPx10_ASAP7_75t_R FILLER_101_619 ();
 DECAPx1_ASAP7_75t_R FILLER_101_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_645 ();
 DECAPx1_ASAP7_75t_R FILLER_101_672 ();
 DECAPx1_ASAP7_75t_R FILLER_101_711 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_736 ();
 FILLER_ASAP7_75t_R FILLER_101_759 ();
 DECAPx10_ASAP7_75t_R FILLER_101_773 ();
 DECAPx6_ASAP7_75t_R FILLER_101_795 ();
 DECAPx1_ASAP7_75t_R FILLER_101_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_820 ();
 DECAPx1_ASAP7_75t_R FILLER_101_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_865 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_101_902 ();
 DECAPx2_ASAP7_75t_R FILLER_101_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_924 ();
 DECAPx2_ASAP7_75t_R FILLER_101_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_101_933 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_2 ();
 DECAPx10_ASAP7_75t_R FILLER_102_22 ();
 DECAPx10_ASAP7_75t_R FILLER_102_44 ();
 DECAPx6_ASAP7_75t_R FILLER_102_66 ();
 DECAPx2_ASAP7_75t_R FILLER_102_80 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_86 ();
 DECAPx6_ASAP7_75t_R FILLER_102_99 ();
 DECAPx1_ASAP7_75t_R FILLER_102_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_126 ();
 DECAPx10_ASAP7_75t_R FILLER_102_130 ();
 DECAPx2_ASAP7_75t_R FILLER_102_152 ();
 FILLER_ASAP7_75t_R FILLER_102_158 ();
 DECAPx6_ASAP7_75t_R FILLER_102_186 ();
 DECAPx2_ASAP7_75t_R FILLER_102_206 ();
 FILLER_ASAP7_75t_R FILLER_102_212 ();
 DECAPx1_ASAP7_75t_R FILLER_102_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_224 ();
 FILLER_ASAP7_75t_R FILLER_102_231 ();
 DECAPx1_ASAP7_75t_R FILLER_102_239 ();
 DECAPx1_ASAP7_75t_R FILLER_102_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_283 ();
 DECAPx4_ASAP7_75t_R FILLER_102_316 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_326 ();
 DECAPx4_ASAP7_75t_R FILLER_102_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_383 ();
 DECAPx4_ASAP7_75t_R FILLER_102_387 ();
 DECAPx10_ASAP7_75t_R FILLER_102_411 ();
 DECAPx4_ASAP7_75t_R FILLER_102_433 ();
 FILLER_ASAP7_75t_R FILLER_102_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_455 ();
 DECAPx10_ASAP7_75t_R FILLER_102_464 ();
 FILLER_ASAP7_75t_R FILLER_102_486 ();
 DECAPx1_ASAP7_75t_R FILLER_102_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_500 ();
 FILLER_ASAP7_75t_R FILLER_102_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_523 ();
 DECAPx4_ASAP7_75t_R FILLER_102_532 ();
 FILLER_ASAP7_75t_R FILLER_102_542 ();
 DECAPx1_ASAP7_75t_R FILLER_102_564 ();
 DECAPx10_ASAP7_75t_R FILLER_102_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_605 ();
 DECAPx4_ASAP7_75t_R FILLER_102_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_623 ();
 DECAPx10_ASAP7_75t_R FILLER_102_630 ();
 DECAPx2_ASAP7_75t_R FILLER_102_652 ();
 DECAPx2_ASAP7_75t_R FILLER_102_667 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_673 ();
 DECAPx1_ASAP7_75t_R FILLER_102_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_684 ();
 DECAPx2_ASAP7_75t_R FILLER_102_688 ();
 FILLER_ASAP7_75t_R FILLER_102_694 ();
 DECAPx2_ASAP7_75t_R FILLER_102_714 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_720 ();
 DECAPx10_ASAP7_75t_R FILLER_102_728 ();
 DECAPx6_ASAP7_75t_R FILLER_102_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_774 ();
 DECAPx10_ASAP7_75t_R FILLER_102_784 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_840 ();
 DECAPx2_ASAP7_75t_R FILLER_102_847 ();
 FILLER_ASAP7_75t_R FILLER_102_853 ();
 FILLER_ASAP7_75t_R FILLER_102_862 ();
 DECAPx2_ASAP7_75t_R FILLER_102_867 ();
 FILLER_ASAP7_75t_R FILLER_102_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_102_887 ();
 DECAPx4_ASAP7_75t_R FILLER_102_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_102_903 ();
 DECAPx1_ASAP7_75t_R FILLER_102_930 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_2 ();
 DECAPx10_ASAP7_75t_R FILLER_103_14 ();
 DECAPx10_ASAP7_75t_R FILLER_103_36 ();
 DECAPx10_ASAP7_75t_R FILLER_103_58 ();
 DECAPx2_ASAP7_75t_R FILLER_103_80 ();
 DECAPx2_ASAP7_75t_R FILLER_103_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_108 ();
 DECAPx10_ASAP7_75t_R FILLER_103_141 ();
 DECAPx6_ASAP7_75t_R FILLER_103_163 ();
 DECAPx6_ASAP7_75t_R FILLER_103_183 ();
 DECAPx2_ASAP7_75t_R FILLER_103_197 ();
 DECAPx4_ASAP7_75t_R FILLER_103_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_220 ();
 DECAPx1_ASAP7_75t_R FILLER_103_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_285 ();
 DECAPx1_ASAP7_75t_R FILLER_103_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_302 ();
 DECAPx10_ASAP7_75t_R FILLER_103_312 ();
 DECAPx4_ASAP7_75t_R FILLER_103_334 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_352 ();
 DECAPx2_ASAP7_75t_R FILLER_103_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_369 ();
 DECAPx4_ASAP7_75t_R FILLER_103_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_406 ();
 DECAPx6_ASAP7_75t_R FILLER_103_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_443 ();
 DECAPx10_ASAP7_75t_R FILLER_103_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_474 ();
 DECAPx4_ASAP7_75t_R FILLER_103_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_499 ();
 DECAPx4_ASAP7_75t_R FILLER_103_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_516 ();
 DECAPx4_ASAP7_75t_R FILLER_103_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_611 ();
 DECAPx2_ASAP7_75t_R FILLER_103_620 ();
 FILLER_ASAP7_75t_R FILLER_103_626 ();
 DECAPx1_ASAP7_75t_R FILLER_103_634 ();
 DECAPx1_ASAP7_75t_R FILLER_103_644 ();
 DECAPx6_ASAP7_75t_R FILLER_103_651 ();
 DECAPx2_ASAP7_75t_R FILLER_103_665 ();
 DECAPx4_ASAP7_75t_R FILLER_103_697 ();
 DECAPx6_ASAP7_75t_R FILLER_103_713 ();
 DECAPx2_ASAP7_75t_R FILLER_103_727 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_752 ();
 DECAPx2_ASAP7_75t_R FILLER_103_758 ();
 DECAPx2_ASAP7_75t_R FILLER_103_772 ();
 DECAPx10_ASAP7_75t_R FILLER_103_789 ();
 DECAPx10_ASAP7_75t_R FILLER_103_811 ();
 DECAPx6_ASAP7_75t_R FILLER_103_833 ();
 FILLER_ASAP7_75t_R FILLER_103_847 ();
 DECAPx2_ASAP7_75t_R FILLER_103_878 ();
 DECAPx6_ASAP7_75t_R FILLER_103_898 ();
 DECAPx2_ASAP7_75t_R FILLER_103_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_918 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_103_922 ();
 DECAPx2_ASAP7_75t_R FILLER_103_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_103_933 ();
 DECAPx10_ASAP7_75t_R FILLER_104_5 ();
 DECAPx10_ASAP7_75t_R FILLER_104_27 ();
 DECAPx10_ASAP7_75t_R FILLER_104_49 ();
 DECAPx2_ASAP7_75t_R FILLER_104_71 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_103 ();
 DECAPx1_ASAP7_75t_R FILLER_104_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_130 ();
 DECAPx6_ASAP7_75t_R FILLER_104_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_174 ();
 DECAPx10_ASAP7_75t_R FILLER_104_189 ();
 DECAPx6_ASAP7_75t_R FILLER_104_229 ();
 DECAPx2_ASAP7_75t_R FILLER_104_243 ();
 DECAPx2_ASAP7_75t_R FILLER_104_255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_261 ();
 FILLER_ASAP7_75t_R FILLER_104_270 ();
 DECAPx10_ASAP7_75t_R FILLER_104_296 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_318 ();
 DECAPx2_ASAP7_75t_R FILLER_104_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_345 ();
 DECAPx10_ASAP7_75t_R FILLER_104_354 ();
 DECAPx10_ASAP7_75t_R FILLER_104_376 ();
 DECAPx6_ASAP7_75t_R FILLER_104_398 ();
 FILLER_ASAP7_75t_R FILLER_104_412 ();
 DECAPx1_ASAP7_75t_R FILLER_104_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_447 ();
 DECAPx2_ASAP7_75t_R FILLER_104_456 ();
 DECAPx1_ASAP7_75t_R FILLER_104_508 ();
 DECAPx2_ASAP7_75t_R FILLER_104_520 ();
 DECAPx1_ASAP7_75t_R FILLER_104_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_541 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_549 ();
 DECAPx1_ASAP7_75t_R FILLER_104_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_576 ();
 DECAPx1_ASAP7_75t_R FILLER_104_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_589 ();
 DECAPx2_ASAP7_75t_R FILLER_104_596 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_623 ();
 DECAPx4_ASAP7_75t_R FILLER_104_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_662 ();
 DECAPx4_ASAP7_75t_R FILLER_104_669 ();
 FILLER_ASAP7_75t_R FILLER_104_685 ();
 DECAPx4_ASAP7_75t_R FILLER_104_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_709 ();
 DECAPx2_ASAP7_75t_R FILLER_104_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_104_723 ();
 DECAPx10_ASAP7_75t_R FILLER_104_730 ();
 DECAPx10_ASAP7_75t_R FILLER_104_752 ();
 DECAPx6_ASAP7_75t_R FILLER_104_774 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_794 ();
 DECAPx10_ASAP7_75t_R FILLER_104_813 ();
 DECAPx6_ASAP7_75t_R FILLER_104_835 ();
 FILLER_ASAP7_75t_R FILLER_104_849 ();
 DECAPx10_ASAP7_75t_R FILLER_104_861 ();
 DECAPx4_ASAP7_75t_R FILLER_104_883 ();
 DECAPx6_ASAP7_75t_R FILLER_104_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_104_933 ();
 DECAPx10_ASAP7_75t_R FILLER_105_2 ();
 DECAPx10_ASAP7_75t_R FILLER_105_24 ();
 DECAPx10_ASAP7_75t_R FILLER_105_46 ();
 DECAPx4_ASAP7_75t_R FILLER_105_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_78 ();
 DECAPx6_ASAP7_75t_R FILLER_105_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_101 ();
 DECAPx10_ASAP7_75t_R FILLER_105_108 ();
 DECAPx2_ASAP7_75t_R FILLER_105_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_136 ();
 FILLER_ASAP7_75t_R FILLER_105_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_191 ();
 DECAPx2_ASAP7_75t_R FILLER_105_198 ();
 DECAPx4_ASAP7_75t_R FILLER_105_236 ();
 DECAPx2_ASAP7_75t_R FILLER_105_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_269 ();
 DECAPx1_ASAP7_75t_R FILLER_105_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_277 ();
 FILLER_ASAP7_75t_R FILLER_105_339 ();
 DECAPx10_ASAP7_75t_R FILLER_105_363 ();
 DECAPx2_ASAP7_75t_R FILLER_105_385 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_391 ();
 DECAPx1_ASAP7_75t_R FILLER_105_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_440 ();
 DECAPx1_ASAP7_75t_R FILLER_105_467 ();
 DECAPx10_ASAP7_75t_R FILLER_105_489 ();
 DECAPx6_ASAP7_75t_R FILLER_105_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_525 ();
 DECAPx4_ASAP7_75t_R FILLER_105_534 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_544 ();
 DECAPx6_ASAP7_75t_R FILLER_105_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_568 ();
 DECAPx4_ASAP7_75t_R FILLER_105_577 ();
 DECAPx6_ASAP7_75t_R FILLER_105_593 ();
 DECAPx2_ASAP7_75t_R FILLER_105_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_613 ();
 DECAPx2_ASAP7_75t_R FILLER_105_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_636 ();
 DECAPx10_ASAP7_75t_R FILLER_105_663 ();
 DECAPx10_ASAP7_75t_R FILLER_105_685 ();
 DECAPx2_ASAP7_75t_R FILLER_105_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_720 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_105_772 ();
 DECAPx6_ASAP7_75t_R FILLER_105_787 ();
 DECAPx4_ASAP7_75t_R FILLER_105_808 ();
 FILLER_ASAP7_75t_R FILLER_105_818 ();
 DECAPx1_ASAP7_75t_R FILLER_105_831 ();
 DECAPx10_ASAP7_75t_R FILLER_105_840 ();
 DECAPx10_ASAP7_75t_R FILLER_105_862 ();
 DECAPx10_ASAP7_75t_R FILLER_105_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_906 ();
 DECAPx1_ASAP7_75t_R FILLER_105_910 ();
 DECAPx1_ASAP7_75t_R FILLER_105_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_105_921 ();
 FILLER_ASAP7_75t_R FILLER_105_927 ();
 DECAPx10_ASAP7_75t_R FILLER_106_2 ();
 DECAPx10_ASAP7_75t_R FILLER_106_24 ();
 DECAPx10_ASAP7_75t_R FILLER_106_46 ();
 DECAPx10_ASAP7_75t_R FILLER_106_68 ();
 DECAPx10_ASAP7_75t_R FILLER_106_90 ();
 DECAPx10_ASAP7_75t_R FILLER_106_112 ();
 DECAPx1_ASAP7_75t_R FILLER_106_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_144 ();
 DECAPx1_ASAP7_75t_R FILLER_106_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_161 ();
 DECAPx4_ASAP7_75t_R FILLER_106_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_205 ();
 DECAPx4_ASAP7_75t_R FILLER_106_211 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_221 ();
 DECAPx2_ASAP7_75t_R FILLER_106_227 ();
 DECAPx1_ASAP7_75t_R FILLER_106_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_250 ();
 DECAPx10_ASAP7_75t_R FILLER_106_257 ();
 DECAPx6_ASAP7_75t_R FILLER_106_279 ();
 DECAPx6_ASAP7_75t_R FILLER_106_302 ();
 FILLER_ASAP7_75t_R FILLER_106_316 ();
 DECAPx1_ASAP7_75t_R FILLER_106_330 ();
 FILLER_ASAP7_75t_R FILLER_106_409 ();
 DECAPx2_ASAP7_75t_R FILLER_106_417 ();
 FILLER_ASAP7_75t_R FILLER_106_423 ();
 DECAPx6_ASAP7_75t_R FILLER_106_428 ();
 DECAPx1_ASAP7_75t_R FILLER_106_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_452 ();
 DECAPx1_ASAP7_75t_R FILLER_106_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_464 ();
 DECAPx10_ASAP7_75t_R FILLER_106_471 ();
 DECAPx2_ASAP7_75t_R FILLER_106_493 ();
 DECAPx10_ASAP7_75t_R FILLER_106_510 ();
 DECAPx10_ASAP7_75t_R FILLER_106_532 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_554 ();
 DECAPx2_ASAP7_75t_R FILLER_106_560 ();
 DECAPx2_ASAP7_75t_R FILLER_106_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_582 ();
 DECAPx10_ASAP7_75t_R FILLER_106_597 ();
 DECAPx10_ASAP7_75t_R FILLER_106_619 ();
 DECAPx1_ASAP7_75t_R FILLER_106_641 ();
 DECAPx1_ASAP7_75t_R FILLER_106_657 ();
 DECAPx1_ASAP7_75t_R FILLER_106_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_674 ();
 DECAPx6_ASAP7_75t_R FILLER_106_678 ();
 DECAPx1_ASAP7_75t_R FILLER_106_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_696 ();
 DECAPx1_ASAP7_75t_R FILLER_106_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_716 ();
 DECAPx2_ASAP7_75t_R FILLER_106_727 ();
 FILLER_ASAP7_75t_R FILLER_106_733 ();
 DECAPx2_ASAP7_75t_R FILLER_106_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_783 ();
 FILLER_ASAP7_75t_R FILLER_106_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_106_872 ();
 DECAPx2_ASAP7_75t_R FILLER_106_889 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_895 ();
 DECAPx4_ASAP7_75t_R FILLER_106_906 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_106_916 ();
 DECAPx10_ASAP7_75t_R FILLER_107_2 ();
 DECAPx10_ASAP7_75t_R FILLER_107_24 ();
 DECAPx10_ASAP7_75t_R FILLER_107_46 ();
 DECAPx6_ASAP7_75t_R FILLER_107_68 ();
 DECAPx1_ASAP7_75t_R FILLER_107_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_86 ();
 DECAPx4_ASAP7_75t_R FILLER_107_90 ();
 FILLER_ASAP7_75t_R FILLER_107_106 ();
 DECAPx1_ASAP7_75t_R FILLER_107_114 ();
 DECAPx6_ASAP7_75t_R FILLER_107_144 ();
 DECAPx2_ASAP7_75t_R FILLER_107_158 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_164 ();
 DECAPx10_ASAP7_75t_R FILLER_107_171 ();
 FILLER_ASAP7_75t_R FILLER_107_222 ();
 DECAPx4_ASAP7_75t_R FILLER_107_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_246 ();
 DECAPx6_ASAP7_75t_R FILLER_107_279 ();
 FILLER_ASAP7_75t_R FILLER_107_293 ();
 DECAPx4_ASAP7_75t_R FILLER_107_302 ();
 FILLER_ASAP7_75t_R FILLER_107_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_348 ();
 FILLER_ASAP7_75t_R FILLER_107_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_391 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_107_415 ();
 DECAPx4_ASAP7_75t_R FILLER_107_425 ();
 DECAPx10_ASAP7_75t_R FILLER_107_465 ();
 DECAPx1_ASAP7_75t_R FILLER_107_487 ();
 DECAPx6_ASAP7_75t_R FILLER_107_517 ();
 FILLER_ASAP7_75t_R FILLER_107_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_542 ();
 DECAPx1_ASAP7_75t_R FILLER_107_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_573 ();
 DECAPx10_ASAP7_75t_R FILLER_107_580 ();
 DECAPx6_ASAP7_75t_R FILLER_107_602 ();
 DECAPx1_ASAP7_75t_R FILLER_107_616 ();
 DECAPx6_ASAP7_75t_R FILLER_107_641 ();
 DECAPx1_ASAP7_75t_R FILLER_107_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_659 ();
 DECAPx6_ASAP7_75t_R FILLER_107_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_715 ();
 DECAPx6_ASAP7_75t_R FILLER_107_722 ();
 DECAPx2_ASAP7_75t_R FILLER_107_741 ();
 DECAPx2_ASAP7_75t_R FILLER_107_753 ();
 FILLER_ASAP7_75t_R FILLER_107_759 ();
 DECAPx1_ASAP7_75t_R FILLER_107_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_771 ();
 DECAPx1_ASAP7_75t_R FILLER_107_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_788 ();
 FILLER_ASAP7_75t_R FILLER_107_805 ();
 DECAPx1_ASAP7_75t_R FILLER_107_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_107_924 ();
 FILLER_ASAP7_75t_R FILLER_107_927 ();
 DECAPx10_ASAP7_75t_R FILLER_108_2 ();
 DECAPx10_ASAP7_75t_R FILLER_108_24 ();
 DECAPx10_ASAP7_75t_R FILLER_108_46 ();
 FILLER_ASAP7_75t_R FILLER_108_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_134 ();
 DECAPx10_ASAP7_75t_R FILLER_108_144 ();
 FILLER_ASAP7_75t_R FILLER_108_166 ();
 DECAPx10_ASAP7_75t_R FILLER_108_174 ();
 DECAPx6_ASAP7_75t_R FILLER_108_202 ();
 DECAPx1_ASAP7_75t_R FILLER_108_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_220 ();
 FILLER_ASAP7_75t_R FILLER_108_247 ();
 DECAPx2_ASAP7_75t_R FILLER_108_293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_325 ();
 DECAPx6_ASAP7_75t_R FILLER_108_331 ();
 FILLER_ASAP7_75t_R FILLER_108_345 ();
 DECAPx2_ASAP7_75t_R FILLER_108_352 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_358 ();
 DECAPx6_ASAP7_75t_R FILLER_108_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_378 ();
 DECAPx6_ASAP7_75t_R FILLER_108_394 ();
 DECAPx1_ASAP7_75t_R FILLER_108_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_461 ();
 DECAPx6_ASAP7_75t_R FILLER_108_469 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_483 ();
 DECAPx1_ASAP7_75t_R FILLER_108_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_502 ();
 FILLER_ASAP7_75t_R FILLER_108_522 ();
 DECAPx10_ASAP7_75t_R FILLER_108_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_584 ();
 DECAPx4_ASAP7_75t_R FILLER_108_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_601 ();
 DECAPx4_ASAP7_75t_R FILLER_108_640 ();
 FILLER_ASAP7_75t_R FILLER_108_679 ();
 DECAPx4_ASAP7_75t_R FILLER_108_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_724 ();
 DECAPx10_ASAP7_75t_R FILLER_108_744 ();
 DECAPx4_ASAP7_75t_R FILLER_108_766 ();
 FILLER_ASAP7_75t_R FILLER_108_776 ();
 DECAPx2_ASAP7_75t_R FILLER_108_800 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_108_806 ();
 DECAPx6_ASAP7_75t_R FILLER_108_819 ();
 DECAPx1_ASAP7_75t_R FILLER_108_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_108_907 ();
 DECAPx10_ASAP7_75t_R FILLER_109_2 ();
 DECAPx10_ASAP7_75t_R FILLER_109_24 ();
 DECAPx10_ASAP7_75t_R FILLER_109_46 ();
 DECAPx1_ASAP7_75t_R FILLER_109_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_72 ();
 DECAPx4_ASAP7_75t_R FILLER_109_111 ();
 DECAPx1_ASAP7_75t_R FILLER_109_127 ();
 DECAPx1_ASAP7_75t_R FILLER_109_137 ();
 FILLER_ASAP7_75t_R FILLER_109_151 ();
 DECAPx1_ASAP7_75t_R FILLER_109_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_189 ();
 DECAPx6_ASAP7_75t_R FILLER_109_216 ();
 DECAPx2_ASAP7_75t_R FILLER_109_230 ();
 DECAPx10_ASAP7_75t_R FILLER_109_239 ();
 DECAPx1_ASAP7_75t_R FILLER_109_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_265 ();
 FILLER_ASAP7_75t_R FILLER_109_272 ();
 DECAPx10_ASAP7_75t_R FILLER_109_311 ();
 DECAPx10_ASAP7_75t_R FILLER_109_333 ();
 DECAPx10_ASAP7_75t_R FILLER_109_355 ();
 DECAPx10_ASAP7_75t_R FILLER_109_377 ();
 DECAPx10_ASAP7_75t_R FILLER_109_399 ();
 DECAPx1_ASAP7_75t_R FILLER_109_421 ();
 DECAPx1_ASAP7_75t_R FILLER_109_428 ();
 DECAPx2_ASAP7_75t_R FILLER_109_435 ();
 FILLER_ASAP7_75t_R FILLER_109_441 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_472 ();
 FILLER_ASAP7_75t_R FILLER_109_481 ();
 DECAPx1_ASAP7_75t_R FILLER_109_491 ();
 DECAPx4_ASAP7_75t_R FILLER_109_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_511 ();
 FILLER_ASAP7_75t_R FILLER_109_520 ();
 DECAPx2_ASAP7_75t_R FILLER_109_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_587 ();
 FILLER_ASAP7_75t_R FILLER_109_614 ();
 DECAPx4_ASAP7_75t_R FILLER_109_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_640 ();
 DECAPx4_ASAP7_75t_R FILLER_109_647 ();
 FILLER_ASAP7_75t_R FILLER_109_657 ();
 DECAPx2_ASAP7_75t_R FILLER_109_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_697 ();
 DECAPx2_ASAP7_75t_R FILLER_109_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_730 ();
 DECAPx1_ASAP7_75t_R FILLER_109_745 ();
 FILLER_ASAP7_75t_R FILLER_109_756 ();
 DECAPx10_ASAP7_75t_R FILLER_109_767 ();
 DECAPx10_ASAP7_75t_R FILLER_109_789 ();
 DECAPx6_ASAP7_75t_R FILLER_109_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_825 ();
 DECAPx10_ASAP7_75t_R FILLER_109_831 ();
 DECAPx4_ASAP7_75t_R FILLER_109_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_109_863 ();
 DECAPx1_ASAP7_75t_R FILLER_109_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_109_924 ();
 FILLER_ASAP7_75t_R FILLER_109_927 ();
 DECAPx10_ASAP7_75t_R FILLER_110_2 ();
 DECAPx10_ASAP7_75t_R FILLER_110_24 ();
 DECAPx10_ASAP7_75t_R FILLER_110_46 ();
 DECAPx1_ASAP7_75t_R FILLER_110_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_85 ();
 DECAPx10_ASAP7_75t_R FILLER_110_98 ();
 DECAPx6_ASAP7_75t_R FILLER_110_120 ();
 FILLER_ASAP7_75t_R FILLER_110_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_142 ();
 DECAPx1_ASAP7_75t_R FILLER_110_159 ();
 DECAPx1_ASAP7_75t_R FILLER_110_169 ();
 DECAPx1_ASAP7_75t_R FILLER_110_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_180 ();
 FILLER_ASAP7_75t_R FILLER_110_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_194 ();
 DECAPx6_ASAP7_75t_R FILLER_110_222 ();
 FILLER_ASAP7_75t_R FILLER_110_236 ();
 DECAPx1_ASAP7_75t_R FILLER_110_244 ();
 DECAPx10_ASAP7_75t_R FILLER_110_254 ();
 DECAPx2_ASAP7_75t_R FILLER_110_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_282 ();
 FILLER_ASAP7_75t_R FILLER_110_289 ();
 DECAPx1_ASAP7_75t_R FILLER_110_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_298 ();
 DECAPx10_ASAP7_75t_R FILLER_110_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_324 ();
 DECAPx1_ASAP7_75t_R FILLER_110_331 ();
 DECAPx1_ASAP7_75t_R FILLER_110_349 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_365 ();
 DECAPx4_ASAP7_75t_R FILLER_110_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_392 ();
 DECAPx1_ASAP7_75t_R FILLER_110_399 ();
 DECAPx6_ASAP7_75t_R FILLER_110_409 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_432 ();
 DECAPx1_ASAP7_75t_R FILLER_110_447 ();
 DECAPx2_ASAP7_75t_R FILLER_110_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_484 ();
 DECAPx4_ASAP7_75t_R FILLER_110_496 ();
 DECAPx2_ASAP7_75t_R FILLER_110_512 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_524 ();
 FILLER_ASAP7_75t_R FILLER_110_535 ();
 DECAPx2_ASAP7_75t_R FILLER_110_540 ();
 FILLER_ASAP7_75t_R FILLER_110_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_554 ();
 DECAPx2_ASAP7_75t_R FILLER_110_560 ();
 DECAPx1_ASAP7_75t_R FILLER_110_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_583 ();
 DECAPx2_ASAP7_75t_R FILLER_110_590 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_110_596 ();
 DECAPx6_ASAP7_75t_R FILLER_110_623 ();
 DECAPx2_ASAP7_75t_R FILLER_110_653 ();
 FILLER_ASAP7_75t_R FILLER_110_659 ();
 DECAPx6_ASAP7_75t_R FILLER_110_667 ();
 DECAPx1_ASAP7_75t_R FILLER_110_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_685 ();
 DECAPx1_ASAP7_75t_R FILLER_110_693 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_697 ();
 DECAPx6_ASAP7_75t_R FILLER_110_712 ();
 DECAPx2_ASAP7_75t_R FILLER_110_726 ();
 DECAPx2_ASAP7_75t_R FILLER_110_739 ();
 DECAPx10_ASAP7_75t_R FILLER_110_771 ();
 DECAPx1_ASAP7_75t_R FILLER_110_793 ();
 DECAPx6_ASAP7_75t_R FILLER_110_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_818 ();
 DECAPx1_ASAP7_75t_R FILLER_110_834 ();
 DECAPx10_ASAP7_75t_R FILLER_110_844 ();
 DECAPx6_ASAP7_75t_R FILLER_110_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_110_906 ();
 FILLER_ASAP7_75t_R FILLER_110_922 ();
 DECAPx10_ASAP7_75t_R FILLER_111_2 ();
 DECAPx10_ASAP7_75t_R FILLER_111_24 ();
 DECAPx10_ASAP7_75t_R FILLER_111_46 ();
 DECAPx6_ASAP7_75t_R FILLER_111_68 ();
 FILLER_ASAP7_75t_R FILLER_111_82 ();
 DECAPx6_ASAP7_75t_R FILLER_111_87 ();
 DECAPx2_ASAP7_75t_R FILLER_111_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_107 ();
 DECAPx6_ASAP7_75t_R FILLER_111_111 ();
 DECAPx4_ASAP7_75t_R FILLER_111_139 ();
 DECAPx4_ASAP7_75t_R FILLER_111_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_165 ();
 FILLER_ASAP7_75t_R FILLER_111_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_228 ();
 DECAPx10_ASAP7_75t_R FILLER_111_258 ();
 DECAPx10_ASAP7_75t_R FILLER_111_280 ();
 DECAPx4_ASAP7_75t_R FILLER_111_302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_365 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_392 ();
 DECAPx2_ASAP7_75t_R FILLER_111_418 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_432 ();
 DECAPx6_ASAP7_75t_R FILLER_111_443 ();
 DECAPx10_ASAP7_75t_R FILLER_111_483 ();
 DECAPx2_ASAP7_75t_R FILLER_111_505 ();
 DECAPx10_ASAP7_75t_R FILLER_111_522 ();
 DECAPx6_ASAP7_75t_R FILLER_111_544 ();
 DECAPx2_ASAP7_75t_R FILLER_111_558 ();
 DECAPx10_ASAP7_75t_R FILLER_111_578 ();
 DECAPx10_ASAP7_75t_R FILLER_111_600 ();
 DECAPx2_ASAP7_75t_R FILLER_111_622 ();
 FILLER_ASAP7_75t_R FILLER_111_628 ();
 DECAPx2_ASAP7_75t_R FILLER_111_646 ();
 DECAPx6_ASAP7_75t_R FILLER_111_662 ();
 DECAPx1_ASAP7_75t_R FILLER_111_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_691 ();
 DECAPx4_ASAP7_75t_R FILLER_111_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_716 ();
 DECAPx1_ASAP7_75t_R FILLER_111_725 ();
 DECAPx6_ASAP7_75t_R FILLER_111_739 ();
 DECAPx1_ASAP7_75t_R FILLER_111_753 ();
 DECAPx10_ASAP7_75t_R FILLER_111_767 ();
 DECAPx1_ASAP7_75t_R FILLER_111_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_111_845 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_111_868 ();
 FILLER_ASAP7_75t_R FILLER_111_927 ();
 DECAPx10_ASAP7_75t_R FILLER_112_2 ();
 DECAPx10_ASAP7_75t_R FILLER_112_24 ();
 DECAPx10_ASAP7_75t_R FILLER_112_46 ();
 DECAPx10_ASAP7_75t_R FILLER_112_68 ();
 DECAPx2_ASAP7_75t_R FILLER_112_90 ();
 DECAPx10_ASAP7_75t_R FILLER_112_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_160 ();
 DECAPx2_ASAP7_75t_R FILLER_112_189 ();
 FILLER_ASAP7_75t_R FILLER_112_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_219 ();
 DECAPx6_ASAP7_75t_R FILLER_112_249 ();
 DECAPx2_ASAP7_75t_R FILLER_112_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_269 ();
 DECAPx4_ASAP7_75t_R FILLER_112_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_293 ();
 DECAPx4_ASAP7_75t_R FILLER_112_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_310 ();
 DECAPx1_ASAP7_75t_R FILLER_112_317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_327 ();
 DECAPx2_ASAP7_75t_R FILLER_112_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_355 ();
 DECAPx2_ASAP7_75t_R FILLER_112_364 ();
 DECAPx10_ASAP7_75t_R FILLER_112_440 ();
 DECAPx2_ASAP7_75t_R FILLER_112_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_470 ();
 DECAPx4_ASAP7_75t_R FILLER_112_482 ();
 DECAPx1_ASAP7_75t_R FILLER_112_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_504 ();
 DECAPx2_ASAP7_75t_R FILLER_112_531 ();
 FILLER_ASAP7_75t_R FILLER_112_537 ();
 DECAPx10_ASAP7_75t_R FILLER_112_547 ();
 DECAPx10_ASAP7_75t_R FILLER_112_569 ();
 DECAPx10_ASAP7_75t_R FILLER_112_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_112_613 ();
 FILLER_ASAP7_75t_R FILLER_112_635 ();
 DECAPx6_ASAP7_75t_R FILLER_112_651 ();
 FILLER_ASAP7_75t_R FILLER_112_671 ();
 DECAPx6_ASAP7_75t_R FILLER_112_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_700 ();
 DECAPx4_ASAP7_75t_R FILLER_112_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_747 ();
 DECAPx2_ASAP7_75t_R FILLER_112_754 ();
 FILLER_ASAP7_75t_R FILLER_112_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_781 ();
 DECAPx2_ASAP7_75t_R FILLER_112_794 ();
 FILLER_ASAP7_75t_R FILLER_112_800 ();
 DECAPx2_ASAP7_75t_R FILLER_112_811 ();
 FILLER_ASAP7_75t_R FILLER_112_817 ();
 FILLER_ASAP7_75t_R FILLER_112_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_112_899 ();
 DECAPx10_ASAP7_75t_R FILLER_113_2 ();
 DECAPx10_ASAP7_75t_R FILLER_113_24 ();
 DECAPx10_ASAP7_75t_R FILLER_113_46 ();
 DECAPx10_ASAP7_75t_R FILLER_113_68 ();
 FILLER_ASAP7_75t_R FILLER_113_90 ();
 FILLER_ASAP7_75t_R FILLER_113_126 ();
 DECAPx2_ASAP7_75t_R FILLER_113_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_140 ();
 DECAPx10_ASAP7_75t_R FILLER_113_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_177 ();
 DECAPx10_ASAP7_75t_R FILLER_113_181 ();
 DECAPx6_ASAP7_75t_R FILLER_113_240 ();
 FILLER_ASAP7_75t_R FILLER_113_254 ();
 FILLER_ASAP7_75t_R FILLER_113_282 ();
 DECAPx6_ASAP7_75t_R FILLER_113_322 ();
 FILLER_ASAP7_75t_R FILLER_113_336 ();
 DECAPx10_ASAP7_75t_R FILLER_113_341 ();
 DECAPx6_ASAP7_75t_R FILLER_113_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_401 ();
 DECAPx6_ASAP7_75t_R FILLER_113_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_422 ();
 DECAPx6_ASAP7_75t_R FILLER_113_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_446 ();
 DECAPx6_ASAP7_75t_R FILLER_113_461 ();
 DECAPx2_ASAP7_75t_R FILLER_113_475 ();
 DECAPx6_ASAP7_75t_R FILLER_113_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_561 ();
 DECAPx2_ASAP7_75t_R FILLER_113_568 ();
 FILLER_ASAP7_75t_R FILLER_113_586 ();
 DECAPx1_ASAP7_75t_R FILLER_113_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_604 ();
 DECAPx10_ASAP7_75t_R FILLER_113_611 ();
 DECAPx10_ASAP7_75t_R FILLER_113_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_655 ();
 DECAPx1_ASAP7_75t_R FILLER_113_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_667 ();
 DECAPx6_ASAP7_75t_R FILLER_113_675 ();
 DECAPx2_ASAP7_75t_R FILLER_113_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_723 ();
 DECAPx2_ASAP7_75t_R FILLER_113_742 ();
 DECAPx6_ASAP7_75t_R FILLER_113_815 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_113_829 ();
 FILLER_ASAP7_75t_R FILLER_113_835 ();
 FILLER_ASAP7_75t_R FILLER_113_863 ();
 FILLER_ASAP7_75t_R FILLER_113_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_113_924 ();
 FILLER_ASAP7_75t_R FILLER_113_927 ();
 DECAPx10_ASAP7_75t_R FILLER_114_2 ();
 DECAPx10_ASAP7_75t_R FILLER_114_24 ();
 DECAPx10_ASAP7_75t_R FILLER_114_46 ();
 DECAPx6_ASAP7_75t_R FILLER_114_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_111 ();
 DECAPx1_ASAP7_75t_R FILLER_114_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_137 ();
 FILLER_ASAP7_75t_R FILLER_114_150 ();
 DECAPx10_ASAP7_75t_R FILLER_114_166 ();
 DECAPx10_ASAP7_75t_R FILLER_114_188 ();
 DECAPx10_ASAP7_75t_R FILLER_114_213 ();
 DECAPx4_ASAP7_75t_R FILLER_114_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_245 ();
 FILLER_ASAP7_75t_R FILLER_114_266 ();
 DECAPx2_ASAP7_75t_R FILLER_114_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_289 ();
 FILLER_ASAP7_75t_R FILLER_114_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_310 ();
 DECAPx2_ASAP7_75t_R FILLER_114_317 ();
 FILLER_ASAP7_75t_R FILLER_114_323 ();
 DECAPx10_ASAP7_75t_R FILLER_114_359 ();
 DECAPx2_ASAP7_75t_R FILLER_114_381 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_387 ();
 DECAPx10_ASAP7_75t_R FILLER_114_393 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_415 ();
 DECAPx1_ASAP7_75t_R FILLER_114_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_433 ();
 DECAPx2_ASAP7_75t_R FILLER_114_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_476 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_491 ();
 FILLER_ASAP7_75t_R FILLER_114_503 ();
 DECAPx6_ASAP7_75t_R FILLER_114_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_552 ();
 FILLER_ASAP7_75t_R FILLER_114_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_611 ();
 DECAPx10_ASAP7_75t_R FILLER_114_620 ();
 DECAPx1_ASAP7_75t_R FILLER_114_642 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_653 ();
 DECAPx6_ASAP7_75t_R FILLER_114_662 ();
 DECAPx1_ASAP7_75t_R FILLER_114_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_680 ();
 DECAPx10_ASAP7_75t_R FILLER_114_687 ();
 DECAPx2_ASAP7_75t_R FILLER_114_709 ();
 FILLER_ASAP7_75t_R FILLER_114_715 ();
 DECAPx6_ASAP7_75t_R FILLER_114_723 ();
 DECAPx10_ASAP7_75t_R FILLER_114_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_765 ();
 FILLER_ASAP7_75t_R FILLER_114_775 ();
 DECAPx4_ASAP7_75t_R FILLER_114_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_806 ();
 DECAPx1_ASAP7_75t_R FILLER_114_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_820 ();
 DECAPx2_ASAP7_75t_R FILLER_114_827 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_114_833 ();
 DECAPx2_ASAP7_75t_R FILLER_114_839 ();
 FILLER_ASAP7_75t_R FILLER_114_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_114_907 ();
 DECAPx10_ASAP7_75t_R FILLER_115_2 ();
 DECAPx10_ASAP7_75t_R FILLER_115_24 ();
 DECAPx10_ASAP7_75t_R FILLER_115_46 ();
 DECAPx6_ASAP7_75t_R FILLER_115_68 ();
 DECAPx1_ASAP7_75t_R FILLER_115_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_86 ();
 DECAPx4_ASAP7_75t_R FILLER_115_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_126 ();
 DECAPx1_ASAP7_75t_R FILLER_115_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_159 ();
 DECAPx1_ASAP7_75t_R FILLER_115_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_172 ();
 DECAPx10_ASAP7_75t_R FILLER_115_188 ();
 DECAPx6_ASAP7_75t_R FILLER_115_210 ();
 DECAPx6_ASAP7_75t_R FILLER_115_236 ();
 DECAPx1_ASAP7_75t_R FILLER_115_250 ();
 DECAPx1_ASAP7_75t_R FILLER_115_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_316 ();
 DECAPx1_ASAP7_75t_R FILLER_115_343 ();
 DECAPx10_ASAP7_75t_R FILLER_115_376 ();
 DECAPx10_ASAP7_75t_R FILLER_115_398 ();
 DECAPx10_ASAP7_75t_R FILLER_115_420 ();
 DECAPx2_ASAP7_75t_R FILLER_115_442 ();
 DECAPx2_ASAP7_75t_R FILLER_115_460 ();
 DECAPx10_ASAP7_75t_R FILLER_115_492 ();
 DECAPx1_ASAP7_75t_R FILLER_115_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_518 ();
 DECAPx1_ASAP7_75t_R FILLER_115_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_534 ();
 DECAPx2_ASAP7_75t_R FILLER_115_549 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_555 ();
 DECAPx2_ASAP7_75t_R FILLER_115_564 ();
 DECAPx2_ASAP7_75t_R FILLER_115_576 ();
 DECAPx10_ASAP7_75t_R FILLER_115_588 ();
 DECAPx4_ASAP7_75t_R FILLER_115_610 ();
 FILLER_ASAP7_75t_R FILLER_115_620 ();
 DECAPx2_ASAP7_75t_R FILLER_115_634 ();
 FILLER_ASAP7_75t_R FILLER_115_640 ();
 DECAPx10_ASAP7_75t_R FILLER_115_694 ();
 FILLER_ASAP7_75t_R FILLER_115_716 ();
 FILLER_ASAP7_75t_R FILLER_115_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_115_752 ();
 DECAPx10_ASAP7_75t_R FILLER_115_758 ();
 DECAPx10_ASAP7_75t_R FILLER_115_780 ();
 DECAPx1_ASAP7_75t_R FILLER_115_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_115_806 ();
 DECAPx6_ASAP7_75t_R FILLER_115_833 ();
 DECAPx1_ASAP7_75t_R FILLER_115_847 ();
 FILLER_ASAP7_75t_R FILLER_115_927 ();
 DECAPx10_ASAP7_75t_R FILLER_116_2 ();
 DECAPx10_ASAP7_75t_R FILLER_116_24 ();
 DECAPx10_ASAP7_75t_R FILLER_116_46 ();
 DECAPx10_ASAP7_75t_R FILLER_116_68 ();
 DECAPx10_ASAP7_75t_R FILLER_116_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_112 ();
 FILLER_ASAP7_75t_R FILLER_116_119 ();
 DECAPx1_ASAP7_75t_R FILLER_116_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_155 ();
 DECAPx2_ASAP7_75t_R FILLER_116_164 ();
 DECAPx4_ASAP7_75t_R FILLER_116_199 ();
 DECAPx2_ASAP7_75t_R FILLER_116_215 ();
 DECAPx2_ASAP7_75t_R FILLER_116_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_253 ();
 DECAPx2_ASAP7_75t_R FILLER_116_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_268 ();
 DECAPx10_ASAP7_75t_R FILLER_116_272 ();
 DECAPx2_ASAP7_75t_R FILLER_116_294 ();
 DECAPx4_ASAP7_75t_R FILLER_116_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_319 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_328 ();
 DECAPx6_ASAP7_75t_R FILLER_116_334 ();
 DECAPx1_ASAP7_75t_R FILLER_116_348 ();
 DECAPx1_ASAP7_75t_R FILLER_116_358 ();
 DECAPx2_ASAP7_75t_R FILLER_116_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_378 ();
 DECAPx2_ASAP7_75t_R FILLER_116_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_391 ();
 DECAPx2_ASAP7_75t_R FILLER_116_395 ();
 FILLER_ASAP7_75t_R FILLER_116_401 ();
 DECAPx1_ASAP7_75t_R FILLER_116_409 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_425 ();
 DECAPx10_ASAP7_75t_R FILLER_116_431 ();
 DECAPx2_ASAP7_75t_R FILLER_116_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_459 ();
 DECAPx6_ASAP7_75t_R FILLER_116_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_478 ();
 DECAPx10_ASAP7_75t_R FILLER_116_484 ();
 DECAPx4_ASAP7_75t_R FILLER_116_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_516 ();
 DECAPx6_ASAP7_75t_R FILLER_116_523 ();
 DECAPx2_ASAP7_75t_R FILLER_116_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_543 ();
 DECAPx1_ASAP7_75t_R FILLER_116_547 ();
 DECAPx10_ASAP7_75t_R FILLER_116_569 ();
 DECAPx6_ASAP7_75t_R FILLER_116_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_645 ();
 FILLER_ASAP7_75t_R FILLER_116_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_670 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_679 ();
 DECAPx2_ASAP7_75t_R FILLER_116_685 ();
 FILLER_ASAP7_75t_R FILLER_116_691 ();
 DECAPx10_ASAP7_75t_R FILLER_116_704 ();
 DECAPx4_ASAP7_75t_R FILLER_116_726 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_736 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_760 ();
 DECAPx6_ASAP7_75t_R FILLER_116_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_791 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_116_807 ();
 DECAPx1_ASAP7_75t_R FILLER_116_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_116_829 ();
 DECAPx1_ASAP7_75t_R FILLER_116_833 ();
 DECAPx10_ASAP7_75t_R FILLER_117_2 ();
 DECAPx10_ASAP7_75t_R FILLER_117_24 ();
 DECAPx10_ASAP7_75t_R FILLER_117_46 ();
 DECAPx10_ASAP7_75t_R FILLER_117_68 ();
 DECAPx6_ASAP7_75t_R FILLER_117_90 ();
 DECAPx2_ASAP7_75t_R FILLER_117_104 ();
 DECAPx10_ASAP7_75t_R FILLER_117_136 ();
 DECAPx4_ASAP7_75t_R FILLER_117_158 ();
 FILLER_ASAP7_75t_R FILLER_117_168 ();
 FILLER_ASAP7_75t_R FILLER_117_176 ();
 DECAPx2_ASAP7_75t_R FILLER_117_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_190 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_213 ();
 DECAPx4_ASAP7_75t_R FILLER_117_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_232 ();
 DECAPx1_ASAP7_75t_R FILLER_117_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_242 ();
 DECAPx10_ASAP7_75t_R FILLER_117_246 ();
 DECAPx10_ASAP7_75t_R FILLER_117_268 ();
 DECAPx10_ASAP7_75t_R FILLER_117_290 ();
 DECAPx2_ASAP7_75t_R FILLER_117_312 ();
 DECAPx10_ASAP7_75t_R FILLER_117_344 ();
 DECAPx1_ASAP7_75t_R FILLER_117_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_402 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_410 ();
 DECAPx6_ASAP7_75t_R FILLER_117_442 ();
 DECAPx2_ASAP7_75t_R FILLER_117_456 ();
 DECAPx10_ASAP7_75t_R FILLER_117_470 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_492 ();
 DECAPx1_ASAP7_75t_R FILLER_117_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_574 ();
 DECAPx6_ASAP7_75t_R FILLER_117_583 ();
 FILLER_ASAP7_75t_R FILLER_117_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_629 ();
 DECAPx10_ASAP7_75t_R FILLER_117_662 ();
 FILLER_ASAP7_75t_R FILLER_117_684 ();
 DECAPx2_ASAP7_75t_R FILLER_117_712 ();
 FILLER_ASAP7_75t_R FILLER_117_718 ();
 DECAPx2_ASAP7_75t_R FILLER_117_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_742 ();
 DECAPx2_ASAP7_75t_R FILLER_117_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_787 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_117_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_117_911 ();
 FILLER_ASAP7_75t_R FILLER_117_927 ();
 DECAPx10_ASAP7_75t_R FILLER_118_2 ();
 DECAPx10_ASAP7_75t_R FILLER_118_24 ();
 DECAPx10_ASAP7_75t_R FILLER_118_46 ();
 DECAPx6_ASAP7_75t_R FILLER_118_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_89 ();
 DECAPx1_ASAP7_75t_R FILLER_118_96 ();
 DECAPx4_ASAP7_75t_R FILLER_118_103 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_122 ();
 DECAPx10_ASAP7_75t_R FILLER_118_128 ();
 DECAPx6_ASAP7_75t_R FILLER_118_150 ();
 FILLER_ASAP7_75t_R FILLER_118_164 ();
 DECAPx2_ASAP7_75t_R FILLER_118_226 ();
 FILLER_ASAP7_75t_R FILLER_118_232 ();
 DECAPx6_ASAP7_75t_R FILLER_118_260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_274 ();
 DECAPx6_ASAP7_75t_R FILLER_118_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_294 ();
 DECAPx6_ASAP7_75t_R FILLER_118_304 ();
 DECAPx1_ASAP7_75t_R FILLER_118_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_337 ();
 DECAPx4_ASAP7_75t_R FILLER_118_344 ();
 FILLER_ASAP7_75t_R FILLER_118_354 ();
 DECAPx2_ASAP7_75t_R FILLER_118_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_388 ();
 DECAPx1_ASAP7_75t_R FILLER_118_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_400 ();
 DECAPx1_ASAP7_75t_R FILLER_118_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_461 ();
 DECAPx2_ASAP7_75t_R FILLER_118_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_476 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_483 ();
 DECAPx4_ASAP7_75t_R FILLER_118_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_530 ();
 DECAPx1_ASAP7_75t_R FILLER_118_537 ();
 DECAPx6_ASAP7_75t_R FILLER_118_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_558 ();
 DECAPx4_ASAP7_75t_R FILLER_118_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_583 ();
 DECAPx4_ASAP7_75t_R FILLER_118_595 ();
 FILLER_ASAP7_75t_R FILLER_118_605 ();
 DECAPx6_ASAP7_75t_R FILLER_118_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_636 ();
 DECAPx2_ASAP7_75t_R FILLER_118_643 ();
 FILLER_ASAP7_75t_R FILLER_118_649 ();
 DECAPx2_ASAP7_75t_R FILLER_118_654 ();
 FILLER_ASAP7_75t_R FILLER_118_660 ();
 DECAPx2_ASAP7_75t_R FILLER_118_674 ();
 FILLER_ASAP7_75t_R FILLER_118_680 ();
 DECAPx4_ASAP7_75t_R FILLER_118_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_713 ();
 DECAPx6_ASAP7_75t_R FILLER_118_725 ();
 DECAPx1_ASAP7_75t_R FILLER_118_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_743 ();
 DECAPx4_ASAP7_75t_R FILLER_118_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_118_783 ();
 DECAPx2_ASAP7_75t_R FILLER_118_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_827 ();
 FILLER_ASAP7_75t_R FILLER_118_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_118_864 ();
 FILLER_ASAP7_75t_R FILLER_118_872 ();
 DECAPx10_ASAP7_75t_R FILLER_119_2 ();
 DECAPx10_ASAP7_75t_R FILLER_119_24 ();
 DECAPx10_ASAP7_75t_R FILLER_119_46 ();
 DECAPx4_ASAP7_75t_R FILLER_119_68 ();
 DECAPx2_ASAP7_75t_R FILLER_119_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_129 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_145 ();
 DECAPx6_ASAP7_75t_R FILLER_119_161 ();
 DECAPx2_ASAP7_75t_R FILLER_119_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_181 ();
 DECAPx6_ASAP7_75t_R FILLER_119_185 ();
 FILLER_ASAP7_75t_R FILLER_119_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_210 ();
 DECAPx2_ASAP7_75t_R FILLER_119_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_252 ();
 FILLER_ASAP7_75t_R FILLER_119_279 ();
 DECAPx6_ASAP7_75t_R FILLER_119_316 ();
 DECAPx1_ASAP7_75t_R FILLER_119_330 ();
 DECAPx4_ASAP7_75t_R FILLER_119_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_384 ();
 DECAPx1_ASAP7_75t_R FILLER_119_388 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_426 ();
 DECAPx4_ASAP7_75t_R FILLER_119_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_443 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_463 ();
 DECAPx1_ASAP7_75t_R FILLER_119_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_500 ();
 DECAPx2_ASAP7_75t_R FILLER_119_516 ();
 FILLER_ASAP7_75t_R FILLER_119_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_550 ();
 DECAPx4_ASAP7_75t_R FILLER_119_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_567 ();
 DECAPx2_ASAP7_75t_R FILLER_119_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_593 ();
 DECAPx2_ASAP7_75t_R FILLER_119_626 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_632 ();
 DECAPx10_ASAP7_75t_R FILLER_119_638 ();
 DECAPx4_ASAP7_75t_R FILLER_119_660 ();
 DECAPx2_ASAP7_75t_R FILLER_119_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_692 ();
 DECAPx2_ASAP7_75t_R FILLER_119_699 ();
 DECAPx2_ASAP7_75t_R FILLER_119_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_119_728 ();
 DECAPx2_ASAP7_75t_R FILLER_119_750 ();
 FILLER_ASAP7_75t_R FILLER_119_756 ();
 DECAPx6_ASAP7_75t_R FILLER_119_761 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_775 ();
 DECAPx6_ASAP7_75t_R FILLER_119_792 ();
 DECAPx10_ASAP7_75t_R FILLER_119_816 ();
 DECAPx4_ASAP7_75t_R FILLER_119_838 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_119_848 ();
 FILLER_ASAP7_75t_R FILLER_119_927 ();
 DECAPx10_ASAP7_75t_R FILLER_120_2 ();
 DECAPx10_ASAP7_75t_R FILLER_120_24 ();
 DECAPx10_ASAP7_75t_R FILLER_120_46 ();
 DECAPx4_ASAP7_75t_R FILLER_120_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_78 ();
 FILLER_ASAP7_75t_R FILLER_120_113 ();
 DECAPx10_ASAP7_75t_R FILLER_120_177 ();
 DECAPx10_ASAP7_75t_R FILLER_120_199 ();
 DECAPx2_ASAP7_75t_R FILLER_120_221 ();
 FILLER_ASAP7_75t_R FILLER_120_227 ();
 DECAPx2_ASAP7_75t_R FILLER_120_235 ();
 FILLER_ASAP7_75t_R FILLER_120_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_254 ();
 DECAPx2_ASAP7_75t_R FILLER_120_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_322 ();
 DECAPx1_ASAP7_75t_R FILLER_120_329 ();
 DECAPx1_ASAP7_75t_R FILLER_120_361 ();
 DECAPx10_ASAP7_75t_R FILLER_120_372 ();
 DECAPx10_ASAP7_75t_R FILLER_120_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_425 ();
 FILLER_ASAP7_75t_R FILLER_120_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_467 ();
 DECAPx6_ASAP7_75t_R FILLER_120_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_488 ();
 DECAPx10_ASAP7_75t_R FILLER_120_499 ();
 DECAPx2_ASAP7_75t_R FILLER_120_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_527 ();
 DECAPx1_ASAP7_75t_R FILLER_120_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_546 ();
 DECAPx10_ASAP7_75t_R FILLER_120_553 ();
 DECAPx2_ASAP7_75t_R FILLER_120_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_588 ();
 DECAPx10_ASAP7_75t_R FILLER_120_605 ();
 DECAPx6_ASAP7_75t_R FILLER_120_627 ();
 DECAPx2_ASAP7_75t_R FILLER_120_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_647 ();
 DECAPx1_ASAP7_75t_R FILLER_120_654 ();
 DECAPx2_ASAP7_75t_R FILLER_120_661 ();
 DECAPx1_ASAP7_75t_R FILLER_120_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_696 ();
 DECAPx1_ASAP7_75t_R FILLER_120_715 ();
 FILLER_ASAP7_75t_R FILLER_120_727 ();
 DECAPx2_ASAP7_75t_R FILLER_120_734 ();
 FILLER_ASAP7_75t_R FILLER_120_740 ();
 DECAPx4_ASAP7_75t_R FILLER_120_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_120_766 ();
 DECAPx4_ASAP7_75t_R FILLER_120_795 ();
 FILLER_ASAP7_75t_R FILLER_120_805 ();
 DECAPx6_ASAP7_75t_R FILLER_120_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_833 ();
 DECAPx6_ASAP7_75t_R FILLER_120_841 ();
 DECAPx2_ASAP7_75t_R FILLER_120_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_120_904 ();
 DECAPx10_ASAP7_75t_R FILLER_121_2 ();
 DECAPx10_ASAP7_75t_R FILLER_121_24 ();
 DECAPx10_ASAP7_75t_R FILLER_121_46 ();
 DECAPx6_ASAP7_75t_R FILLER_121_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_82 ();
 FILLER_ASAP7_75t_R FILLER_121_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_118 ();
 DECAPx1_ASAP7_75t_R FILLER_121_125 ();
 FILLER_ASAP7_75t_R FILLER_121_137 ();
 FILLER_ASAP7_75t_R FILLER_121_150 ();
 DECAPx4_ASAP7_75t_R FILLER_121_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_181 ();
 DECAPx4_ASAP7_75t_R FILLER_121_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_206 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_210 ();
 DECAPx1_ASAP7_75t_R FILLER_121_221 ();
 DECAPx6_ASAP7_75t_R FILLER_121_237 ();
 DECAPx1_ASAP7_75t_R FILLER_121_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_271 ();
 DECAPx1_ASAP7_75t_R FILLER_121_288 ();
 DECAPx2_ASAP7_75t_R FILLER_121_312 ();
 FILLER_ASAP7_75t_R FILLER_121_347 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_359 ();
 DECAPx1_ASAP7_75t_R FILLER_121_388 ();
 DECAPx1_ASAP7_75t_R FILLER_121_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_403 ();
 DECAPx1_ASAP7_75t_R FILLER_121_407 ();
 DECAPx2_ASAP7_75t_R FILLER_121_419 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_425 ();
 DECAPx10_ASAP7_75t_R FILLER_121_465 ();
 DECAPx1_ASAP7_75t_R FILLER_121_487 ();
 DECAPx10_ASAP7_75t_R FILLER_121_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_519 ();
 DECAPx10_ASAP7_75t_R FILLER_121_528 ();
 DECAPx10_ASAP7_75t_R FILLER_121_550 ();
 DECAPx2_ASAP7_75t_R FILLER_121_572 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_578 ();
 DECAPx10_ASAP7_75t_R FILLER_121_594 ();
 DECAPx2_ASAP7_75t_R FILLER_121_616 ();
 DECAPx4_ASAP7_75t_R FILLER_121_630 ();
 DECAPx2_ASAP7_75t_R FILLER_121_669 ();
 FILLER_ASAP7_75t_R FILLER_121_675 ();
 DECAPx10_ASAP7_75t_R FILLER_121_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_711 ();
 DECAPx2_ASAP7_75t_R FILLER_121_718 ();
 FILLER_ASAP7_75t_R FILLER_121_724 ();
 FILLER_ASAP7_75t_R FILLER_121_741 ();
 DECAPx2_ASAP7_75t_R FILLER_121_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_759 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_777 ();
 DECAPx2_ASAP7_75t_R FILLER_121_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_796 ();
 DECAPx6_ASAP7_75t_R FILLER_121_802 ();
 DECAPx1_ASAP7_75t_R FILLER_121_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_820 ();
 DECAPx2_ASAP7_75t_R FILLER_121_857 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_121_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_121_933 ();
 DECAPx10_ASAP7_75t_R FILLER_122_2 ();
 DECAPx10_ASAP7_75t_R FILLER_122_24 ();
 DECAPx10_ASAP7_75t_R FILLER_122_46 ();
 DECAPx10_ASAP7_75t_R FILLER_122_68 ();
 DECAPx10_ASAP7_75t_R FILLER_122_90 ();
 DECAPx10_ASAP7_75t_R FILLER_122_112 ();
 DECAPx6_ASAP7_75t_R FILLER_122_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_160 ();
 DECAPx1_ASAP7_75t_R FILLER_122_167 ();
 DECAPx1_ASAP7_75t_R FILLER_122_183 ();
 FILLER_ASAP7_75t_R FILLER_122_209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_219 ();
 DECAPx6_ASAP7_75t_R FILLER_122_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_265 ();
 DECAPx2_ASAP7_75t_R FILLER_122_271 ();
 FILLER_ASAP7_75t_R FILLER_122_277 ();
 DECAPx4_ASAP7_75t_R FILLER_122_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_328 ();
 DECAPx10_ASAP7_75t_R FILLER_122_338 ();
 DECAPx1_ASAP7_75t_R FILLER_122_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_364 ();
 DECAPx1_ASAP7_75t_R FILLER_122_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_388 ();
 DECAPx4_ASAP7_75t_R FILLER_122_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_428 ();
 DECAPx6_ASAP7_75t_R FILLER_122_444 ();
 DECAPx1_ASAP7_75t_R FILLER_122_458 ();
 DECAPx4_ASAP7_75t_R FILLER_122_464 ();
 FILLER_ASAP7_75t_R FILLER_122_474 ();
 DECAPx6_ASAP7_75t_R FILLER_122_490 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_122_504 ();
 DECAPx2_ASAP7_75t_R FILLER_122_515 ();
 DECAPx4_ASAP7_75t_R FILLER_122_530 ();
 FILLER_ASAP7_75t_R FILLER_122_540 ();
 DECAPx2_ASAP7_75t_R FILLER_122_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_563 ();
 DECAPx1_ASAP7_75t_R FILLER_122_571 ();
 FILLER_ASAP7_75t_R FILLER_122_581 ();
 DECAPx6_ASAP7_75t_R FILLER_122_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_605 ();
 DECAPx10_ASAP7_75t_R FILLER_122_656 ();
 DECAPx6_ASAP7_75t_R FILLER_122_678 ();
 DECAPx1_ASAP7_75t_R FILLER_122_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_696 ();
 DECAPx6_ASAP7_75t_R FILLER_122_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_718 ();
 DECAPx6_ASAP7_75t_R FILLER_122_725 ();
 DECAPx2_ASAP7_75t_R FILLER_122_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_745 ();
 DECAPx10_ASAP7_75t_R FILLER_122_772 ();
 DECAPx2_ASAP7_75t_R FILLER_122_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_828 ();
 DECAPx2_ASAP7_75t_R FILLER_122_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_122_933 ();
 DECAPx10_ASAP7_75t_R FILLER_123_2 ();
 DECAPx10_ASAP7_75t_R FILLER_123_24 ();
 DECAPx10_ASAP7_75t_R FILLER_123_46 ();
 DECAPx10_ASAP7_75t_R FILLER_123_68 ();
 DECAPx10_ASAP7_75t_R FILLER_123_90 ();
 DECAPx4_ASAP7_75t_R FILLER_123_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_122 ();
 DECAPx10_ASAP7_75t_R FILLER_123_128 ();
 DECAPx10_ASAP7_75t_R FILLER_123_150 ();
 DECAPx6_ASAP7_75t_R FILLER_123_172 ();
 DECAPx2_ASAP7_75t_R FILLER_123_186 ();
 DECAPx10_ASAP7_75t_R FILLER_123_243 ();
 DECAPx6_ASAP7_75t_R FILLER_123_265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_316 ();
 DECAPx10_ASAP7_75t_R FILLER_123_324 ();
 DECAPx10_ASAP7_75t_R FILLER_123_346 ();
 DECAPx10_ASAP7_75t_R FILLER_123_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_390 ();
 DECAPx10_ASAP7_75t_R FILLER_123_399 ();
 DECAPx10_ASAP7_75t_R FILLER_123_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_443 ();
 DECAPx10_ASAP7_75t_R FILLER_123_478 ();
 DECAPx1_ASAP7_75t_R FILLER_123_500 ();
 FILLER_ASAP7_75t_R FILLER_123_530 ();
 DECAPx1_ASAP7_75t_R FILLER_123_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_601 ();
 DECAPx6_ASAP7_75t_R FILLER_123_646 ();
 DECAPx4_ASAP7_75t_R FILLER_123_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_123_687 ();
 DECAPx1_ASAP7_75t_R FILLER_123_703 ();
 DECAPx10_ASAP7_75t_R FILLER_123_716 ();
 DECAPx4_ASAP7_75t_R FILLER_123_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_748 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_758 ();
 DECAPx6_ASAP7_75t_R FILLER_123_770 ();
 DECAPx1_ASAP7_75t_R FILLER_123_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_123_848 ();
 FILLER_ASAP7_75t_R FILLER_123_903 ();
 FILLER_ASAP7_75t_R FILLER_123_932 ();
 DECAPx10_ASAP7_75t_R FILLER_124_2 ();
 DECAPx10_ASAP7_75t_R FILLER_124_24 ();
 DECAPx10_ASAP7_75t_R FILLER_124_46 ();
 DECAPx4_ASAP7_75t_R FILLER_124_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_87 ();
 DECAPx1_ASAP7_75t_R FILLER_124_93 ();
 DECAPx6_ASAP7_75t_R FILLER_124_100 ();
 DECAPx1_ASAP7_75t_R FILLER_124_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_118 ();
 FILLER_ASAP7_75t_R FILLER_124_125 ();
 DECAPx10_ASAP7_75t_R FILLER_124_135 ();
 DECAPx10_ASAP7_75t_R FILLER_124_157 ();
 DECAPx6_ASAP7_75t_R FILLER_124_179 ();
 DECAPx2_ASAP7_75t_R FILLER_124_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_199 ();
 DECAPx2_ASAP7_75t_R FILLER_124_206 ();
 DECAPx10_ASAP7_75t_R FILLER_124_215 ();
 DECAPx4_ASAP7_75t_R FILLER_124_237 ();
 FILLER_ASAP7_75t_R FILLER_124_247 ();
 DECAPx2_ASAP7_75t_R FILLER_124_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_261 ();
 DECAPx10_ASAP7_75t_R FILLER_124_268 ();
 DECAPx2_ASAP7_75t_R FILLER_124_290 ();
 DECAPx2_ASAP7_75t_R FILLER_124_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_305 ();
 DECAPx6_ASAP7_75t_R FILLER_124_314 ();
 DECAPx2_ASAP7_75t_R FILLER_124_328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_357 ();
 DECAPx2_ASAP7_75t_R FILLER_124_367 ();
 DECAPx2_ASAP7_75t_R FILLER_124_376 ();
 DECAPx10_ASAP7_75t_R FILLER_124_388 ();
 DECAPx1_ASAP7_75t_R FILLER_124_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_414 ();
 FILLER_ASAP7_75t_R FILLER_124_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_436 ();
 DECAPx1_ASAP7_75t_R FILLER_124_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_464 ();
 DECAPx4_ASAP7_75t_R FILLER_124_473 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_483 ();
 DECAPx2_ASAP7_75t_R FILLER_124_498 ();
 DECAPx4_ASAP7_75t_R FILLER_124_550 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_560 ();
 DECAPx10_ASAP7_75t_R FILLER_124_568 ();
 DECAPx2_ASAP7_75t_R FILLER_124_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_596 ();
 DECAPx10_ASAP7_75t_R FILLER_124_603 ();
 DECAPx10_ASAP7_75t_R FILLER_124_625 ();
 DECAPx2_ASAP7_75t_R FILLER_124_647 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_689 ();
 FILLER_ASAP7_75t_R FILLER_124_702 ();
 DECAPx2_ASAP7_75t_R FILLER_124_707 ();
 FILLER_ASAP7_75t_R FILLER_124_713 ();
 DECAPx2_ASAP7_75t_R FILLER_124_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_124_727 ();
 DECAPx1_ASAP7_75t_R FILLER_124_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_751 ();
 DECAPx10_ASAP7_75t_R FILLER_124_762 ();
 DECAPx2_ASAP7_75t_R FILLER_124_784 ();
 FILLER_ASAP7_75t_R FILLER_124_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_798 ();
 DECAPx1_ASAP7_75t_R FILLER_124_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_806 ();
 DECAPx2_ASAP7_75t_R FILLER_124_827 ();
 DECAPx4_ASAP7_75t_R FILLER_124_841 ();
 FILLER_ASAP7_75t_R FILLER_124_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_124_907 ();
 DECAPx10_ASAP7_75t_R FILLER_125_2 ();
 DECAPx10_ASAP7_75t_R FILLER_125_24 ();
 DECAPx10_ASAP7_75t_R FILLER_125_46 ();
 DECAPx2_ASAP7_75t_R FILLER_125_68 ();
 FILLER_ASAP7_75t_R FILLER_125_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_102 ();
 FILLER_ASAP7_75t_R FILLER_125_151 ();
 DECAPx4_ASAP7_75t_R FILLER_125_162 ();
 DECAPx10_ASAP7_75t_R FILLER_125_187 ();
 DECAPx10_ASAP7_75t_R FILLER_125_209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_275 ();
 DECAPx1_ASAP7_75t_R FILLER_125_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_288 ();
 DECAPx4_ASAP7_75t_R FILLER_125_299 ();
 FILLER_ASAP7_75t_R FILLER_125_309 ();
 DECAPx1_ASAP7_75t_R FILLER_125_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_321 ();
 DECAPx2_ASAP7_75t_R FILLER_125_389 ();
 FILLER_ASAP7_75t_R FILLER_125_395 ();
 DECAPx2_ASAP7_75t_R FILLER_125_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_469 ();
 DECAPx10_ASAP7_75t_R FILLER_125_522 ();
 DECAPx1_ASAP7_75t_R FILLER_125_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_548 ();
 DECAPx6_ASAP7_75t_R FILLER_125_576 ();
 DECAPx2_ASAP7_75t_R FILLER_125_590 ();
 DECAPx6_ASAP7_75t_R FILLER_125_603 ();
 FILLER_ASAP7_75t_R FILLER_125_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_636 ();
 DECAPx1_ASAP7_75t_R FILLER_125_651 ();
 FILLER_ASAP7_75t_R FILLER_125_670 ();
 FILLER_ASAP7_75t_R FILLER_125_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_690 ();
 FILLER_ASAP7_75t_R FILLER_125_703 ();
 DECAPx2_ASAP7_75t_R FILLER_125_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_729 ();
 DECAPx4_ASAP7_75t_R FILLER_125_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_750 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_125_783 ();
 DECAPx10_ASAP7_75t_R FILLER_125_792 ();
 DECAPx6_ASAP7_75t_R FILLER_125_814 ();
 DECAPx1_ASAP7_75t_R FILLER_125_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_839 ();
 DECAPx2_ASAP7_75t_R FILLER_125_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_125_909 ();
 FILLER_ASAP7_75t_R FILLER_125_927 ();
 DECAPx10_ASAP7_75t_R FILLER_126_2 ();
 DECAPx10_ASAP7_75t_R FILLER_126_24 ();
 DECAPx10_ASAP7_75t_R FILLER_126_46 ();
 DECAPx2_ASAP7_75t_R FILLER_126_68 ();
 FILLER_ASAP7_75t_R FILLER_126_100 ();
 FILLER_ASAP7_75t_R FILLER_126_122 ();
 FILLER_ASAP7_75t_R FILLER_126_136 ();
 DECAPx10_ASAP7_75t_R FILLER_126_199 ();
 DECAPx2_ASAP7_75t_R FILLER_126_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_274 ();
 DECAPx6_ASAP7_75t_R FILLER_126_295 ();
 FILLER_ASAP7_75t_R FILLER_126_309 ();
 FILLER_ASAP7_75t_R FILLER_126_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_348 ();
 DECAPx2_ASAP7_75t_R FILLER_126_355 ();
 DECAPx1_ASAP7_75t_R FILLER_126_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_371 ();
 DECAPx6_ASAP7_75t_R FILLER_126_375 ();
 DECAPx2_ASAP7_75t_R FILLER_126_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_412 ();
 DECAPx2_ASAP7_75t_R FILLER_126_421 ();
 FILLER_ASAP7_75t_R FILLER_126_427 ();
 DECAPx10_ASAP7_75t_R FILLER_126_435 ();
 DECAPx1_ASAP7_75t_R FILLER_126_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_461 ();
 DECAPx4_ASAP7_75t_R FILLER_126_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_477 ();
 DECAPx1_ASAP7_75t_R FILLER_126_486 ();
 DECAPx2_ASAP7_75t_R FILLER_126_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_510 ();
 DECAPx10_ASAP7_75t_R FILLER_126_514 ();
 DECAPx10_ASAP7_75t_R FILLER_126_536 ();
 DECAPx6_ASAP7_75t_R FILLER_126_558 ();
 DECAPx2_ASAP7_75t_R FILLER_126_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_585 ();
 DECAPx4_ASAP7_75t_R FILLER_126_604 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_614 ();
 DECAPx10_ASAP7_75t_R FILLER_126_624 ();
 DECAPx6_ASAP7_75t_R FILLER_126_646 ();
 DECAPx1_ASAP7_75t_R FILLER_126_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_664 ();
 DECAPx2_ASAP7_75t_R FILLER_126_671 ();
 FILLER_ASAP7_75t_R FILLER_126_677 ();
 DECAPx4_ASAP7_75t_R FILLER_126_691 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_126_701 ();
 DECAPx6_ASAP7_75t_R FILLER_126_741 ();
 DECAPx2_ASAP7_75t_R FILLER_126_755 ();
 DECAPx10_ASAP7_75t_R FILLER_126_794 ();
 DECAPx6_ASAP7_75t_R FILLER_126_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_830 ();
 DECAPx6_ASAP7_75t_R FILLER_126_843 ();
 DECAPx2_ASAP7_75t_R FILLER_126_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_126_863 ();
 DECAPx1_ASAP7_75t_R FILLER_126_869 ();
 FILLER_ASAP7_75t_R FILLER_126_901 ();
 DECAPx10_ASAP7_75t_R FILLER_127_2 ();
 DECAPx10_ASAP7_75t_R FILLER_127_24 ();
 DECAPx10_ASAP7_75t_R FILLER_127_46 ();
 DECAPx4_ASAP7_75t_R FILLER_127_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_87 ();
 DECAPx10_ASAP7_75t_R FILLER_127_112 ();
 DECAPx6_ASAP7_75t_R FILLER_127_134 ();
 FILLER_ASAP7_75t_R FILLER_127_148 ();
 DECAPx4_ASAP7_75t_R FILLER_127_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_181 ();
 DECAPx1_ASAP7_75t_R FILLER_127_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_202 ();
 DECAPx1_ASAP7_75t_R FILLER_127_209 ();
 DECAPx1_ASAP7_75t_R FILLER_127_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_289 ();
 FILLER_ASAP7_75t_R FILLER_127_298 ();
 DECAPx2_ASAP7_75t_R FILLER_127_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_317 ();
 DECAPx6_ASAP7_75t_R FILLER_127_326 ();
 FILLER_ASAP7_75t_R FILLER_127_340 ();
 DECAPx10_ASAP7_75t_R FILLER_127_345 ();
 DECAPx1_ASAP7_75t_R FILLER_127_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_380 ();
 DECAPx10_ASAP7_75t_R FILLER_127_398 ();
 DECAPx2_ASAP7_75t_R FILLER_127_420 ();
 FILLER_ASAP7_75t_R FILLER_127_426 ();
 DECAPx6_ASAP7_75t_R FILLER_127_434 ();
 DECAPx1_ASAP7_75t_R FILLER_127_448 ();
 DECAPx10_ASAP7_75t_R FILLER_127_488 ();
 DECAPx4_ASAP7_75t_R FILLER_127_510 ();
 FILLER_ASAP7_75t_R FILLER_127_520 ();
 DECAPx10_ASAP7_75t_R FILLER_127_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_576 ();
 DECAPx1_ASAP7_75t_R FILLER_127_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_609 ();
 DECAPx10_ASAP7_75t_R FILLER_127_616 ();
 FILLER_ASAP7_75t_R FILLER_127_638 ();
 DECAPx10_ASAP7_75t_R FILLER_127_656 ();
 DECAPx10_ASAP7_75t_R FILLER_127_678 ();
 DECAPx10_ASAP7_75t_R FILLER_127_700 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_722 ();
 DECAPx6_ASAP7_75t_R FILLER_127_749 ();
 FILLER_ASAP7_75t_R FILLER_127_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_768 ();
 DECAPx4_ASAP7_75t_R FILLER_127_815 ();
 FILLER_ASAP7_75t_R FILLER_127_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_127_837 ();
 DECAPx2_ASAP7_75t_R FILLER_127_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_855 ();
 FILLER_ASAP7_75t_R FILLER_127_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_127_924 ();
 FILLER_ASAP7_75t_R FILLER_127_927 ();
 DECAPx10_ASAP7_75t_R FILLER_128_2 ();
 DECAPx10_ASAP7_75t_R FILLER_128_24 ();
 DECAPx10_ASAP7_75t_R FILLER_128_46 ();
 DECAPx6_ASAP7_75t_R FILLER_128_68 ();
 DECAPx2_ASAP7_75t_R FILLER_128_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_88 ();
 DECAPx10_ASAP7_75t_R FILLER_128_92 ();
 DECAPx10_ASAP7_75t_R FILLER_128_114 ();
 DECAPx10_ASAP7_75t_R FILLER_128_136 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_227 ();
 DECAPx6_ASAP7_75t_R FILLER_128_237 ();
 FILLER_ASAP7_75t_R FILLER_128_251 ();
 DECAPx1_ASAP7_75t_R FILLER_128_259 ();
 DECAPx6_ASAP7_75t_R FILLER_128_266 ();
 DECAPx1_ASAP7_75t_R FILLER_128_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_284 ();
 DECAPx4_ASAP7_75t_R FILLER_128_319 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_329 ();
 DECAPx6_ASAP7_75t_R FILLER_128_344 ();
 FILLER_ASAP7_75t_R FILLER_128_358 ();
 FILLER_ASAP7_75t_R FILLER_128_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_376 ();
 DECAPx1_ASAP7_75t_R FILLER_128_387 ();
 DECAPx2_ASAP7_75t_R FILLER_128_405 ();
 FILLER_ASAP7_75t_R FILLER_128_411 ();
 DECAPx10_ASAP7_75t_R FILLER_128_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_443 ();
 DECAPx2_ASAP7_75t_R FILLER_128_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_473 ();
 DECAPx4_ASAP7_75t_R FILLER_128_484 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_494 ();
 DECAPx2_ASAP7_75t_R FILLER_128_507 ();
 FILLER_ASAP7_75t_R FILLER_128_513 ();
 DECAPx1_ASAP7_75t_R FILLER_128_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_527 ();
 FILLER_ASAP7_75t_R FILLER_128_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_553 ();
 DECAPx1_ASAP7_75t_R FILLER_128_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_589 ();
 DECAPx1_ASAP7_75t_R FILLER_128_608 ();
 DECAPx2_ASAP7_75t_R FILLER_128_636 ();
 DECAPx4_ASAP7_75t_R FILLER_128_665 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_675 ();
 DECAPx2_ASAP7_75t_R FILLER_128_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_696 ();
 DECAPx6_ASAP7_75t_R FILLER_128_705 ();
 DECAPx1_ASAP7_75t_R FILLER_128_719 ();
 DECAPx4_ASAP7_75t_R FILLER_128_732 ();
 FILLER_ASAP7_75t_R FILLER_128_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_764 ();
 DECAPx4_ASAP7_75t_R FILLER_128_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_782 ();
 DECAPx2_ASAP7_75t_R FILLER_128_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_792 ();
 DECAPx1_ASAP7_75t_R FILLER_128_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_128_884 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_128_907 ();
 DECAPx10_ASAP7_75t_R FILLER_129_2 ();
 DECAPx10_ASAP7_75t_R FILLER_129_24 ();
 DECAPx10_ASAP7_75t_R FILLER_129_46 ();
 DECAPx10_ASAP7_75t_R FILLER_129_68 ();
 DECAPx10_ASAP7_75t_R FILLER_129_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_119 ();
 DECAPx2_ASAP7_75t_R FILLER_129_130 ();
 FILLER_ASAP7_75t_R FILLER_129_136 ();
 FILLER_ASAP7_75t_R FILLER_129_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_192 ();
 DECAPx2_ASAP7_75t_R FILLER_129_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_207 ();
 FILLER_ASAP7_75t_R FILLER_129_214 ();
 DECAPx10_ASAP7_75t_R FILLER_129_219 ();
 DECAPx10_ASAP7_75t_R FILLER_129_241 ();
 DECAPx10_ASAP7_75t_R FILLER_129_263 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_285 ();
 DECAPx6_ASAP7_75t_R FILLER_129_309 ();
 DECAPx1_ASAP7_75t_R FILLER_129_323 ();
 DECAPx1_ASAP7_75t_R FILLER_129_353 ();
 DECAPx1_ASAP7_75t_R FILLER_129_383 ();
 FILLER_ASAP7_75t_R FILLER_129_393 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_420 ();
 DECAPx4_ASAP7_75t_R FILLER_129_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_469 ();
 DECAPx2_ASAP7_75t_R FILLER_129_474 ();
 DECAPx2_ASAP7_75t_R FILLER_129_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_492 ();
 DECAPx2_ASAP7_75t_R FILLER_129_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_531 ();
 DECAPx6_ASAP7_75t_R FILLER_129_548 ();
 DECAPx6_ASAP7_75t_R FILLER_129_574 ();
 DECAPx2_ASAP7_75t_R FILLER_129_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_594 ();
 DECAPx2_ASAP7_75t_R FILLER_129_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_627 ();
 DECAPx2_ASAP7_75t_R FILLER_129_634 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_640 ();
 DECAPx6_ASAP7_75t_R FILLER_129_653 ();
 DECAPx1_ASAP7_75t_R FILLER_129_667 ();
 DECAPx4_ASAP7_75t_R FILLER_129_677 ();
 DECAPx6_ASAP7_75t_R FILLER_129_719 ();
 DECAPx1_ASAP7_75t_R FILLER_129_733 ();
 DECAPx6_ASAP7_75t_R FILLER_129_783 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_835 ();
 FILLER_ASAP7_75t_R FILLER_129_841 ();
 DECAPx2_ASAP7_75t_R FILLER_129_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_129_852 ();
 DECAPx2_ASAP7_75t_R FILLER_129_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_129_873 ();
 FILLER_ASAP7_75t_R FILLER_129_894 ();
 DECAPx1_ASAP7_75t_R FILLER_129_916 ();
 FILLER_ASAP7_75t_R FILLER_129_927 ();
 DECAPx10_ASAP7_75t_R FILLER_130_2 ();
 DECAPx10_ASAP7_75t_R FILLER_130_24 ();
 DECAPx10_ASAP7_75t_R FILLER_130_46 ();
 DECAPx6_ASAP7_75t_R FILLER_130_68 ();
 DECAPx2_ASAP7_75t_R FILLER_130_82 ();
 DECAPx2_ASAP7_75t_R FILLER_130_94 ();
 FILLER_ASAP7_75t_R FILLER_130_100 ();
 FILLER_ASAP7_75t_R FILLER_130_163 ();
 DECAPx10_ASAP7_75t_R FILLER_130_174 ();
 DECAPx4_ASAP7_75t_R FILLER_130_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_206 ();
 DECAPx2_ASAP7_75t_R FILLER_130_213 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_219 ();
 DECAPx10_ASAP7_75t_R FILLER_130_228 ();
 DECAPx10_ASAP7_75t_R FILLER_130_250 ();
 DECAPx10_ASAP7_75t_R FILLER_130_272 ();
 DECAPx6_ASAP7_75t_R FILLER_130_294 ();
 DECAPx2_ASAP7_75t_R FILLER_130_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_320 ();
 DECAPx6_ASAP7_75t_R FILLER_130_326 ();
 FILLER_ASAP7_75t_R FILLER_130_340 ();
 DECAPx6_ASAP7_75t_R FILLER_130_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_359 ();
 DECAPx1_ASAP7_75t_R FILLER_130_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_370 ();
 DECAPx10_ASAP7_75t_R FILLER_130_374 ();
 DECAPx10_ASAP7_75t_R FILLER_130_396 ();
 FILLER_ASAP7_75t_R FILLER_130_418 ();
 DECAPx1_ASAP7_75t_R FILLER_130_458 ();
 DECAPx10_ASAP7_75t_R FILLER_130_464 ();
 DECAPx4_ASAP7_75t_R FILLER_130_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_496 ();
 DECAPx10_ASAP7_75t_R FILLER_130_510 ();
 FILLER_ASAP7_75t_R FILLER_130_532 ();
 DECAPx10_ASAP7_75t_R FILLER_130_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_559 ();
 DECAPx6_ASAP7_75t_R FILLER_130_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_591 ();
 DECAPx1_ASAP7_75t_R FILLER_130_595 ();
 DECAPx4_ASAP7_75t_R FILLER_130_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_615 ();
 DECAPx10_ASAP7_75t_R FILLER_130_624 ();
 DECAPx4_ASAP7_75t_R FILLER_130_646 ();
 FILLER_ASAP7_75t_R FILLER_130_656 ();
 DECAPx2_ASAP7_75t_R FILLER_130_704 ();
 FILLER_ASAP7_75t_R FILLER_130_730 ();
 DECAPx4_ASAP7_75t_R FILLER_130_738 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_748 ();
 DECAPx4_ASAP7_75t_R FILLER_130_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_130_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_777 ();
 DECAPx6_ASAP7_75t_R FILLER_130_788 ();
 DECAPx2_ASAP7_75t_R FILLER_130_802 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_808 ();
 DECAPx10_ASAP7_75t_R FILLER_130_835 ();
 DECAPx6_ASAP7_75t_R FILLER_130_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_130_892 ();
 DECAPx10_ASAP7_75t_R FILLER_131_2 ();
 DECAPx10_ASAP7_75t_R FILLER_131_24 ();
 DECAPx10_ASAP7_75t_R FILLER_131_46 ();
 DECAPx2_ASAP7_75t_R FILLER_131_68 ();
 FILLER_ASAP7_75t_R FILLER_131_74 ();
 DECAPx2_ASAP7_75t_R FILLER_131_102 ();
 FILLER_ASAP7_75t_R FILLER_131_114 ();
 DECAPx4_ASAP7_75t_R FILLER_131_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_141 ();
 DECAPx10_ASAP7_75t_R FILLER_131_151 ();
 DECAPx10_ASAP7_75t_R FILLER_131_173 ();
 DECAPx4_ASAP7_75t_R FILLER_131_195 ();
 DECAPx2_ASAP7_75t_R FILLER_131_245 ();
 FILLER_ASAP7_75t_R FILLER_131_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_265 ();
 DECAPx1_ASAP7_75t_R FILLER_131_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_286 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_293 ();
 DECAPx2_ASAP7_75t_R FILLER_131_300 ();
 FILLER_ASAP7_75t_R FILLER_131_306 ();
 DECAPx6_ASAP7_75t_R FILLER_131_337 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_351 ();
 DECAPx2_ASAP7_75t_R FILLER_131_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_366 ();
 DECAPx2_ASAP7_75t_R FILLER_131_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_388 ();
 DECAPx2_ASAP7_75t_R FILLER_131_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_401 ();
 DECAPx10_ASAP7_75t_R FILLER_131_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_430 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_465 ();
 DECAPx4_ASAP7_75t_R FILLER_131_495 ();
 DECAPx2_ASAP7_75t_R FILLER_131_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_517 ();
 DECAPx10_ASAP7_75t_R FILLER_131_544 ();
 DECAPx1_ASAP7_75t_R FILLER_131_566 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_579 ();
 DECAPx10_ASAP7_75t_R FILLER_131_592 ();
 DECAPx6_ASAP7_75t_R FILLER_131_614 ();
 DECAPx1_ASAP7_75t_R FILLER_131_628 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_641 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_647 ();
 DECAPx10_ASAP7_75t_R FILLER_131_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_715 ();
 FILLER_ASAP7_75t_R FILLER_131_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_734 ();
 DECAPx6_ASAP7_75t_R FILLER_131_749 ();
 FILLER_ASAP7_75t_R FILLER_131_763 ();
 DECAPx6_ASAP7_75t_R FILLER_131_797 ();
 DECAPx1_ASAP7_75t_R FILLER_131_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_815 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_821 ();
 DECAPx6_ASAP7_75t_R FILLER_131_827 ();
 DECAPx1_ASAP7_75t_R FILLER_131_841 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_845 ();
 DECAPx2_ASAP7_75t_R FILLER_131_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_131_869 ();
 FILLER_ASAP7_75t_R FILLER_131_885 ();
 FILLER_ASAP7_75t_R FILLER_131_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_131_924 ();
 DECAPx10_ASAP7_75t_R FILLER_132_2 ();
 DECAPx10_ASAP7_75t_R FILLER_132_24 ();
 DECAPx10_ASAP7_75t_R FILLER_132_46 ();
 DECAPx6_ASAP7_75t_R FILLER_132_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_93 ();
 DECAPx6_ASAP7_75t_R FILLER_132_100 ();
 DECAPx2_ASAP7_75t_R FILLER_132_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_120 ();
 DECAPx1_ASAP7_75t_R FILLER_132_129 ();
 DECAPx10_ASAP7_75t_R FILLER_132_139 ();
 DECAPx6_ASAP7_75t_R FILLER_132_161 ();
 FILLER_ASAP7_75t_R FILLER_132_175 ();
 FILLER_ASAP7_75t_R FILLER_132_184 ();
 DECAPx1_ASAP7_75t_R FILLER_132_192 ();
 DECAPx4_ASAP7_75t_R FILLER_132_202 ();
 DECAPx4_ASAP7_75t_R FILLER_132_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_237 ();
 DECAPx4_ASAP7_75t_R FILLER_132_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_251 ();
 FILLER_ASAP7_75t_R FILLER_132_280 ();
 DECAPx1_ASAP7_75t_R FILLER_132_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_312 ();
 DECAPx6_ASAP7_75t_R FILLER_132_319 ();
 DECAPx1_ASAP7_75t_R FILLER_132_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_347 ();
 DECAPx2_ASAP7_75t_R FILLER_132_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_392 ();
 FILLER_ASAP7_75t_R FILLER_132_401 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_409 ();
 DECAPx1_ASAP7_75t_R FILLER_132_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_424 ();
 DECAPx10_ASAP7_75t_R FILLER_132_429 ();
 DECAPx4_ASAP7_75t_R FILLER_132_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_461 ();
 DECAPx4_ASAP7_75t_R FILLER_132_464 ();
 FILLER_ASAP7_75t_R FILLER_132_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_486 ();
 DECAPx10_ASAP7_75t_R FILLER_132_493 ();
 DECAPx1_ASAP7_75t_R FILLER_132_515 ();
 DECAPx2_ASAP7_75t_R FILLER_132_526 ();
 FILLER_ASAP7_75t_R FILLER_132_532 ();
 DECAPx2_ASAP7_75t_R FILLER_132_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_565 ();
 DECAPx6_ASAP7_75t_R FILLER_132_596 ();
 FILLER_ASAP7_75t_R FILLER_132_610 ();
 DECAPx1_ASAP7_75t_R FILLER_132_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_623 ();
 FILLER_ASAP7_75t_R FILLER_132_656 ();
 DECAPx1_ASAP7_75t_R FILLER_132_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_669 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_679 ();
 DECAPx6_ASAP7_75t_R FILLER_132_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_705 ();
 DECAPx4_ASAP7_75t_R FILLER_132_712 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_722 ();
 DECAPx10_ASAP7_75t_R FILLER_132_754 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_132_776 ();
 DECAPx4_ASAP7_75t_R FILLER_132_808 ();
 DECAPx10_ASAP7_75t_R FILLER_132_823 ();
 DECAPx1_ASAP7_75t_R FILLER_132_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_132_886 ();
 FILLER_ASAP7_75t_R FILLER_132_906 ();
 DECAPx10_ASAP7_75t_R FILLER_133_2 ();
 DECAPx10_ASAP7_75t_R FILLER_133_24 ();
 DECAPx10_ASAP7_75t_R FILLER_133_46 ();
 DECAPx10_ASAP7_75t_R FILLER_133_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_90 ();
 DECAPx6_ASAP7_75t_R FILLER_133_111 ();
 DECAPx2_ASAP7_75t_R FILLER_133_125 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_131 ();
 DECAPx2_ASAP7_75t_R FILLER_133_152 ();
 DECAPx4_ASAP7_75t_R FILLER_133_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_210 ();
 DECAPx4_ASAP7_75t_R FILLER_133_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_227 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_273 ();
 DECAPx6_ASAP7_75t_R FILLER_133_283 ();
 DECAPx10_ASAP7_75t_R FILLER_133_300 ();
 DECAPx2_ASAP7_75t_R FILLER_133_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_328 ();
 DECAPx1_ASAP7_75t_R FILLER_133_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_372 ();
 DECAPx2_ASAP7_75t_R FILLER_133_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_433 ();
 DECAPx2_ASAP7_75t_R FILLER_133_444 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_450 ();
 DECAPx6_ASAP7_75t_R FILLER_133_462 ();
 DECAPx1_ASAP7_75t_R FILLER_133_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_480 ();
 DECAPx2_ASAP7_75t_R FILLER_133_484 ();
 DECAPx1_ASAP7_75t_R FILLER_133_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_502 ();
 FILLER_ASAP7_75t_R FILLER_133_511 ();
 FILLER_ASAP7_75t_R FILLER_133_519 ();
 DECAPx6_ASAP7_75t_R FILLER_133_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_541 ();
 FILLER_ASAP7_75t_R FILLER_133_549 ();
 DECAPx2_ASAP7_75t_R FILLER_133_568 ();
 DECAPx1_ASAP7_75t_R FILLER_133_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_629 ();
 FILLER_ASAP7_75t_R FILLER_133_638 ();
 DECAPx4_ASAP7_75t_R FILLER_133_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_674 ();
 DECAPx6_ASAP7_75t_R FILLER_133_686 ();
 FILLER_ASAP7_75t_R FILLER_133_706 ();
 DECAPx4_ASAP7_75t_R FILLER_133_716 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_734 ();
 DECAPx2_ASAP7_75t_R FILLER_133_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_759 ();
 DECAPx1_ASAP7_75t_R FILLER_133_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_771 ();
 DECAPx4_ASAP7_75t_R FILLER_133_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_785 ();
 FILLER_ASAP7_75t_R FILLER_133_798 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_133_806 ();
 DECAPx6_ASAP7_75t_R FILLER_133_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_857 ();
 DECAPx4_ASAP7_75t_R FILLER_133_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_871 ();
 DECAPx10_ASAP7_75t_R FILLER_133_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_133_899 ();
 DECAPx10_ASAP7_75t_R FILLER_134_2 ();
 DECAPx10_ASAP7_75t_R FILLER_134_24 ();
 DECAPx10_ASAP7_75t_R FILLER_134_46 ();
 DECAPx10_ASAP7_75t_R FILLER_134_68 ();
 DECAPx2_ASAP7_75t_R FILLER_134_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_96 ();
 DECAPx1_ASAP7_75t_R FILLER_134_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_127 ();
 DECAPx10_ASAP7_75t_R FILLER_134_134 ();
 DECAPx4_ASAP7_75t_R FILLER_134_156 ();
 FILLER_ASAP7_75t_R FILLER_134_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_217 ();
 DECAPx10_ASAP7_75t_R FILLER_134_268 ();
 DECAPx6_ASAP7_75t_R FILLER_134_290 ();
 DECAPx1_ASAP7_75t_R FILLER_134_304 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_320 ();
 DECAPx6_ASAP7_75t_R FILLER_134_341 ();
 DECAPx2_ASAP7_75t_R FILLER_134_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_361 ();
 DECAPx2_ASAP7_75t_R FILLER_134_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_410 ();
 FILLER_ASAP7_75t_R FILLER_134_414 ();
 DECAPx2_ASAP7_75t_R FILLER_134_419 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_425 ();
 DECAPx1_ASAP7_75t_R FILLER_134_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_464 ();
 DECAPx1_ASAP7_75t_R FILLER_134_471 ();
 FILLER_ASAP7_75t_R FILLER_134_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_518 ();
 FILLER_ASAP7_75t_R FILLER_134_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_585 ();
 FILLER_ASAP7_75t_R FILLER_134_597 ();
 DECAPx2_ASAP7_75t_R FILLER_134_613 ();
 DECAPx4_ASAP7_75t_R FILLER_134_635 ();
 FILLER_ASAP7_75t_R FILLER_134_645 ();
 DECAPx10_ASAP7_75t_R FILLER_134_659 ();
 DECAPx4_ASAP7_75t_R FILLER_134_681 ();
 DECAPx4_ASAP7_75t_R FILLER_134_699 ();
 DECAPx10_ASAP7_75t_R FILLER_134_715 ();
 DECAPx6_ASAP7_75t_R FILLER_134_737 ();
 DECAPx4_ASAP7_75t_R FILLER_134_783 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_134_839 ();
 FILLER_ASAP7_75t_R FILLER_134_849 ();
 DECAPx10_ASAP7_75t_R FILLER_134_862 ();
 DECAPx2_ASAP7_75t_R FILLER_134_884 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_134_890 ();
 DECAPx10_ASAP7_75t_R FILLER_135_2 ();
 DECAPx10_ASAP7_75t_R FILLER_135_24 ();
 DECAPx10_ASAP7_75t_R FILLER_135_46 ();
 DECAPx6_ASAP7_75t_R FILLER_135_68 ();
 DECAPx1_ASAP7_75t_R FILLER_135_82 ();
 DECAPx4_ASAP7_75t_R FILLER_135_95 ();
 DECAPx4_ASAP7_75t_R FILLER_135_134 ();
 FILLER_ASAP7_75t_R FILLER_135_144 ();
 DECAPx4_ASAP7_75t_R FILLER_135_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_168 ();
 DECAPx1_ASAP7_75t_R FILLER_135_177 ();
 DECAPx6_ASAP7_75t_R FILLER_135_196 ();
 DECAPx1_ASAP7_75t_R FILLER_135_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_220 ();
 DECAPx1_ASAP7_75t_R FILLER_135_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_237 ();
 DECAPx1_ASAP7_75t_R FILLER_135_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_266 ();
 DECAPx2_ASAP7_75t_R FILLER_135_273 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_299 ();
 DECAPx10_ASAP7_75t_R FILLER_135_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_391 ();
 DECAPx1_ASAP7_75t_R FILLER_135_414 ();
 DECAPx4_ASAP7_75t_R FILLER_135_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_434 ();
 FILLER_ASAP7_75t_R FILLER_135_440 ();
 DECAPx4_ASAP7_75t_R FILLER_135_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_455 ();
 DECAPx1_ASAP7_75t_R FILLER_135_486 ();
 FILLER_ASAP7_75t_R FILLER_135_496 ();
 DECAPx2_ASAP7_75t_R FILLER_135_510 ();
 DECAPx1_ASAP7_75t_R FILLER_135_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_560 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_583 ();
 DECAPx1_ASAP7_75t_R FILLER_135_592 ();
 DECAPx10_ASAP7_75t_R FILLER_135_611 ();
 DECAPx10_ASAP7_75t_R FILLER_135_633 ();
 FILLER_ASAP7_75t_R FILLER_135_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_673 ();
 DECAPx10_ASAP7_75t_R FILLER_135_689 ();
 DECAPx2_ASAP7_75t_R FILLER_135_711 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_738 ();
 DECAPx4_ASAP7_75t_R FILLER_135_749 ();
 FILLER_ASAP7_75t_R FILLER_135_759 ();
 DECAPx10_ASAP7_75t_R FILLER_135_775 ();
 FILLER_ASAP7_75t_R FILLER_135_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_832 ();
 FILLER_ASAP7_75t_R FILLER_135_859 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_135_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_135_933 ();
 DECAPx10_ASAP7_75t_R FILLER_136_2 ();
 DECAPx10_ASAP7_75t_R FILLER_136_24 ();
 DECAPx10_ASAP7_75t_R FILLER_136_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_68 ();
 DECAPx6_ASAP7_75t_R FILLER_136_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_117 ();
 DECAPx6_ASAP7_75t_R FILLER_136_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_145 ();
 DECAPx2_ASAP7_75t_R FILLER_136_149 ();
 FILLER_ASAP7_75t_R FILLER_136_155 ();
 DECAPx10_ASAP7_75t_R FILLER_136_172 ();
 DECAPx10_ASAP7_75t_R FILLER_136_194 ();
 DECAPx10_ASAP7_75t_R FILLER_136_216 ();
 DECAPx6_ASAP7_75t_R FILLER_136_238 ();
 DECAPx1_ASAP7_75t_R FILLER_136_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_256 ();
 DECAPx1_ASAP7_75t_R FILLER_136_283 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_313 ();
 DECAPx2_ASAP7_75t_R FILLER_136_319 ();
 FILLER_ASAP7_75t_R FILLER_136_347 ();
 DECAPx2_ASAP7_75t_R FILLER_136_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_373 ();
 DECAPx2_ASAP7_75t_R FILLER_136_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_406 ();
 DECAPx2_ASAP7_75t_R FILLER_136_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_439 ();
 FILLER_ASAP7_75t_R FILLER_136_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_461 ();
 DECAPx6_ASAP7_75t_R FILLER_136_464 ();
 DECAPx2_ASAP7_75t_R FILLER_136_478 ();
 DECAPx10_ASAP7_75t_R FILLER_136_498 ();
 DECAPx4_ASAP7_75t_R FILLER_136_520 ();
 DECAPx4_ASAP7_75t_R FILLER_136_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_569 ();
 DECAPx6_ASAP7_75t_R FILLER_136_578 ();
 DECAPx4_ASAP7_75t_R FILLER_136_598 ();
 DECAPx6_ASAP7_75t_R FILLER_136_620 ();
 DECAPx1_ASAP7_75t_R FILLER_136_634 ();
 DECAPx1_ASAP7_75t_R FILLER_136_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_655 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_666 ();
 DECAPx2_ASAP7_75t_R FILLER_136_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_691 ();
 FILLER_ASAP7_75t_R FILLER_136_704 ();
 FILLER_ASAP7_75t_R FILLER_136_714 ();
 DECAPx4_ASAP7_75t_R FILLER_136_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_762 ();
 DECAPx10_ASAP7_75t_R FILLER_136_766 ();
 DECAPx10_ASAP7_75t_R FILLER_136_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_810 ();
 DECAPx2_ASAP7_75t_R FILLER_136_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_820 ();
 DECAPx2_ASAP7_75t_R FILLER_136_826 ();
 FILLER_ASAP7_75t_R FILLER_136_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_136_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_136_928 ();
 DECAPx10_ASAP7_75t_R FILLER_137_2 ();
 DECAPx10_ASAP7_75t_R FILLER_137_24 ();
 DECAPx10_ASAP7_75t_R FILLER_137_46 ();
 DECAPx4_ASAP7_75t_R FILLER_137_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_78 ();
 DECAPx10_ASAP7_75t_R FILLER_137_90 ();
 DECAPx6_ASAP7_75t_R FILLER_137_112 ();
 FILLER_ASAP7_75t_R FILLER_137_126 ();
 DECAPx10_ASAP7_75t_R FILLER_137_180 ();
 DECAPx6_ASAP7_75t_R FILLER_137_202 ();
 DECAPx1_ASAP7_75t_R FILLER_137_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_226 ();
 DECAPx10_ASAP7_75t_R FILLER_137_233 ();
 FILLER_ASAP7_75t_R FILLER_137_255 ();
 DECAPx2_ASAP7_75t_R FILLER_137_263 ();
 FILLER_ASAP7_75t_R FILLER_137_269 ();
 DECAPx2_ASAP7_75t_R FILLER_137_274 ();
 FILLER_ASAP7_75t_R FILLER_137_280 ();
 FILLER_ASAP7_75t_R FILLER_137_299 ();
 DECAPx10_ASAP7_75t_R FILLER_137_304 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_326 ();
 DECAPx10_ASAP7_75t_R FILLER_137_353 ();
 DECAPx4_ASAP7_75t_R FILLER_137_375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_385 ();
 FILLER_ASAP7_75t_R FILLER_137_420 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_451 ();
 DECAPx10_ASAP7_75t_R FILLER_137_468 ();
 DECAPx2_ASAP7_75t_R FILLER_137_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_502 ();
 DECAPx10_ASAP7_75t_R FILLER_137_515 ();
 DECAPx4_ASAP7_75t_R FILLER_137_537 ();
 DECAPx6_ASAP7_75t_R FILLER_137_550 ();
 DECAPx1_ASAP7_75t_R FILLER_137_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_568 ();
 DECAPx4_ASAP7_75t_R FILLER_137_572 ();
 DECAPx6_ASAP7_75t_R FILLER_137_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_608 ();
 DECAPx1_ASAP7_75t_R FILLER_137_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_621 ();
 DECAPx6_ASAP7_75t_R FILLER_137_631 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_645 ();
 DECAPx2_ASAP7_75t_R FILLER_137_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_658 ();
 DECAPx1_ASAP7_75t_R FILLER_137_666 ();
 DECAPx6_ASAP7_75t_R FILLER_137_701 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_715 ();
 FILLER_ASAP7_75t_R FILLER_137_729 ();
 DECAPx4_ASAP7_75t_R FILLER_137_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_752 ();
 FILLER_ASAP7_75t_R FILLER_137_765 ();
 DECAPx4_ASAP7_75t_R FILLER_137_783 ();
 DECAPx10_ASAP7_75t_R FILLER_137_799 ();
 DECAPx10_ASAP7_75t_R FILLER_137_821 ();
 DECAPx2_ASAP7_75t_R FILLER_137_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_849 ();
 FILLER_ASAP7_75t_R FILLER_137_855 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_137_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_137_895 ();
 FILLER_ASAP7_75t_R FILLER_137_932 ();
 DECAPx10_ASAP7_75t_R FILLER_138_2 ();
 DECAPx10_ASAP7_75t_R FILLER_138_24 ();
 DECAPx10_ASAP7_75t_R FILLER_138_46 ();
 DECAPx10_ASAP7_75t_R FILLER_138_68 ();
 DECAPx2_ASAP7_75t_R FILLER_138_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_96 ();
 DECAPx10_ASAP7_75t_R FILLER_138_103 ();
 DECAPx6_ASAP7_75t_R FILLER_138_125 ();
 DECAPx1_ASAP7_75t_R FILLER_138_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_143 ();
 DECAPx1_ASAP7_75t_R FILLER_138_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_154 ();
 FILLER_ASAP7_75t_R FILLER_138_161 ();
 DECAPx6_ASAP7_75t_R FILLER_138_172 ();
 FILLER_ASAP7_75t_R FILLER_138_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_194 ();
 DECAPx1_ASAP7_75t_R FILLER_138_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_204 ();
 DECAPx1_ASAP7_75t_R FILLER_138_208 ();
 DECAPx1_ASAP7_75t_R FILLER_138_218 ();
 DECAPx2_ASAP7_75t_R FILLER_138_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_254 ();
 DECAPx6_ASAP7_75t_R FILLER_138_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_295 ();
 DECAPx10_ASAP7_75t_R FILLER_138_302 ();
 DECAPx2_ASAP7_75t_R FILLER_138_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_330 ();
 DECAPx10_ASAP7_75t_R FILLER_138_346 ();
 DECAPx1_ASAP7_75t_R FILLER_138_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_379 ();
 FILLER_ASAP7_75t_R FILLER_138_410 ();
 DECAPx2_ASAP7_75t_R FILLER_138_456 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_464 ();
 DECAPx10_ASAP7_75t_R FILLER_138_473 ();
 DECAPx4_ASAP7_75t_R FILLER_138_495 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_505 ();
 DECAPx2_ASAP7_75t_R FILLER_138_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_520 ();
 DECAPx10_ASAP7_75t_R FILLER_138_528 ();
 DECAPx4_ASAP7_75t_R FILLER_138_550 ();
 FILLER_ASAP7_75t_R FILLER_138_560 ();
 DECAPx4_ASAP7_75t_R FILLER_138_577 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_587 ();
 DECAPx2_ASAP7_75t_R FILLER_138_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_608 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_138_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_677 ();
 DECAPx2_ASAP7_75t_R FILLER_138_688 ();
 FILLER_ASAP7_75t_R FILLER_138_694 ();
 DECAPx6_ASAP7_75t_R FILLER_138_712 ();
 DECAPx2_ASAP7_75t_R FILLER_138_726 ();
 FILLER_ASAP7_75t_R FILLER_138_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_775 ();
 FILLER_ASAP7_75t_R FILLER_138_790 ();
 DECAPx10_ASAP7_75t_R FILLER_138_818 ();
 DECAPx4_ASAP7_75t_R FILLER_138_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_850 ();
 FILLER_ASAP7_75t_R FILLER_138_856 ();
 DECAPx1_ASAP7_75t_R FILLER_138_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_138_933 ();
 DECAPx10_ASAP7_75t_R FILLER_139_2 ();
 DECAPx10_ASAP7_75t_R FILLER_139_24 ();
 DECAPx10_ASAP7_75t_R FILLER_139_46 ();
 DECAPx6_ASAP7_75t_R FILLER_139_68 ();
 DECAPx1_ASAP7_75t_R FILLER_139_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_86 ();
 FILLER_ASAP7_75t_R FILLER_139_115 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_123 ();
 DECAPx6_ASAP7_75t_R FILLER_139_134 ();
 FILLER_ASAP7_75t_R FILLER_139_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_211 ();
 DECAPx1_ASAP7_75t_R FILLER_139_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_224 ();
 DECAPx1_ASAP7_75t_R FILLER_139_259 ();
 DECAPx10_ASAP7_75t_R FILLER_139_272 ();
 FILLER_ASAP7_75t_R FILLER_139_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_304 ();
 DECAPx2_ASAP7_75t_R FILLER_139_311 ();
 DECAPx6_ASAP7_75t_R FILLER_139_323 ();
 DECAPx2_ASAP7_75t_R FILLER_139_337 ();
 DECAPx2_ASAP7_75t_R FILLER_139_346 ();
 DECAPx1_ASAP7_75t_R FILLER_139_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_362 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_371 ();
 FILLER_ASAP7_75t_R FILLER_139_402 ();
 DECAPx2_ASAP7_75t_R FILLER_139_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_437 ();
 DECAPx1_ASAP7_75t_R FILLER_139_452 ();
 DECAPx6_ASAP7_75t_R FILLER_139_491 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_514 ();
 DECAPx4_ASAP7_75t_R FILLER_139_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_551 ();
 DECAPx2_ASAP7_75t_R FILLER_139_560 ();
 FILLER_ASAP7_75t_R FILLER_139_566 ();
 DECAPx2_ASAP7_75t_R FILLER_139_588 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_635 ();
 DECAPx2_ASAP7_75t_R FILLER_139_644 ();
 FILLER_ASAP7_75t_R FILLER_139_650 ();
 DECAPx2_ASAP7_75t_R FILLER_139_658 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_664 ();
 DECAPx6_ASAP7_75t_R FILLER_139_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_689 ();
 FILLER_ASAP7_75t_R FILLER_139_701 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_722 ();
 DECAPx10_ASAP7_75t_R FILLER_139_728 ();
 DECAPx1_ASAP7_75t_R FILLER_139_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_760 ();
 FILLER_ASAP7_75t_R FILLER_139_804 ();
 FILLER_ASAP7_75t_R FILLER_139_836 ();
 DECAPx10_ASAP7_75t_R FILLER_139_841 ();
 DECAPx2_ASAP7_75t_R FILLER_139_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_139_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_139_924 ();
 FILLER_ASAP7_75t_R FILLER_139_932 ();
 DECAPx10_ASAP7_75t_R FILLER_140_2 ();
 DECAPx10_ASAP7_75t_R FILLER_140_24 ();
 DECAPx10_ASAP7_75t_R FILLER_140_46 ();
 DECAPx2_ASAP7_75t_R FILLER_140_68 ();
 FILLER_ASAP7_75t_R FILLER_140_74 ();
 DECAPx2_ASAP7_75t_R FILLER_140_102 ();
 FILLER_ASAP7_75t_R FILLER_140_108 ();
 DECAPx6_ASAP7_75t_R FILLER_140_148 ();
 DECAPx1_ASAP7_75t_R FILLER_140_162 ();
 FILLER_ASAP7_75t_R FILLER_140_181 ();
 DECAPx10_ASAP7_75t_R FILLER_140_252 ();
 DECAPx6_ASAP7_75t_R FILLER_140_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_288 ();
 DECAPx1_ASAP7_75t_R FILLER_140_295 ();
 FILLER_ASAP7_75t_R FILLER_140_305 ();
 FILLER_ASAP7_75t_R FILLER_140_343 ();
 DECAPx10_ASAP7_75t_R FILLER_140_385 ();
 DECAPx4_ASAP7_75t_R FILLER_140_407 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_417 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_436 ();
 DECAPx1_ASAP7_75t_R FILLER_140_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_461 ();
 DECAPx2_ASAP7_75t_R FILLER_140_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_530 ();
 FILLER_ASAP7_75t_R FILLER_140_544 ();
 DECAPx4_ASAP7_75t_R FILLER_140_564 ();
 FILLER_ASAP7_75t_R FILLER_140_574 ();
 DECAPx2_ASAP7_75t_R FILLER_140_596 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_602 ();
 DECAPx2_ASAP7_75t_R FILLER_140_625 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_631 ();
 DECAPx6_ASAP7_75t_R FILLER_140_646 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_678 ();
 DECAPx6_ASAP7_75t_R FILLER_140_685 ();
 DECAPx1_ASAP7_75t_R FILLER_140_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_703 ();
 DECAPx10_ASAP7_75t_R FILLER_140_736 ();
 DECAPx10_ASAP7_75t_R FILLER_140_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_140_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_140_811 ();
 DECAPx1_ASAP7_75t_R FILLER_140_821 ();
 FILLER_ASAP7_75t_R FILLER_140_851 ();
 FILLER_ASAP7_75t_R FILLER_140_879 ();
 FILLER_ASAP7_75t_R FILLER_140_906 ();
 DECAPx10_ASAP7_75t_R FILLER_141_2 ();
 DECAPx10_ASAP7_75t_R FILLER_141_24 ();
 DECAPx10_ASAP7_75t_R FILLER_141_46 ();
 DECAPx6_ASAP7_75t_R FILLER_141_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_88 ();
 DECAPx6_ASAP7_75t_R FILLER_141_94 ();
 DECAPx1_ASAP7_75t_R FILLER_141_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_119 ();
 DECAPx2_ASAP7_75t_R FILLER_141_162 ();
 FILLER_ASAP7_75t_R FILLER_141_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_176 ();
 DECAPx2_ASAP7_75t_R FILLER_141_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_191 ();
 DECAPx10_ASAP7_75t_R FILLER_141_224 ();
 DECAPx6_ASAP7_75t_R FILLER_141_246 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_260 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_269 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_278 ();
 DECAPx1_ASAP7_75t_R FILLER_141_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_319 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_369 ();
 DECAPx4_ASAP7_75t_R FILLER_141_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_398 ();
 DECAPx4_ASAP7_75t_R FILLER_141_409 ();
 DECAPx2_ASAP7_75t_R FILLER_141_446 ();
 FILLER_ASAP7_75t_R FILLER_141_452 ();
 FILLER_ASAP7_75t_R FILLER_141_460 ();
 FILLER_ASAP7_75t_R FILLER_141_470 ();
 DECAPx1_ASAP7_75t_R FILLER_141_484 ();
 DECAPx1_ASAP7_75t_R FILLER_141_496 ();
 DECAPx2_ASAP7_75t_R FILLER_141_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_521 ();
 FILLER_ASAP7_75t_R FILLER_141_559 ();
 DECAPx4_ASAP7_75t_R FILLER_141_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_601 ();
 DECAPx6_ASAP7_75t_R FILLER_141_618 ();
 DECAPx2_ASAP7_75t_R FILLER_141_632 ();
 FILLER_ASAP7_75t_R FILLER_141_648 ();
 DECAPx6_ASAP7_75t_R FILLER_141_656 ();
 DECAPx2_ASAP7_75t_R FILLER_141_670 ();
 DECAPx4_ASAP7_75t_R FILLER_141_702 ();
 FILLER_ASAP7_75t_R FILLER_141_712 ();
 DECAPx10_ASAP7_75t_R FILLER_141_762 ();
 DECAPx4_ASAP7_75t_R FILLER_141_784 ();
 DECAPx10_ASAP7_75t_R FILLER_141_797 ();
 DECAPx1_ASAP7_75t_R FILLER_141_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_141_902 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_141_908 ();
 FILLER_ASAP7_75t_R FILLER_141_923 ();
 FILLER_ASAP7_75t_R FILLER_141_927 ();
 DECAPx10_ASAP7_75t_R FILLER_142_2 ();
 DECAPx10_ASAP7_75t_R FILLER_142_24 ();
 DECAPx10_ASAP7_75t_R FILLER_142_46 ();
 DECAPx6_ASAP7_75t_R FILLER_142_68 ();
 DECAPx2_ASAP7_75t_R FILLER_142_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_88 ();
 DECAPx6_ASAP7_75t_R FILLER_142_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_109 ();
 DECAPx10_ASAP7_75t_R FILLER_142_154 ();
 DECAPx10_ASAP7_75t_R FILLER_142_176 ();
 DECAPx10_ASAP7_75t_R FILLER_142_198 ();
 DECAPx6_ASAP7_75t_R FILLER_142_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_234 ();
 DECAPx6_ASAP7_75t_R FILLER_142_240 ();
 FILLER_ASAP7_75t_R FILLER_142_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_271 ();
 DECAPx1_ASAP7_75t_R FILLER_142_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_284 ();
 DECAPx1_ASAP7_75t_R FILLER_142_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_295 ();
 DECAPx2_ASAP7_75t_R FILLER_142_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_305 ();
 FILLER_ASAP7_75t_R FILLER_142_314 ();
 DECAPx1_ASAP7_75t_R FILLER_142_323 ();
 FILLER_ASAP7_75t_R FILLER_142_344 ();
 DECAPx6_ASAP7_75t_R FILLER_142_371 ();
 DECAPx1_ASAP7_75t_R FILLER_142_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_416 ();
 DECAPx1_ASAP7_75t_R FILLER_142_426 ();
 DECAPx10_ASAP7_75t_R FILLER_142_436 ();
 DECAPx1_ASAP7_75t_R FILLER_142_458 ();
 DECAPx6_ASAP7_75t_R FILLER_142_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_478 ();
 DECAPx1_ASAP7_75t_R FILLER_142_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_557 ();
 DECAPx10_ASAP7_75t_R FILLER_142_576 ();
 DECAPx10_ASAP7_75t_R FILLER_142_598 ();
 DECAPx10_ASAP7_75t_R FILLER_142_620 ();
 DECAPx1_ASAP7_75t_R FILLER_142_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_646 ();
 DECAPx6_ASAP7_75t_R FILLER_142_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_679 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_686 ();
 DECAPx1_ASAP7_75t_R FILLER_142_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_765 ();
 DECAPx1_ASAP7_75t_R FILLER_142_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_794 ();
 FILLER_ASAP7_75t_R FILLER_142_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_142_864 ();
 DECAPx2_ASAP7_75t_R FILLER_142_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_142_895 ();
 FILLER_ASAP7_75t_R FILLER_142_906 ();
 DECAPx10_ASAP7_75t_R FILLER_143_2 ();
 DECAPx10_ASAP7_75t_R FILLER_143_24 ();
 DECAPx10_ASAP7_75t_R FILLER_143_46 ();
 DECAPx4_ASAP7_75t_R FILLER_143_68 ();
 FILLER_ASAP7_75t_R FILLER_143_78 ();
 FILLER_ASAP7_75t_R FILLER_143_106 ();
 DECAPx2_ASAP7_75t_R FILLER_143_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_156 ();
 DECAPx10_ASAP7_75t_R FILLER_143_169 ();
 DECAPx10_ASAP7_75t_R FILLER_143_191 ();
 DECAPx2_ASAP7_75t_R FILLER_143_213 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_248 ();
 DECAPx10_ASAP7_75t_R FILLER_143_286 ();
 DECAPx10_ASAP7_75t_R FILLER_143_308 ();
 DECAPx4_ASAP7_75t_R FILLER_143_330 ();
 FILLER_ASAP7_75t_R FILLER_143_346 ();
 DECAPx6_ASAP7_75t_R FILLER_143_354 ();
 DECAPx1_ASAP7_75t_R FILLER_143_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_379 ();
 FILLER_ASAP7_75t_R FILLER_143_388 ();
 DECAPx2_ASAP7_75t_R FILLER_143_396 ();
 FILLER_ASAP7_75t_R FILLER_143_402 ();
 FILLER_ASAP7_75t_R FILLER_143_407 ();
 DECAPx10_ASAP7_75t_R FILLER_143_415 ();
 DECAPx2_ASAP7_75t_R FILLER_143_437 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_443 ();
 DECAPx10_ASAP7_75t_R FILLER_143_452 ();
 DECAPx10_ASAP7_75t_R FILLER_143_474 ();
 FILLER_ASAP7_75t_R FILLER_143_496 ();
 DECAPx2_ASAP7_75t_R FILLER_143_504 ();
 FILLER_ASAP7_75t_R FILLER_143_510 ();
 DECAPx10_ASAP7_75t_R FILLER_143_518 ();
 DECAPx6_ASAP7_75t_R FILLER_143_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_554 ();
 DECAPx2_ASAP7_75t_R FILLER_143_565 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_571 ();
 DECAPx1_ASAP7_75t_R FILLER_143_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_586 ();
 DECAPx4_ASAP7_75t_R FILLER_143_596 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_606 ();
 DECAPx2_ASAP7_75t_R FILLER_143_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_656 ();
 DECAPx10_ASAP7_75t_R FILLER_143_673 ();
 DECAPx10_ASAP7_75t_R FILLER_143_695 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_143_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_736 ();
 DECAPx6_ASAP7_75t_R FILLER_143_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_815 ();
 DECAPx6_ASAP7_75t_R FILLER_143_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_143_848 ();
 FILLER_ASAP7_75t_R FILLER_143_864 ();
 DECAPx1_ASAP7_75t_R FILLER_143_880 ();
 FILLER_ASAP7_75t_R FILLER_143_901 ();
 FILLER_ASAP7_75t_R FILLER_143_927 ();
 DECAPx10_ASAP7_75t_R FILLER_144_2 ();
 DECAPx10_ASAP7_75t_R FILLER_144_24 ();
 DECAPx10_ASAP7_75t_R FILLER_144_46 ();
 DECAPx6_ASAP7_75t_R FILLER_144_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_91 ();
 DECAPx2_ASAP7_75t_R FILLER_144_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_141 ();
 DECAPx2_ASAP7_75t_R FILLER_144_148 ();
 FILLER_ASAP7_75t_R FILLER_144_154 ();
 DECAPx10_ASAP7_75t_R FILLER_144_164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_186 ();
 DECAPx1_ASAP7_75t_R FILLER_144_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_208 ();
 DECAPx2_ASAP7_75t_R FILLER_144_217 ();
 FILLER_ASAP7_75t_R FILLER_144_223 ();
 FILLER_ASAP7_75t_R FILLER_144_263 ();
 DECAPx2_ASAP7_75t_R FILLER_144_268 ();
 FILLER_ASAP7_75t_R FILLER_144_274 ();
 DECAPx10_ASAP7_75t_R FILLER_144_282 ();
 DECAPx2_ASAP7_75t_R FILLER_144_304 ();
 FILLER_ASAP7_75t_R FILLER_144_310 ();
 DECAPx1_ASAP7_75t_R FILLER_144_326 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_387 ();
 DECAPx1_ASAP7_75t_R FILLER_144_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_407 ();
 DECAPx10_ASAP7_75t_R FILLER_144_416 ();
 DECAPx2_ASAP7_75t_R FILLER_144_438 ();
 FILLER_ASAP7_75t_R FILLER_144_444 ();
 DECAPx1_ASAP7_75t_R FILLER_144_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_461 ();
 DECAPx2_ASAP7_75t_R FILLER_144_464 ();
 DECAPx10_ASAP7_75t_R FILLER_144_478 ();
 DECAPx4_ASAP7_75t_R FILLER_144_500 ();
 FILLER_ASAP7_75t_R FILLER_144_510 ();
 DECAPx2_ASAP7_75t_R FILLER_144_531 ();
 FILLER_ASAP7_75t_R FILLER_144_537 ();
 DECAPx2_ASAP7_75t_R FILLER_144_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_555 ();
 DECAPx2_ASAP7_75t_R FILLER_144_562 ();
 FILLER_ASAP7_75t_R FILLER_144_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_581 ();
 FILLER_ASAP7_75t_R FILLER_144_612 ();
 DECAPx1_ASAP7_75t_R FILLER_144_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_659 ();
 DECAPx10_ASAP7_75t_R FILLER_144_666 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_144_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_703 ();
 DECAPx2_ASAP7_75t_R FILLER_144_714 ();
 FILLER_ASAP7_75t_R FILLER_144_720 ();
 DECAPx10_ASAP7_75t_R FILLER_144_727 ();
 DECAPx4_ASAP7_75t_R FILLER_144_749 ();
 FILLER_ASAP7_75t_R FILLER_144_769 ();
 DECAPx10_ASAP7_75t_R FILLER_144_811 ();
 DECAPx6_ASAP7_75t_R FILLER_144_833 ();
 DECAPx2_ASAP7_75t_R FILLER_144_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_144_933 ();
 DECAPx10_ASAP7_75t_R FILLER_145_2 ();
 DECAPx10_ASAP7_75t_R FILLER_145_24 ();
 DECAPx10_ASAP7_75t_R FILLER_145_46 ();
 DECAPx10_ASAP7_75t_R FILLER_145_68 ();
 DECAPx10_ASAP7_75t_R FILLER_145_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_112 ();
 DECAPx4_ASAP7_75t_R FILLER_145_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_157 ();
 DECAPx2_ASAP7_75t_R FILLER_145_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_172 ();
 FILLER_ASAP7_75t_R FILLER_145_223 ();
 FILLER_ASAP7_75t_R FILLER_145_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_239 ();
 DECAPx2_ASAP7_75t_R FILLER_145_249 ();
 FILLER_ASAP7_75t_R FILLER_145_255 ();
 DECAPx10_ASAP7_75t_R FILLER_145_260 ();
 DECAPx2_ASAP7_75t_R FILLER_145_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_288 ();
 FILLER_ASAP7_75t_R FILLER_145_295 ();
 FILLER_ASAP7_75t_R FILLER_145_300 ();
 DECAPx1_ASAP7_75t_R FILLER_145_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_319 ();
 FILLER_ASAP7_75t_R FILLER_145_333 ();
 DECAPx1_ASAP7_75t_R FILLER_145_341 ();
 DECAPx4_ASAP7_75t_R FILLER_145_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_388 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_418 ();
 DECAPx6_ASAP7_75t_R FILLER_145_427 ();
 DECAPx1_ASAP7_75t_R FILLER_145_455 ();
 FILLER_ASAP7_75t_R FILLER_145_469 ();
 DECAPx6_ASAP7_75t_R FILLER_145_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_507 ();
 DECAPx6_ASAP7_75t_R FILLER_145_534 ();
 DECAPx1_ASAP7_75t_R FILLER_145_548 ();
 DECAPx10_ASAP7_75t_R FILLER_145_557 ();
 FILLER_ASAP7_75t_R FILLER_145_579 ();
 FILLER_ASAP7_75t_R FILLER_145_593 ();
 DECAPx4_ASAP7_75t_R FILLER_145_601 ();
 DECAPx2_ASAP7_75t_R FILLER_145_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_637 ();
 DECAPx4_ASAP7_75t_R FILLER_145_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_664 ();
 DECAPx6_ASAP7_75t_R FILLER_145_689 ();
 FILLER_ASAP7_75t_R FILLER_145_703 ();
 DECAPx10_ASAP7_75t_R FILLER_145_731 ();
 DECAPx10_ASAP7_75t_R FILLER_145_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_781 ();
 DECAPx10_ASAP7_75t_R FILLER_145_785 ();
 DECAPx1_ASAP7_75t_R FILLER_145_807 ();
 DECAPx6_ASAP7_75t_R FILLER_145_819 ();
 FILLER_ASAP7_75t_R FILLER_145_833 ();
 DECAPx6_ASAP7_75t_R FILLER_145_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_145_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_883 ();
 DECAPx2_ASAP7_75t_R FILLER_145_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_145_933 ();
 DECAPx10_ASAP7_75t_R FILLER_146_2 ();
 DECAPx10_ASAP7_75t_R FILLER_146_24 ();
 DECAPx10_ASAP7_75t_R FILLER_146_46 ();
 DECAPx10_ASAP7_75t_R FILLER_146_68 ();
 DECAPx10_ASAP7_75t_R FILLER_146_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_112 ();
 FILLER_ASAP7_75t_R FILLER_146_121 ();
 DECAPx6_ASAP7_75t_R FILLER_146_129 ();
 DECAPx6_ASAP7_75t_R FILLER_146_146 ();
 DECAPx2_ASAP7_75t_R FILLER_146_160 ();
 DECAPx4_ASAP7_75t_R FILLER_146_198 ();
 DECAPx10_ASAP7_75t_R FILLER_146_220 ();
 DECAPx10_ASAP7_75t_R FILLER_146_242 ();
 DECAPx2_ASAP7_75t_R FILLER_146_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_312 ();
 DECAPx10_ASAP7_75t_R FILLER_146_335 ();
 DECAPx1_ASAP7_75t_R FILLER_146_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_361 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_368 ();
 FILLER_ASAP7_75t_R FILLER_146_377 ();
 DECAPx1_ASAP7_75t_R FILLER_146_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_389 ();
 DECAPx2_ASAP7_75t_R FILLER_146_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_402 ();
 DECAPx6_ASAP7_75t_R FILLER_146_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_420 ();
 FILLER_ASAP7_75t_R FILLER_146_429 ();
 DECAPx1_ASAP7_75t_R FILLER_146_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_461 ();
 FILLER_ASAP7_75t_R FILLER_146_464 ();
 DECAPx10_ASAP7_75t_R FILLER_146_499 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_521 ();
 DECAPx1_ASAP7_75t_R FILLER_146_531 ();
 DECAPx2_ASAP7_75t_R FILLER_146_549 ();
 DECAPx2_ASAP7_75t_R FILLER_146_558 ();
 FILLER_ASAP7_75t_R FILLER_146_564 ();
 FILLER_ASAP7_75t_R FILLER_146_573 ();
 DECAPx1_ASAP7_75t_R FILLER_146_582 ();
 DECAPx10_ASAP7_75t_R FILLER_146_589 ();
 DECAPx10_ASAP7_75t_R FILLER_146_611 ();
 DECAPx10_ASAP7_75t_R FILLER_146_633 ();
 DECAPx2_ASAP7_75t_R FILLER_146_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_661 ();
 DECAPx1_ASAP7_75t_R FILLER_146_670 ();
 DECAPx1_ASAP7_75t_R FILLER_146_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_688 ();
 FILLER_ASAP7_75t_R FILLER_146_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_719 ();
 DECAPx2_ASAP7_75t_R FILLER_146_723 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_729 ();
 FILLER_ASAP7_75t_R FILLER_146_735 ();
 DECAPx10_ASAP7_75t_R FILLER_146_750 ();
 DECAPx10_ASAP7_75t_R FILLER_146_772 ();
 DECAPx2_ASAP7_75t_R FILLER_146_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_800 ();
 DECAPx6_ASAP7_75t_R FILLER_146_859 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_146_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_146_915 ();
 DECAPx10_ASAP7_75t_R FILLER_147_2 ();
 DECAPx10_ASAP7_75t_R FILLER_147_24 ();
 DECAPx10_ASAP7_75t_R FILLER_147_46 ();
 DECAPx10_ASAP7_75t_R FILLER_147_68 ();
 DECAPx4_ASAP7_75t_R FILLER_147_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_100 ();
 DECAPx1_ASAP7_75t_R FILLER_147_107 ();
 DECAPx10_ASAP7_75t_R FILLER_147_137 ();
 DECAPx1_ASAP7_75t_R FILLER_147_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_176 ();
 DECAPx10_ASAP7_75t_R FILLER_147_191 ();
 DECAPx4_ASAP7_75t_R FILLER_147_213 ();
 FILLER_ASAP7_75t_R FILLER_147_223 ();
 DECAPx6_ASAP7_75t_R FILLER_147_245 ();
 DECAPx1_ASAP7_75t_R FILLER_147_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_263 ();
 DECAPx2_ASAP7_75t_R FILLER_147_278 ();
 FILLER_ASAP7_75t_R FILLER_147_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_292 ();
 DECAPx6_ASAP7_75t_R FILLER_147_298 ();
 DECAPx1_ASAP7_75t_R FILLER_147_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_323 ();
 DECAPx10_ASAP7_75t_R FILLER_147_330 ();
 DECAPx10_ASAP7_75t_R FILLER_147_352 ();
 DECAPx10_ASAP7_75t_R FILLER_147_374 ();
 DECAPx6_ASAP7_75t_R FILLER_147_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_453 ();
 DECAPx6_ASAP7_75t_R FILLER_147_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_474 ();
 DECAPx6_ASAP7_75t_R FILLER_147_505 ();
 FILLER_ASAP7_75t_R FILLER_147_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_539 ();
 DECAPx10_ASAP7_75t_R FILLER_147_569 ();
 DECAPx10_ASAP7_75t_R FILLER_147_591 ();
 DECAPx6_ASAP7_75t_R FILLER_147_613 ();
 DECAPx4_ASAP7_75t_R FILLER_147_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_645 ();
 DECAPx10_ASAP7_75t_R FILLER_147_655 ();
 DECAPx1_ASAP7_75t_R FILLER_147_677 ();
 DECAPx6_ASAP7_75t_R FILLER_147_687 ();
 DECAPx4_ASAP7_75t_R FILLER_147_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_716 ();
 FILLER_ASAP7_75t_R FILLER_147_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_778 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_809 ();
 DECAPx1_ASAP7_75t_R FILLER_147_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_820 ();
 DECAPx6_ASAP7_75t_R FILLER_147_824 ();
 DECAPx2_ASAP7_75t_R FILLER_147_848 ();
 DECAPx1_ASAP7_75t_R FILLER_147_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_865 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_147_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_147_919 ();
 FILLER_ASAP7_75t_R FILLER_147_927 ();
 DECAPx10_ASAP7_75t_R FILLER_148_2 ();
 DECAPx10_ASAP7_75t_R FILLER_148_24 ();
 DECAPx10_ASAP7_75t_R FILLER_148_46 ();
 DECAPx10_ASAP7_75t_R FILLER_148_68 ();
 FILLER_ASAP7_75t_R FILLER_148_90 ();
 DECAPx2_ASAP7_75t_R FILLER_148_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_124 ();
 DECAPx6_ASAP7_75t_R FILLER_148_128 ();
 DECAPx2_ASAP7_75t_R FILLER_148_148 ();
 FILLER_ASAP7_75t_R FILLER_148_154 ();
 DECAPx10_ASAP7_75t_R FILLER_148_164 ();
 DECAPx2_ASAP7_75t_R FILLER_148_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_202 ();
 DECAPx2_ASAP7_75t_R FILLER_148_215 ();
 DECAPx4_ASAP7_75t_R FILLER_148_247 ();
 DECAPx10_ASAP7_75t_R FILLER_148_275 ();
 FILLER_ASAP7_75t_R FILLER_148_297 ();
 DECAPx4_ASAP7_75t_R FILLER_148_302 ();
 DECAPx4_ASAP7_75t_R FILLER_148_318 ();
 FILLER_ASAP7_75t_R FILLER_148_340 ();
 DECAPx1_ASAP7_75t_R FILLER_148_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_360 ();
 DECAPx1_ASAP7_75t_R FILLER_148_369 ();
 DECAPx10_ASAP7_75t_R FILLER_148_376 ();
 DECAPx6_ASAP7_75t_R FILLER_148_398 ();
 DECAPx1_ASAP7_75t_R FILLER_148_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_416 ();
 DECAPx4_ASAP7_75t_R FILLER_148_446 ();
 FILLER_ASAP7_75t_R FILLER_148_470 ();
 DECAPx4_ASAP7_75t_R FILLER_148_475 ();
 FILLER_ASAP7_75t_R FILLER_148_485 ();
 DECAPx4_ASAP7_75t_R FILLER_148_513 ();
 FILLER_ASAP7_75t_R FILLER_148_523 ();
 DECAPx2_ASAP7_75t_R FILLER_148_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_543 ();
 DECAPx2_ASAP7_75t_R FILLER_148_552 ();
 DECAPx6_ASAP7_75t_R FILLER_148_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_609 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_148_623 ();
 DECAPx2_ASAP7_75t_R FILLER_148_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_642 ();
 DECAPx6_ASAP7_75t_R FILLER_148_663 ();
 FILLER_ASAP7_75t_R FILLER_148_677 ();
 DECAPx4_ASAP7_75t_R FILLER_148_694 ();
 DECAPx2_ASAP7_75t_R FILLER_148_713 ();
 DECAPx1_ASAP7_75t_R FILLER_148_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_744 ();
 FILLER_ASAP7_75t_R FILLER_148_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_763 ();
 DECAPx1_ASAP7_75t_R FILLER_148_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_820 ();
 DECAPx2_ASAP7_75t_R FILLER_148_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_837 ();
 DECAPx2_ASAP7_75t_R FILLER_148_844 ();
 FILLER_ASAP7_75t_R FILLER_148_850 ();
 FILLER_ASAP7_75t_R FILLER_148_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_148_913 ();
 DECAPx10_ASAP7_75t_R FILLER_149_2 ();
 DECAPx10_ASAP7_75t_R FILLER_149_24 ();
 DECAPx10_ASAP7_75t_R FILLER_149_46 ();
 DECAPx10_ASAP7_75t_R FILLER_149_68 ();
 DECAPx2_ASAP7_75t_R FILLER_149_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_103 ();
 DECAPx10_ASAP7_75t_R FILLER_149_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_131 ();
 DECAPx10_ASAP7_75t_R FILLER_149_164 ();
 DECAPx2_ASAP7_75t_R FILLER_149_186 ();
 FILLER_ASAP7_75t_R FILLER_149_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_253 ();
 DECAPx4_ASAP7_75t_R FILLER_149_280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_299 ();
 DECAPx10_ASAP7_75t_R FILLER_149_384 ();
 DECAPx10_ASAP7_75t_R FILLER_149_406 ();
 DECAPx2_ASAP7_75t_R FILLER_149_428 ();
 FILLER_ASAP7_75t_R FILLER_149_434 ();
 DECAPx4_ASAP7_75t_R FILLER_149_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_456 ();
 DECAPx2_ASAP7_75t_R FILLER_149_483 ();
 DECAPx2_ASAP7_75t_R FILLER_149_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_512 ();
 FILLER_ASAP7_75t_R FILLER_149_518 ();
 DECAPx4_ASAP7_75t_R FILLER_149_542 ();
 FILLER_ASAP7_75t_R FILLER_149_588 ();
 DECAPx2_ASAP7_75t_R FILLER_149_627 ();
 DECAPx6_ASAP7_75t_R FILLER_149_667 ();
 DECAPx1_ASAP7_75t_R FILLER_149_693 ();
 DECAPx6_ASAP7_75t_R FILLER_149_725 ();
 DECAPx1_ASAP7_75t_R FILLER_149_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_743 ();
 DECAPx2_ASAP7_75t_R FILLER_149_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_149_765 ();
 FILLER_ASAP7_75t_R FILLER_149_777 ();
 FILLER_ASAP7_75t_R FILLER_149_782 ();
 DECAPx10_ASAP7_75t_R FILLER_149_811 ();
 DECAPx6_ASAP7_75t_R FILLER_149_833 ();
 DECAPx1_ASAP7_75t_R FILLER_149_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_149_851 ();
 DECAPx4_ASAP7_75t_R FILLER_149_868 ();
 DECAPx1_ASAP7_75t_R FILLER_149_881 ();
 FILLER_ASAP7_75t_R FILLER_149_932 ();
 DECAPx10_ASAP7_75t_R FILLER_150_2 ();
 DECAPx10_ASAP7_75t_R FILLER_150_24 ();
 DECAPx10_ASAP7_75t_R FILLER_150_46 ();
 DECAPx10_ASAP7_75t_R FILLER_150_68 ();
 DECAPx6_ASAP7_75t_R FILLER_150_90 ();
 DECAPx2_ASAP7_75t_R FILLER_150_104 ();
 DECAPx6_ASAP7_75t_R FILLER_150_116 ();
 DECAPx2_ASAP7_75t_R FILLER_150_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_136 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_143 ();
 FILLER_ASAP7_75t_R FILLER_150_149 ();
 DECAPx2_ASAP7_75t_R FILLER_150_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_176 ();
 DECAPx1_ASAP7_75t_R FILLER_150_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_238 ();
 DECAPx1_ASAP7_75t_R FILLER_150_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_306 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_313 ();
 DECAPx6_ASAP7_75t_R FILLER_150_319 ();
 DECAPx1_ASAP7_75t_R FILLER_150_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_337 ();
 DECAPx1_ASAP7_75t_R FILLER_150_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_385 ();
 DECAPx6_ASAP7_75t_R FILLER_150_420 ();
 DECAPx2_ASAP7_75t_R FILLER_150_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_440 ();
 DECAPx1_ASAP7_75t_R FILLER_150_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_468 ();
 DECAPx10_ASAP7_75t_R FILLER_150_475 ();
 DECAPx4_ASAP7_75t_R FILLER_150_497 ();
 DECAPx1_ASAP7_75t_R FILLER_150_529 ();
 DECAPx2_ASAP7_75t_R FILLER_150_549 ();
 FILLER_ASAP7_75t_R FILLER_150_571 ();
 DECAPx4_ASAP7_75t_R FILLER_150_585 ();
 FILLER_ASAP7_75t_R FILLER_150_595 ();
 DECAPx1_ASAP7_75t_R FILLER_150_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_630 ();
 DECAPx2_ASAP7_75t_R FILLER_150_641 ();
 DECAPx1_ASAP7_75t_R FILLER_150_656 ();
 DECAPx4_ASAP7_75t_R FILLER_150_677 ();
 FILLER_ASAP7_75t_R FILLER_150_692 ();
 DECAPx10_ASAP7_75t_R FILLER_150_727 ();
 DECAPx2_ASAP7_75t_R FILLER_150_749 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_755 ();
 DECAPx4_ASAP7_75t_R FILLER_150_782 ();
 DECAPx6_ASAP7_75t_R FILLER_150_797 ();
 FILLER_ASAP7_75t_R FILLER_150_811 ();
 DECAPx1_ASAP7_75t_R FILLER_150_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_150_824 ();
 DECAPx10_ASAP7_75t_R FILLER_150_851 ();
 DECAPx4_ASAP7_75t_R FILLER_150_873 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_150_883 ();
 DECAPx1_ASAP7_75t_R FILLER_150_897 ();
 DECAPx10_ASAP7_75t_R FILLER_151_2 ();
 DECAPx10_ASAP7_75t_R FILLER_151_24 ();
 DECAPx10_ASAP7_75t_R FILLER_151_46 ();
 DECAPx6_ASAP7_75t_R FILLER_151_68 ();
 DECAPx2_ASAP7_75t_R FILLER_151_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_88 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_95 ();
 FILLER_ASAP7_75t_R FILLER_151_104 ();
 DECAPx1_ASAP7_75t_R FILLER_151_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_124 ();
 DECAPx6_ASAP7_75t_R FILLER_151_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_151 ();
 FILLER_ASAP7_75t_R FILLER_151_162 ();
 DECAPx1_ASAP7_75t_R FILLER_151_190 ();
 DECAPx2_ASAP7_75t_R FILLER_151_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_206 ();
 DECAPx1_ASAP7_75t_R FILLER_151_213 ();
 FILLER_ASAP7_75t_R FILLER_151_229 ();
 FILLER_ASAP7_75t_R FILLER_151_238 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_248 ();
 DECAPx6_ASAP7_75t_R FILLER_151_259 ();
 DECAPx1_ASAP7_75t_R FILLER_151_273 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_285 ();
 DECAPx4_ASAP7_75t_R FILLER_151_297 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_307 ();
 DECAPx2_ASAP7_75t_R FILLER_151_322 ();
 FILLER_ASAP7_75t_R FILLER_151_328 ();
 DECAPx1_ASAP7_75t_R FILLER_151_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_340 ();
 DECAPx1_ASAP7_75t_R FILLER_151_344 ();
 DECAPx6_ASAP7_75t_R FILLER_151_351 ();
 DECAPx2_ASAP7_75t_R FILLER_151_365 ();
 FILLER_ASAP7_75t_R FILLER_151_416 ();
 DECAPx1_ASAP7_75t_R FILLER_151_470 ();
 DECAPx2_ASAP7_75t_R FILLER_151_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_531 ();
 FILLER_ASAP7_75t_R FILLER_151_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_565 ();
 DECAPx10_ASAP7_75t_R FILLER_151_576 ();
 DECAPx2_ASAP7_75t_R FILLER_151_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_604 ();
 DECAPx6_ASAP7_75t_R FILLER_151_617 ();
 FILLER_ASAP7_75t_R FILLER_151_631 ();
 DECAPx1_ASAP7_75t_R FILLER_151_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_645 ();
 FILLER_ASAP7_75t_R FILLER_151_665 ();
 DECAPx1_ASAP7_75t_R FILLER_151_683 ();
 DECAPx1_ASAP7_75t_R FILLER_151_735 ();
 DECAPx10_ASAP7_75t_R FILLER_151_780 ();
 DECAPx2_ASAP7_75t_R FILLER_151_802 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_151_808 ();
 DECAPx1_ASAP7_75t_R FILLER_151_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_857 ();
 DECAPx6_ASAP7_75t_R FILLER_151_864 ();
 DECAPx1_ASAP7_75t_R FILLER_151_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_151_924 ();
 FILLER_ASAP7_75t_R FILLER_151_927 ();
 DECAPx10_ASAP7_75t_R FILLER_152_2 ();
 DECAPx10_ASAP7_75t_R FILLER_152_24 ();
 DECAPx10_ASAP7_75t_R FILLER_152_46 ();
 DECAPx6_ASAP7_75t_R FILLER_152_68 ();
 DECAPx1_ASAP7_75t_R FILLER_152_119 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_139 ();
 DECAPx4_ASAP7_75t_R FILLER_152_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_158 ();
 FILLER_ASAP7_75t_R FILLER_152_167 ();
 DECAPx10_ASAP7_75t_R FILLER_152_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_211 ();
 DECAPx10_ASAP7_75t_R FILLER_152_246 ();
 DECAPx2_ASAP7_75t_R FILLER_152_268 ();
 FILLER_ASAP7_75t_R FILLER_152_274 ();
 FILLER_ASAP7_75t_R FILLER_152_302 ();
 DECAPx1_ASAP7_75t_R FILLER_152_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_375 ();
 FILLER_ASAP7_75t_R FILLER_152_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_461 ();
 DECAPx2_ASAP7_75t_R FILLER_152_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_531 ();
 DECAPx6_ASAP7_75t_R FILLER_152_566 ();
 FILLER_ASAP7_75t_R FILLER_152_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_585 ();
 DECAPx10_ASAP7_75t_R FILLER_152_592 ();
 DECAPx4_ASAP7_75t_R FILLER_152_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_624 ();
 DECAPx10_ASAP7_75t_R FILLER_152_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_665 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_152_673 ();
 DECAPx10_ASAP7_75t_R FILLER_152_686 ();
 DECAPx2_ASAP7_75t_R FILLER_152_708 ();
 DECAPx10_ASAP7_75t_R FILLER_152_717 ();
 DECAPx6_ASAP7_75t_R FILLER_152_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_753 ();
 DECAPx10_ASAP7_75t_R FILLER_152_757 ();
 DECAPx6_ASAP7_75t_R FILLER_152_779 ();
 DECAPx1_ASAP7_75t_R FILLER_152_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_797 ();
 DECAPx1_ASAP7_75t_R FILLER_152_810 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_814 ();
 FILLER_ASAP7_75t_R FILLER_152_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_835 ();
 DECAPx4_ASAP7_75t_R FILLER_152_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_152_902 ();
 DECAPx10_ASAP7_75t_R FILLER_153_2 ();
 DECAPx10_ASAP7_75t_R FILLER_153_24 ();
 DECAPx10_ASAP7_75t_R FILLER_153_46 ();
 DECAPx10_ASAP7_75t_R FILLER_153_68 ();
 DECAPx2_ASAP7_75t_R FILLER_153_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_96 ();
 DECAPx6_ASAP7_75t_R FILLER_153_100 ();
 DECAPx2_ASAP7_75t_R FILLER_153_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_120 ();
 DECAPx6_ASAP7_75t_R FILLER_153_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_176 ();
 DECAPx10_ASAP7_75t_R FILLER_153_190 ();
 DECAPx10_ASAP7_75t_R FILLER_153_212 ();
 DECAPx4_ASAP7_75t_R FILLER_153_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_251 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_258 ();
 FILLER_ASAP7_75t_R FILLER_153_265 ();
 DECAPx2_ASAP7_75t_R FILLER_153_273 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_288 ();
 DECAPx10_ASAP7_75t_R FILLER_153_294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_316 ();
 DECAPx1_ASAP7_75t_R FILLER_153_322 ();
 DECAPx2_ASAP7_75t_R FILLER_153_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_390 ();
 DECAPx6_ASAP7_75t_R FILLER_153_394 ();
 DECAPx1_ASAP7_75t_R FILLER_153_408 ();
 DECAPx4_ASAP7_75t_R FILLER_153_446 ();
 FILLER_ASAP7_75t_R FILLER_153_456 ();
 DECAPx10_ASAP7_75t_R FILLER_153_468 ();
 DECAPx10_ASAP7_75t_R FILLER_153_516 ();
 DECAPx4_ASAP7_75t_R FILLER_153_538 ();
 DECAPx6_ASAP7_75t_R FILLER_153_559 ();
 FILLER_ASAP7_75t_R FILLER_153_573 ();
 DECAPx6_ASAP7_75t_R FILLER_153_596 ();
 DECAPx2_ASAP7_75t_R FILLER_153_616 ();
 FILLER_ASAP7_75t_R FILLER_153_622 ();
 DECAPx10_ASAP7_75t_R FILLER_153_636 ();
 DECAPx6_ASAP7_75t_R FILLER_153_658 ();
 FILLER_ASAP7_75t_R FILLER_153_672 ();
 DECAPx2_ASAP7_75t_R FILLER_153_683 ();
 FILLER_ASAP7_75t_R FILLER_153_689 ();
 DECAPx10_ASAP7_75t_R FILLER_153_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_153_729 ();
 DECAPx10_ASAP7_75t_R FILLER_153_739 ();
 DECAPx4_ASAP7_75t_R FILLER_153_761 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_771 ();
 FILLER_ASAP7_75t_R FILLER_153_784 ();
 DECAPx2_ASAP7_75t_R FILLER_153_819 ();
 DECAPx4_ASAP7_75t_R FILLER_153_828 ();
 FILLER_ASAP7_75t_R FILLER_153_838 ();
 FILLER_ASAP7_75t_R FILLER_153_854 ();
 DECAPx6_ASAP7_75t_R FILLER_153_888 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_153_902 ();
 FILLER_ASAP7_75t_R FILLER_153_932 ();
 DECAPx10_ASAP7_75t_R FILLER_154_2 ();
 DECAPx10_ASAP7_75t_R FILLER_154_24 ();
 DECAPx10_ASAP7_75t_R FILLER_154_46 ();
 DECAPx4_ASAP7_75t_R FILLER_154_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_87 ();
 DECAPx10_ASAP7_75t_R FILLER_154_97 ();
 DECAPx6_ASAP7_75t_R FILLER_154_119 ();
 DECAPx1_ASAP7_75t_R FILLER_154_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_144 ();
 DECAPx10_ASAP7_75t_R FILLER_154_150 ();
 DECAPx10_ASAP7_75t_R FILLER_154_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_194 ();
 FILLER_ASAP7_75t_R FILLER_154_238 ();
 DECAPx1_ASAP7_75t_R FILLER_154_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_252 ();
 DECAPx1_ASAP7_75t_R FILLER_154_261 ();
 DECAPx10_ASAP7_75t_R FILLER_154_271 ();
 DECAPx10_ASAP7_75t_R FILLER_154_293 ();
 DECAPx6_ASAP7_75t_R FILLER_154_315 ();
 FILLER_ASAP7_75t_R FILLER_154_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_361 ();
 DECAPx10_ASAP7_75t_R FILLER_154_368 ();
 DECAPx10_ASAP7_75t_R FILLER_154_390 ();
 DECAPx1_ASAP7_75t_R FILLER_154_412 ();
 DECAPx10_ASAP7_75t_R FILLER_154_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_461 ();
 DECAPx10_ASAP7_75t_R FILLER_154_464 ();
 DECAPx1_ASAP7_75t_R FILLER_154_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_490 ();
 DECAPx10_ASAP7_75t_R FILLER_154_511 ();
 DECAPx10_ASAP7_75t_R FILLER_154_533 ();
 DECAPx4_ASAP7_75t_R FILLER_154_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_580 ();
 DECAPx4_ASAP7_75t_R FILLER_154_596 ();
 FILLER_ASAP7_75t_R FILLER_154_614 ();
 DECAPx6_ASAP7_75t_R FILLER_154_625 ();
 DECAPx4_ASAP7_75t_R FILLER_154_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_154_667 ();
 DECAPx4_ASAP7_75t_R FILLER_154_688 ();
 FILLER_ASAP7_75t_R FILLER_154_698 ();
 DECAPx4_ASAP7_75t_R FILLER_154_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_716 ();
 DECAPx2_ASAP7_75t_R FILLER_154_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_749 ();
 DECAPx10_ASAP7_75t_R FILLER_154_811 ();
 DECAPx2_ASAP7_75t_R FILLER_154_833 ();
 FILLER_ASAP7_75t_R FILLER_154_839 ();
 FILLER_ASAP7_75t_R FILLER_154_867 ();
 DECAPx4_ASAP7_75t_R FILLER_154_882 ();
 FILLER_ASAP7_75t_R FILLER_154_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_154_907 ();
 DECAPx10_ASAP7_75t_R FILLER_155_2 ();
 DECAPx10_ASAP7_75t_R FILLER_155_24 ();
 DECAPx10_ASAP7_75t_R FILLER_155_46 ();
 DECAPx2_ASAP7_75t_R FILLER_155_68 ();
 FILLER_ASAP7_75t_R FILLER_155_74 ();
 DECAPx10_ASAP7_75t_R FILLER_155_112 ();
 DECAPx2_ASAP7_75t_R FILLER_155_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_140 ();
 DECAPx6_ASAP7_75t_R FILLER_155_152 ();
 DECAPx1_ASAP7_75t_R FILLER_155_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_170 ();
 DECAPx2_ASAP7_75t_R FILLER_155_177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_183 ();
 FILLER_ASAP7_75t_R FILLER_155_226 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_257 ();
 DECAPx2_ASAP7_75t_R FILLER_155_289 ();
 FILLER_ASAP7_75t_R FILLER_155_301 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_306 ();
 DECAPx1_ASAP7_75t_R FILLER_155_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_339 ();
 DECAPx6_ASAP7_75t_R FILLER_155_346 ();
 DECAPx1_ASAP7_75t_R FILLER_155_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_364 ();
 DECAPx1_ASAP7_75t_R FILLER_155_371 ();
 DECAPx6_ASAP7_75t_R FILLER_155_381 ();
 DECAPx1_ASAP7_75t_R FILLER_155_395 ();
 DECAPx10_ASAP7_75t_R FILLER_155_402 ();
 FILLER_ASAP7_75t_R FILLER_155_424 ();
 DECAPx4_ASAP7_75t_R FILLER_155_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_439 ();
 DECAPx1_ASAP7_75t_R FILLER_155_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_470 ();
 DECAPx10_ASAP7_75t_R FILLER_155_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_517 ();
 DECAPx2_ASAP7_75t_R FILLER_155_535 ();
 DECAPx2_ASAP7_75t_R FILLER_155_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_553 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_564 ();
 DECAPx6_ASAP7_75t_R FILLER_155_582 ();
 FILLER_ASAP7_75t_R FILLER_155_596 ();
 DECAPx1_ASAP7_75t_R FILLER_155_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_611 ();
 FILLER_ASAP7_75t_R FILLER_155_619 ();
 DECAPx4_ASAP7_75t_R FILLER_155_629 ();
 FILLER_ASAP7_75t_R FILLER_155_639 ();
 DECAPx1_ASAP7_75t_R FILLER_155_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_675 ();
 DECAPx4_ASAP7_75t_R FILLER_155_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_695 ();
 FILLER_ASAP7_75t_R FILLER_155_714 ();
 DECAPx1_ASAP7_75t_R FILLER_155_719 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_782 ();
 DECAPx10_ASAP7_75t_R FILLER_155_800 ();
 DECAPx1_ASAP7_75t_R FILLER_155_822 ();
 DECAPx6_ASAP7_75t_R FILLER_155_839 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_853 ();
 DECAPx10_ASAP7_75t_R FILLER_155_862 ();
 DECAPx2_ASAP7_75t_R FILLER_155_884 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_155_890 ();
 FILLER_ASAP7_75t_R FILLER_155_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_155_933 ();
 DECAPx10_ASAP7_75t_R FILLER_156_2 ();
 DECAPx10_ASAP7_75t_R FILLER_156_24 ();
 DECAPx10_ASAP7_75t_R FILLER_156_46 ();
 DECAPx4_ASAP7_75t_R FILLER_156_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_128 ();
 DECAPx2_ASAP7_75t_R FILLER_156_158 ();
 FILLER_ASAP7_75t_R FILLER_156_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_226 ();
 DECAPx1_ASAP7_75t_R FILLER_156_235 ();
 DECAPx1_ASAP7_75t_R FILLER_156_248 ();
 DECAPx1_ASAP7_75t_R FILLER_156_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_268 ();
 FILLER_ASAP7_75t_R FILLER_156_286 ();
 FILLER_ASAP7_75t_R FILLER_156_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_334 ();
 DECAPx1_ASAP7_75t_R FILLER_156_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_345 ();
 DECAPx4_ASAP7_75t_R FILLER_156_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_362 ();
 FILLER_ASAP7_75t_R FILLER_156_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_383 ();
 DECAPx2_ASAP7_75t_R FILLER_156_413 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_419 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_435 ();
 FILLER_ASAP7_75t_R FILLER_156_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_461 ();
 DECAPx1_ASAP7_75t_R FILLER_156_464 ();
 DECAPx6_ASAP7_75t_R FILLER_156_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_503 ();
 DECAPx1_ASAP7_75t_R FILLER_156_549 ();
 FILLER_ASAP7_75t_R FILLER_156_570 ();
 DECAPx4_ASAP7_75t_R FILLER_156_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_590 ();
 DECAPx4_ASAP7_75t_R FILLER_156_619 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_629 ();
 DECAPx1_ASAP7_75t_R FILLER_156_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_644 ();
 FILLER_ASAP7_75t_R FILLER_156_674 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_685 ();
 DECAPx1_ASAP7_75t_R FILLER_156_700 ();
 DECAPx4_ASAP7_75t_R FILLER_156_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_753 ();
 DECAPx6_ASAP7_75t_R FILLER_156_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_781 ();
 DECAPx10_ASAP7_75t_R FILLER_156_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_156_819 ();
 DECAPx10_ASAP7_75t_R FILLER_156_846 ();
 DECAPx4_ASAP7_75t_R FILLER_156_868 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_156_878 ();
 DECAPx10_ASAP7_75t_R FILLER_157_2 ();
 DECAPx10_ASAP7_75t_R FILLER_157_24 ();
 DECAPx10_ASAP7_75t_R FILLER_157_46 ();
 DECAPx4_ASAP7_75t_R FILLER_157_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_144 ();
 FILLER_ASAP7_75t_R FILLER_157_175 ();
 DECAPx6_ASAP7_75t_R FILLER_157_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_201 ();
 DECAPx2_ASAP7_75t_R FILLER_157_208 ();
 DECAPx6_ASAP7_75t_R FILLER_157_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_231 ();
 DECAPx10_ASAP7_75t_R FILLER_157_246 ();
 DECAPx1_ASAP7_75t_R FILLER_157_268 ();
 FILLER_ASAP7_75t_R FILLER_157_280 ();
 DECAPx1_ASAP7_75t_R FILLER_157_288 ();
 DECAPx1_ASAP7_75t_R FILLER_157_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_349 ();
 DECAPx1_ASAP7_75t_R FILLER_157_457 ();
 DECAPx2_ASAP7_75t_R FILLER_157_469 ();
 DECAPx4_ASAP7_75t_R FILLER_157_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_518 ();
 DECAPx1_ASAP7_75t_R FILLER_157_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_526 ();
 FILLER_ASAP7_75t_R FILLER_157_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_556 ();
 DECAPx10_ASAP7_75t_R FILLER_157_565 ();
 DECAPx2_ASAP7_75t_R FILLER_157_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_593 ();
 DECAPx6_ASAP7_75t_R FILLER_157_604 ();
 DECAPx6_ASAP7_75t_R FILLER_157_624 ();
 DECAPx2_ASAP7_75t_R FILLER_157_638 ();
 DECAPx4_ASAP7_75t_R FILLER_157_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_663 ();
 DECAPx6_ASAP7_75t_R FILLER_157_670 ();
 DECAPx2_ASAP7_75t_R FILLER_157_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_690 ();
 DECAPx4_ASAP7_75t_R FILLER_157_702 ();
 DECAPx10_ASAP7_75t_R FILLER_157_721 ();
 DECAPx2_ASAP7_75t_R FILLER_157_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_749 ();
 DECAPx10_ASAP7_75t_R FILLER_157_761 ();
 DECAPx10_ASAP7_75t_R FILLER_157_783 ();
 FILLER_ASAP7_75t_R FILLER_157_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_837 ();
 DECAPx2_ASAP7_75t_R FILLER_157_848 ();
 FILLER_ASAP7_75t_R FILLER_157_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_157_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_157_924 ();
 FILLER_ASAP7_75t_R FILLER_157_932 ();
 DECAPx10_ASAP7_75t_R FILLER_158_2 ();
 DECAPx10_ASAP7_75t_R FILLER_158_24 ();
 DECAPx10_ASAP7_75t_R FILLER_158_46 ();
 DECAPx10_ASAP7_75t_R FILLER_158_68 ();
 DECAPx1_ASAP7_75t_R FILLER_158_90 ();
 DECAPx2_ASAP7_75t_R FILLER_158_97 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_103 ();
 DECAPx2_ASAP7_75t_R FILLER_158_125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_131 ();
 DECAPx2_ASAP7_75t_R FILLER_158_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_152 ();
 DECAPx10_ASAP7_75t_R FILLER_158_171 ();
 DECAPx10_ASAP7_75t_R FILLER_158_193 ();
 DECAPx6_ASAP7_75t_R FILLER_158_215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_229 ();
 DECAPx6_ASAP7_75t_R FILLER_158_258 ();
 DECAPx1_ASAP7_75t_R FILLER_158_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_276 ();
 DECAPx6_ASAP7_75t_R FILLER_158_283 ();
 DECAPx1_ASAP7_75t_R FILLER_158_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_301 ();
 DECAPx1_ASAP7_75t_R FILLER_158_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_329 ();
 FILLER_ASAP7_75t_R FILLER_158_336 ();
 DECAPx2_ASAP7_75t_R FILLER_158_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_347 ();
 DECAPx1_ASAP7_75t_R FILLER_158_356 ();
 FILLER_ASAP7_75t_R FILLER_158_366 ();
 FILLER_ASAP7_75t_R FILLER_158_411 ();
 DECAPx6_ASAP7_75t_R FILLER_158_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_461 ();
 FILLER_ASAP7_75t_R FILLER_158_464 ();
 DECAPx10_ASAP7_75t_R FILLER_158_472 ();
 DECAPx1_ASAP7_75t_R FILLER_158_494 ();
 DECAPx10_ASAP7_75t_R FILLER_158_504 ();
 DECAPx10_ASAP7_75t_R FILLER_158_526 ();
 DECAPx10_ASAP7_75t_R FILLER_158_548 ();
 DECAPx6_ASAP7_75t_R FILLER_158_570 ();
 DECAPx2_ASAP7_75t_R FILLER_158_584 ();
 DECAPx6_ASAP7_75t_R FILLER_158_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_610 ();
 DECAPx10_ASAP7_75t_R FILLER_158_618 ();
 DECAPx10_ASAP7_75t_R FILLER_158_640 ();
 DECAPx10_ASAP7_75t_R FILLER_158_662 ();
 DECAPx10_ASAP7_75t_R FILLER_158_684 ();
 DECAPx6_ASAP7_75t_R FILLER_158_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_720 ();
 DECAPx6_ASAP7_75t_R FILLER_158_739 ();
 DECAPx1_ASAP7_75t_R FILLER_158_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_158_801 ();
 DECAPx1_ASAP7_75t_R FILLER_158_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_158_920 ();
 DECAPx10_ASAP7_75t_R FILLER_159_2 ();
 DECAPx10_ASAP7_75t_R FILLER_159_24 ();
 DECAPx10_ASAP7_75t_R FILLER_159_46 ();
 DECAPx10_ASAP7_75t_R FILLER_159_68 ();
 DECAPx6_ASAP7_75t_R FILLER_159_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_104 ();
 DECAPx4_ASAP7_75t_R FILLER_159_112 ();
 FILLER_ASAP7_75t_R FILLER_159_122 ();
 DECAPx2_ASAP7_75t_R FILLER_159_153 ();
 FILLER_ASAP7_75t_R FILLER_159_159 ();
 DECAPx6_ASAP7_75t_R FILLER_159_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_181 ();
 DECAPx4_ASAP7_75t_R FILLER_159_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_200 ();
 DECAPx10_ASAP7_75t_R FILLER_159_207 ();
 DECAPx6_ASAP7_75t_R FILLER_159_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_243 ();
 DECAPx10_ASAP7_75t_R FILLER_159_269 ();
 DECAPx4_ASAP7_75t_R FILLER_159_291 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_301 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_312 ();
 DECAPx1_ASAP7_75t_R FILLER_159_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_345 ();
 DECAPx10_ASAP7_75t_R FILLER_159_358 ();
 DECAPx1_ASAP7_75t_R FILLER_159_380 ();
 DECAPx6_ASAP7_75t_R FILLER_159_390 ();
 FILLER_ASAP7_75t_R FILLER_159_404 ();
 DECAPx6_ASAP7_75t_R FILLER_159_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_423 ();
 DECAPx10_ASAP7_75t_R FILLER_159_437 ();
 DECAPx2_ASAP7_75t_R FILLER_159_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_465 ();
 DECAPx2_ASAP7_75t_R FILLER_159_479 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_485 ();
 DECAPx6_ASAP7_75t_R FILLER_159_495 ();
 DECAPx2_ASAP7_75t_R FILLER_159_509 ();
 DECAPx6_ASAP7_75t_R FILLER_159_529 ();
 FILLER_ASAP7_75t_R FILLER_159_551 ();
 DECAPx4_ASAP7_75t_R FILLER_159_556 ();
 FILLER_ASAP7_75t_R FILLER_159_566 ();
 DECAPx2_ASAP7_75t_R FILLER_159_574 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_580 ();
 DECAPx6_ASAP7_75t_R FILLER_159_590 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_604 ();
 DECAPx1_ASAP7_75t_R FILLER_159_613 ();
 DECAPx10_ASAP7_75t_R FILLER_159_639 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_661 ();
 DECAPx10_ASAP7_75t_R FILLER_159_670 ();
 DECAPx2_ASAP7_75t_R FILLER_159_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_698 ();
 DECAPx2_ASAP7_75t_R FILLER_159_709 ();
 FILLER_ASAP7_75t_R FILLER_159_715 ();
 DECAPx2_ASAP7_75t_R FILLER_159_763 ();
 FILLER_ASAP7_75t_R FILLER_159_769 ();
 DECAPx1_ASAP7_75t_R FILLER_159_803 ();
 DECAPx10_ASAP7_75t_R FILLER_159_826 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_159_848 ();
 DECAPx1_ASAP7_75t_R FILLER_159_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_159_861 ();
 DECAPx10_ASAP7_75t_R FILLER_159_865 ();
 DECAPx2_ASAP7_75t_R FILLER_159_887 ();
 DECAPx10_ASAP7_75t_R FILLER_160_2 ();
 DECAPx10_ASAP7_75t_R FILLER_160_24 ();
 DECAPx10_ASAP7_75t_R FILLER_160_46 ();
 DECAPx10_ASAP7_75t_R FILLER_160_68 ();
 DECAPx10_ASAP7_75t_R FILLER_160_90 ();
 DECAPx2_ASAP7_75t_R FILLER_160_118 ();
 DECAPx2_ASAP7_75t_R FILLER_160_130 ();
 FILLER_ASAP7_75t_R FILLER_160_136 ();
 DECAPx10_ASAP7_75t_R FILLER_160_141 ();
 DECAPx6_ASAP7_75t_R FILLER_160_163 ();
 FILLER_ASAP7_75t_R FILLER_160_177 ();
 DECAPx10_ASAP7_75t_R FILLER_160_217 ();
 DECAPx6_ASAP7_75t_R FILLER_160_239 ();
 DECAPx2_ASAP7_75t_R FILLER_160_253 ();
 DECAPx1_ASAP7_75t_R FILLER_160_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_269 ();
 DECAPx1_ASAP7_75t_R FILLER_160_281 ();
 DECAPx1_ASAP7_75t_R FILLER_160_303 ();
 DECAPx10_ASAP7_75t_R FILLER_160_345 ();
 DECAPx4_ASAP7_75t_R FILLER_160_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_377 ();
 DECAPx10_ASAP7_75t_R FILLER_160_404 ();
 DECAPx6_ASAP7_75t_R FILLER_160_426 ();
 DECAPx2_ASAP7_75t_R FILLER_160_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_446 ();
 DECAPx2_ASAP7_75t_R FILLER_160_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_484 ();
 DECAPx6_ASAP7_75t_R FILLER_160_504 ();
 DECAPx2_ASAP7_75t_R FILLER_160_529 ();
 FILLER_ASAP7_75t_R FILLER_160_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_563 ();
 DECAPx1_ASAP7_75t_R FILLER_160_567 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_584 ();
 DECAPx10_ASAP7_75t_R FILLER_160_598 ();
 DECAPx10_ASAP7_75t_R FILLER_160_620 ();
 DECAPx2_ASAP7_75t_R FILLER_160_642 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_662 ();
 FILLER_ASAP7_75t_R FILLER_160_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_160_696 ();
 DECAPx2_ASAP7_75t_R FILLER_160_708 ();
 FILLER_ASAP7_75t_R FILLER_160_748 ();
 FILLER_ASAP7_75t_R FILLER_160_795 ();
 DECAPx10_ASAP7_75t_R FILLER_160_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_160_825 ();
 DECAPx10_ASAP7_75t_R FILLER_160_836 ();
 DECAPx4_ASAP7_75t_R FILLER_160_858 ();
 DECAPx1_ASAP7_75t_R FILLER_160_894 ();
 DECAPx10_ASAP7_75t_R FILLER_161_2 ();
 DECAPx10_ASAP7_75t_R FILLER_161_24 ();
 DECAPx10_ASAP7_75t_R FILLER_161_46 ();
 DECAPx4_ASAP7_75t_R FILLER_161_68 ();
 FILLER_ASAP7_75t_R FILLER_161_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_95 ();
 DECAPx2_ASAP7_75t_R FILLER_161_104 ();
 DECAPx2_ASAP7_75t_R FILLER_161_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_122 ();
 DECAPx10_ASAP7_75t_R FILLER_161_129 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_151 ();
 DECAPx4_ASAP7_75t_R FILLER_161_184 ();
 FILLER_ASAP7_75t_R FILLER_161_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_202 ();
 FILLER_ASAP7_75t_R FILLER_161_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_308 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_326 ();
 DECAPx2_ASAP7_75t_R FILLER_161_353 ();
 FILLER_ASAP7_75t_R FILLER_161_359 ();
 DECAPx6_ASAP7_75t_R FILLER_161_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_381 ();
 DECAPx4_ASAP7_75t_R FILLER_161_407 ();
 FILLER_ASAP7_75t_R FILLER_161_417 ();
 DECAPx10_ASAP7_75t_R FILLER_161_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_485 ();
 DECAPx2_ASAP7_75t_R FILLER_161_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_510 ();
 DECAPx1_ASAP7_75t_R FILLER_161_537 ();
 FILLER_ASAP7_75t_R FILLER_161_556 ();
 DECAPx1_ASAP7_75t_R FILLER_161_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_590 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_603 ();
 DECAPx4_ASAP7_75t_R FILLER_161_613 ();
 DECAPx2_ASAP7_75t_R FILLER_161_646 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_161_652 ();
 DECAPx2_ASAP7_75t_R FILLER_161_667 ();
 FILLER_ASAP7_75t_R FILLER_161_673 ();
 DECAPx6_ASAP7_75t_R FILLER_161_712 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_766 ();
 DECAPx2_ASAP7_75t_R FILLER_161_776 ();
 DECAPx1_ASAP7_75t_R FILLER_161_793 ();
 DECAPx6_ASAP7_75t_R FILLER_161_802 ();
 FILLER_ASAP7_75t_R FILLER_161_816 ();
 DECAPx10_ASAP7_75t_R FILLER_161_844 ();
 FILLER_ASAP7_75t_R FILLER_161_866 ();
 FILLER_ASAP7_75t_R FILLER_161_883 ();
 FILLER_ASAP7_75t_R FILLER_161_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_161_921 ();
 FILLER_ASAP7_75t_R FILLER_161_927 ();
 DECAPx10_ASAP7_75t_R FILLER_162_2 ();
 DECAPx10_ASAP7_75t_R FILLER_162_24 ();
 DECAPx10_ASAP7_75t_R FILLER_162_46 ();
 DECAPx2_ASAP7_75t_R FILLER_162_68 ();
 FILLER_ASAP7_75t_R FILLER_162_74 ();
 DECAPx10_ASAP7_75t_R FILLER_162_124 ();
 DECAPx2_ASAP7_75t_R FILLER_162_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_197 ();
 FILLER_ASAP7_75t_R FILLER_162_204 ();
 DECAPx2_ASAP7_75t_R FILLER_162_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_258 ();
 DECAPx10_ASAP7_75t_R FILLER_162_279 ();
 DECAPx10_ASAP7_75t_R FILLER_162_301 ();
 DECAPx6_ASAP7_75t_R FILLER_162_323 ();
 DECAPx1_ASAP7_75t_R FILLER_162_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_341 ();
 FILLER_ASAP7_75t_R FILLER_162_345 ();
 DECAPx4_ASAP7_75t_R FILLER_162_379 ();
 FILLER_ASAP7_75t_R FILLER_162_389 ();
 DECAPx2_ASAP7_75t_R FILLER_162_397 ();
 FILLER_ASAP7_75t_R FILLER_162_403 ();
 FILLER_ASAP7_75t_R FILLER_162_472 ();
 DECAPx1_ASAP7_75t_R FILLER_162_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_492 ();
 DECAPx10_ASAP7_75t_R FILLER_162_519 ();
 DECAPx10_ASAP7_75t_R FILLER_162_541 ();
 DECAPx10_ASAP7_75t_R FILLER_162_563 ();
 DECAPx1_ASAP7_75t_R FILLER_162_585 ();
 DECAPx1_ASAP7_75t_R FILLER_162_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_607 ();
 FILLER_ASAP7_75t_R FILLER_162_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_643 ();
 DECAPx4_ASAP7_75t_R FILLER_162_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_665 ();
 DECAPx1_ASAP7_75t_R FILLER_162_672 ();
 DECAPx2_ASAP7_75t_R FILLER_162_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_688 ();
 DECAPx1_ASAP7_75t_R FILLER_162_697 ();
 DECAPx10_ASAP7_75t_R FILLER_162_707 ();
 DECAPx1_ASAP7_75t_R FILLER_162_729 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_733 ();
 DECAPx6_ASAP7_75t_R FILLER_162_739 ();
 DECAPx2_ASAP7_75t_R FILLER_162_753 ();
 DECAPx4_ASAP7_75t_R FILLER_162_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_162_777 ();
 FILLER_ASAP7_75t_R FILLER_162_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_832 ();
 DECAPx2_ASAP7_75t_R FILLER_162_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_842 ();
 FILLER_ASAP7_75t_R FILLER_162_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_881 ();
 DECAPx1_ASAP7_75t_R FILLER_162_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_162_903 ();
 DECAPx10_ASAP7_75t_R FILLER_163_2 ();
 DECAPx10_ASAP7_75t_R FILLER_163_24 ();
 DECAPx10_ASAP7_75t_R FILLER_163_46 ();
 DECAPx6_ASAP7_75t_R FILLER_163_68 ();
 DECAPx1_ASAP7_75t_R FILLER_163_94 ();
 DECAPx2_ASAP7_75t_R FILLER_163_104 ();
 FILLER_ASAP7_75t_R FILLER_163_110 ();
 FILLER_ASAP7_75t_R FILLER_163_138 ();
 DECAPx2_ASAP7_75t_R FILLER_163_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_160 ();
 FILLER_ASAP7_75t_R FILLER_163_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_216 ();
 DECAPx10_ASAP7_75t_R FILLER_163_236 ();
 DECAPx4_ASAP7_75t_R FILLER_163_258 ();
 DECAPx2_ASAP7_75t_R FILLER_163_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_283 ();
 DECAPx10_ASAP7_75t_R FILLER_163_292 ();
 FILLER_ASAP7_75t_R FILLER_163_314 ();
 DECAPx10_ASAP7_75t_R FILLER_163_328 ();
 DECAPx2_ASAP7_75t_R FILLER_163_350 ();
 FILLER_ASAP7_75t_R FILLER_163_356 ();
 DECAPx4_ASAP7_75t_R FILLER_163_390 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_400 ();
 FILLER_ASAP7_75t_R FILLER_163_419 ();
 DECAPx10_ASAP7_75t_R FILLER_163_468 ();
 DECAPx4_ASAP7_75t_R FILLER_163_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_500 ();
 DECAPx6_ASAP7_75t_R FILLER_163_510 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_524 ();
 DECAPx10_ASAP7_75t_R FILLER_163_539 ();
 DECAPx4_ASAP7_75t_R FILLER_163_561 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_571 ();
 DECAPx4_ASAP7_75t_R FILLER_163_588 ();
 DECAPx1_ASAP7_75t_R FILLER_163_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_608 ();
 DECAPx1_ASAP7_75t_R FILLER_163_621 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_163_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_644 ();
 DECAPx10_ASAP7_75t_R FILLER_163_669 ();
 DECAPx6_ASAP7_75t_R FILLER_163_691 ();
 DECAPx10_ASAP7_75t_R FILLER_163_734 ();
 DECAPx10_ASAP7_75t_R FILLER_163_756 ();
 DECAPx4_ASAP7_75t_R FILLER_163_778 ();
 DECAPx4_ASAP7_75t_R FILLER_163_823 ();
 DECAPx1_ASAP7_75t_R FILLER_163_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_163_907 ();
 FILLER_ASAP7_75t_R FILLER_163_927 ();
 DECAPx10_ASAP7_75t_R FILLER_164_2 ();
 DECAPx10_ASAP7_75t_R FILLER_164_24 ();
 DECAPx10_ASAP7_75t_R FILLER_164_46 ();
 DECAPx2_ASAP7_75t_R FILLER_164_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_74 ();
 DECAPx6_ASAP7_75t_R FILLER_164_106 ();
 DECAPx1_ASAP7_75t_R FILLER_164_163 ();
 DECAPx10_ASAP7_75t_R FILLER_164_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_192 ();
 DECAPx10_ASAP7_75t_R FILLER_164_215 ();
 DECAPx10_ASAP7_75t_R FILLER_164_237 ();
 DECAPx10_ASAP7_75t_R FILLER_164_259 ();
 DECAPx2_ASAP7_75t_R FILLER_164_310 ();
 DECAPx1_ASAP7_75t_R FILLER_164_324 ();
 DECAPx4_ASAP7_75t_R FILLER_164_354 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_364 ();
 DECAPx2_ASAP7_75t_R FILLER_164_380 ();
 FILLER_ASAP7_75t_R FILLER_164_402 ();
 DECAPx2_ASAP7_75t_R FILLER_164_410 ();
 FILLER_ASAP7_75t_R FILLER_164_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_435 ();
 DECAPx1_ASAP7_75t_R FILLER_164_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_443 ();
 DECAPx4_ASAP7_75t_R FILLER_164_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_461 ();
 DECAPx4_ASAP7_75t_R FILLER_164_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_474 ();
 DECAPx2_ASAP7_75t_R FILLER_164_490 ();
 DECAPx2_ASAP7_75t_R FILLER_164_502 ();
 FILLER_ASAP7_75t_R FILLER_164_508 ();
 DECAPx4_ASAP7_75t_R FILLER_164_542 ();
 DECAPx10_ASAP7_75t_R FILLER_164_564 ();
 DECAPx10_ASAP7_75t_R FILLER_164_586 ();
 DECAPx10_ASAP7_75t_R FILLER_164_608 ();
 DECAPx1_ASAP7_75t_R FILLER_164_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_634 ();
 DECAPx10_ASAP7_75t_R FILLER_164_656 ();
 DECAPx10_ASAP7_75t_R FILLER_164_678 ();
 DECAPx4_ASAP7_75t_R FILLER_164_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_164_710 ();
 DECAPx6_ASAP7_75t_R FILLER_164_739 ();
 DECAPx2_ASAP7_75t_R FILLER_164_753 ();
 DECAPx10_ASAP7_75t_R FILLER_164_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_814 ();
 DECAPx2_ASAP7_75t_R FILLER_164_818 ();
 DECAPx4_ASAP7_75t_R FILLER_164_834 ();
 FILLER_ASAP7_75t_R FILLER_164_853 ();
 FILLERxp5_ASAP7_75t_R FILLER_164_887 ();
 DECAPx10_ASAP7_75t_R FILLER_165_2 ();
 DECAPx10_ASAP7_75t_R FILLER_165_24 ();
 DECAPx10_ASAP7_75t_R FILLER_165_46 ();
 DECAPx10_ASAP7_75t_R FILLER_165_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_90 ();
 DECAPx10_ASAP7_75t_R FILLER_165_94 ();
 DECAPx6_ASAP7_75t_R FILLER_165_116 ();
 DECAPx2_ASAP7_75t_R FILLER_165_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_142 ();
 DECAPx1_ASAP7_75t_R FILLER_165_146 ();
 DECAPx4_ASAP7_75t_R FILLER_165_153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_172 ();
 DECAPx6_ASAP7_75t_R FILLER_165_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_193 ();
 DECAPx10_ASAP7_75t_R FILLER_165_211 ();
 DECAPx1_ASAP7_75t_R FILLER_165_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_237 ();
 FILLER_ASAP7_75t_R FILLER_165_260 ();
 FILLER_ASAP7_75t_R FILLER_165_268 ();
 DECAPx1_ASAP7_75t_R FILLER_165_285 ();
 DECAPx2_ASAP7_75t_R FILLER_165_298 ();
 FILLER_ASAP7_75t_R FILLER_165_304 ();
 DECAPx1_ASAP7_75t_R FILLER_165_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_316 ();
 DECAPx10_ASAP7_75t_R FILLER_165_361 ();
 DECAPx2_ASAP7_75t_R FILLER_165_383 ();
 DECAPx10_ASAP7_75t_R FILLER_165_402 ();
 DECAPx10_ASAP7_75t_R FILLER_165_424 ();
 DECAPx6_ASAP7_75t_R FILLER_165_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_460 ();
 DECAPx10_ASAP7_75t_R FILLER_165_477 ();
 DECAPx10_ASAP7_75t_R FILLER_165_499 ();
 DECAPx4_ASAP7_75t_R FILLER_165_521 ();
 FILLER_ASAP7_75t_R FILLER_165_537 ();
 DECAPx6_ASAP7_75t_R FILLER_165_575 ();
 DECAPx2_ASAP7_75t_R FILLER_165_600 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_606 ();
 DECAPx6_ASAP7_75t_R FILLER_165_620 ();
 DECAPx2_ASAP7_75t_R FILLER_165_634 ();
 DECAPx6_ASAP7_75t_R FILLER_165_646 ();
 DECAPx1_ASAP7_75t_R FILLER_165_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_664 ();
 FILLER_ASAP7_75t_R FILLER_165_670 ();
 DECAPx4_ASAP7_75t_R FILLER_165_687 ();
 DECAPx2_ASAP7_75t_R FILLER_165_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_731 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_165_754 ();
 DECAPx10_ASAP7_75t_R FILLER_165_783 ();
 DECAPx4_ASAP7_75t_R FILLER_165_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_815 ();
 DECAPx10_ASAP7_75t_R FILLER_165_842 ();
 DECAPx6_ASAP7_75t_R FILLER_165_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_165_924 ();
 FILLER_ASAP7_75t_R FILLER_165_932 ();
 DECAPx10_ASAP7_75t_R FILLER_166_2 ();
 DECAPx10_ASAP7_75t_R FILLER_166_24 ();
 DECAPx10_ASAP7_75t_R FILLER_166_46 ();
 DECAPx10_ASAP7_75t_R FILLER_166_68 ();
 DECAPx6_ASAP7_75t_R FILLER_166_90 ();
 DECAPx1_ASAP7_75t_R FILLER_166_104 ();
 DECAPx10_ASAP7_75t_R FILLER_166_123 ();
 DECAPx1_ASAP7_75t_R FILLER_166_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_161 ();
 DECAPx2_ASAP7_75t_R FILLER_166_188 ();
 DECAPx2_ASAP7_75t_R FILLER_166_220 ();
 FILLER_ASAP7_75t_R FILLER_166_226 ();
 FILLER_ASAP7_75t_R FILLER_166_234 ();
 DECAPx6_ASAP7_75t_R FILLER_166_280 ();
 DECAPx1_ASAP7_75t_R FILLER_166_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_298 ();
 FILLER_ASAP7_75t_R FILLER_166_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_354 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_361 ();
 DECAPx6_ASAP7_75t_R FILLER_166_367 ();
 DECAPx2_ASAP7_75t_R FILLER_166_381 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_387 ();
 DECAPx2_ASAP7_75t_R FILLER_166_418 ();
 DECAPx2_ASAP7_75t_R FILLER_166_434 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_472 ();
 DECAPx4_ASAP7_75t_R FILLER_166_483 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_493 ();
 DECAPx10_ASAP7_75t_R FILLER_166_504 ();
 DECAPx4_ASAP7_75t_R FILLER_166_526 ();
 DECAPx4_ASAP7_75t_R FILLER_166_584 ();
 DECAPx2_ASAP7_75t_R FILLER_166_602 ();
 DECAPx2_ASAP7_75t_R FILLER_166_614 ();
 DECAPx6_ASAP7_75t_R FILLER_166_638 ();
 DECAPx1_ASAP7_75t_R FILLER_166_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_686 ();
 DECAPx6_ASAP7_75t_R FILLER_166_695 ();
 FILLER_ASAP7_75t_R FILLER_166_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_717 ();
 DECAPx1_ASAP7_75t_R FILLER_166_744 ();
 DECAPx10_ASAP7_75t_R FILLER_166_800 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_822 ();
 DECAPx10_ASAP7_75t_R FILLER_166_836 ();
 DECAPx6_ASAP7_75t_R FILLER_166_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_166_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_166_918 ();
 DECAPx10_ASAP7_75t_R FILLER_167_2 ();
 DECAPx10_ASAP7_75t_R FILLER_167_24 ();
 DECAPx10_ASAP7_75t_R FILLER_167_46 ();
 DECAPx6_ASAP7_75t_R FILLER_167_68 ();
 FILLER_ASAP7_75t_R FILLER_167_82 ();
 DECAPx6_ASAP7_75t_R FILLER_167_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_104 ();
 DECAPx6_ASAP7_75t_R FILLER_167_131 ();
 DECAPx10_ASAP7_75t_R FILLER_167_151 ();
 FILLER_ASAP7_75t_R FILLER_167_173 ();
 DECAPx10_ASAP7_75t_R FILLER_167_185 ();
 FILLER_ASAP7_75t_R FILLER_167_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_212 ();
 FILLER_ASAP7_75t_R FILLER_167_223 ();
 DECAPx2_ASAP7_75t_R FILLER_167_251 ();
 DECAPx2_ASAP7_75t_R FILLER_167_263 ();
 DECAPx6_ASAP7_75t_R FILLER_167_272 ();
 FILLER_ASAP7_75t_R FILLER_167_286 ();
 FILLER_ASAP7_75t_R FILLER_167_308 ();
 DECAPx10_ASAP7_75t_R FILLER_167_317 ();
 DECAPx6_ASAP7_75t_R FILLER_167_339 ();
 DECAPx2_ASAP7_75t_R FILLER_167_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_392 ();
 FILLER_ASAP7_75t_R FILLER_167_411 ();
 DECAPx2_ASAP7_75t_R FILLER_167_448 ();
 DECAPx1_ASAP7_75t_R FILLER_167_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_484 ();
 DECAPx1_ASAP7_75t_R FILLER_167_518 ();
 DECAPx10_ASAP7_75t_R FILLER_167_532 ();
 DECAPx4_ASAP7_75t_R FILLER_167_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_564 ();
 FILLER_ASAP7_75t_R FILLER_167_574 ();
 FILLER_ASAP7_75t_R FILLER_167_594 ();
 DECAPx4_ASAP7_75t_R FILLER_167_613 ();
 FILLER_ASAP7_75t_R FILLER_167_623 ();
 DECAPx6_ASAP7_75t_R FILLER_167_633 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_167_647 ();
 DECAPx6_ASAP7_75t_R FILLER_167_659 ();
 DECAPx1_ASAP7_75t_R FILLER_167_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_684 ();
 DECAPx10_ASAP7_75t_R FILLER_167_714 ();
 DECAPx2_ASAP7_75t_R FILLER_167_755 ();
 FILLER_ASAP7_75t_R FILLER_167_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_786 ();
 DECAPx10_ASAP7_75t_R FILLER_167_790 ();
 DECAPx6_ASAP7_75t_R FILLER_167_812 ();
 DECAPx1_ASAP7_75t_R FILLER_167_832 ();
 DECAPx2_ASAP7_75t_R FILLER_167_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_167_919 ();
 FILLER_ASAP7_75t_R FILLER_167_927 ();
 DECAPx10_ASAP7_75t_R FILLER_168_2 ();
 DECAPx10_ASAP7_75t_R FILLER_168_24 ();
 DECAPx10_ASAP7_75t_R FILLER_168_46 ();
 DECAPx4_ASAP7_75t_R FILLER_168_68 ();
 FILLER_ASAP7_75t_R FILLER_168_78 ();
 DECAPx6_ASAP7_75t_R FILLER_168_106 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_126 ();
 FILLER_ASAP7_75t_R FILLER_168_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_160 ();
 FILLER_ASAP7_75t_R FILLER_168_189 ();
 DECAPx4_ASAP7_75t_R FILLER_168_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_210 ();
 DECAPx10_ASAP7_75t_R FILLER_168_242 ();
 DECAPx6_ASAP7_75t_R FILLER_168_264 ();
 FILLER_ASAP7_75t_R FILLER_168_278 ();
 DECAPx6_ASAP7_75t_R FILLER_168_306 ();
 FILLER_ASAP7_75t_R FILLER_168_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_344 ();
 DECAPx1_ASAP7_75t_R FILLER_168_359 ();
 DECAPx1_ASAP7_75t_R FILLER_168_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_381 ();
 DECAPx2_ASAP7_75t_R FILLER_168_388 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_394 ();
 FILLER_ASAP7_75t_R FILLER_168_432 ();
 DECAPx4_ASAP7_75t_R FILLER_168_450 ();
 FILLER_ASAP7_75t_R FILLER_168_460 ();
 DECAPx1_ASAP7_75t_R FILLER_168_464 ();
 DECAPx2_ASAP7_75t_R FILLER_168_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_477 ();
 DECAPx1_ASAP7_75t_R FILLER_168_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_503 ();
 FILLER_ASAP7_75t_R FILLER_168_522 ();
 DECAPx1_ASAP7_75t_R FILLER_168_534 ();
 DECAPx10_ASAP7_75t_R FILLER_168_544 ();
 DECAPx1_ASAP7_75t_R FILLER_168_566 ();
 FILLER_ASAP7_75t_R FILLER_168_577 ();
 DECAPx1_ASAP7_75t_R FILLER_168_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_598 ();
 DECAPx10_ASAP7_75t_R FILLER_168_610 ();
 DECAPx1_ASAP7_75t_R FILLER_168_650 ();
 DECAPx2_ASAP7_75t_R FILLER_168_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_691 ();
 DECAPx10_ASAP7_75t_R FILLER_168_707 ();
 DECAPx10_ASAP7_75t_R FILLER_168_729 ();
 DECAPx10_ASAP7_75t_R FILLER_168_751 ();
 DECAPx2_ASAP7_75t_R FILLER_168_773 ();
 DECAPx2_ASAP7_75t_R FILLER_168_785 ();
 FILLER_ASAP7_75t_R FILLER_168_791 ();
 DECAPx2_ASAP7_75t_R FILLER_168_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_168_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_168_887 ();
 FILLER_ASAP7_75t_R FILLER_168_896 ();
 DECAPx10_ASAP7_75t_R FILLER_169_2 ();
 DECAPx10_ASAP7_75t_R FILLER_169_24 ();
 DECAPx10_ASAP7_75t_R FILLER_169_46 ();
 DECAPx6_ASAP7_75t_R FILLER_169_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_94 ();
 FILLER_ASAP7_75t_R FILLER_169_104 ();
 DECAPx2_ASAP7_75t_R FILLER_169_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_139 ();
 FILLER_ASAP7_75t_R FILLER_169_146 ();
 DECAPx2_ASAP7_75t_R FILLER_169_151 ();
 DECAPx1_ASAP7_75t_R FILLER_169_209 ();
 DECAPx10_ASAP7_75t_R FILLER_169_223 ();
 DECAPx4_ASAP7_75t_R FILLER_169_245 ();
 FILLER_ASAP7_75t_R FILLER_169_255 ();
 DECAPx6_ASAP7_75t_R FILLER_169_263 ();
 DECAPx2_ASAP7_75t_R FILLER_169_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_283 ();
 DECAPx6_ASAP7_75t_R FILLER_169_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_332 ();
 FILLER_ASAP7_75t_R FILLER_169_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_409 ();
 DECAPx10_ASAP7_75t_R FILLER_169_444 ();
 DECAPx10_ASAP7_75t_R FILLER_169_466 ();
 DECAPx4_ASAP7_75t_R FILLER_169_488 ();
 FILLER_ASAP7_75t_R FILLER_169_498 ();
 DECAPx4_ASAP7_75t_R FILLER_169_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_526 ();
 DECAPx10_ASAP7_75t_R FILLER_169_535 ();
 DECAPx10_ASAP7_75t_R FILLER_169_557 ();
 DECAPx4_ASAP7_75t_R FILLER_169_579 ();
 FILLER_ASAP7_75t_R FILLER_169_589 ();
 DECAPx6_ASAP7_75t_R FILLER_169_597 ();
 DECAPx2_ASAP7_75t_R FILLER_169_611 ();
 DECAPx6_ASAP7_75t_R FILLER_169_627 ();
 FILLER_ASAP7_75t_R FILLER_169_641 ();
 DECAPx1_ASAP7_75t_R FILLER_169_649 ();
 DECAPx10_ASAP7_75t_R FILLER_169_659 ();
 DECAPx1_ASAP7_75t_R FILLER_169_681 ();
 DECAPx6_ASAP7_75t_R FILLER_169_689 ();
 FILLER_ASAP7_75t_R FILLER_169_703 ();
 FILLER_ASAP7_75t_R FILLER_169_724 ();
 DECAPx10_ASAP7_75t_R FILLER_169_731 ();
 FILLER_ASAP7_75t_R FILLER_169_753 ();
 DECAPx10_ASAP7_75t_R FILLER_169_758 ();
 FILLER_ASAP7_75t_R FILLER_169_780 ();
 FILLER_ASAP7_75t_R FILLER_169_798 ();
 DECAPx2_ASAP7_75t_R FILLER_169_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_835 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_169_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_169_921 ();
 FILLER_ASAP7_75t_R FILLER_169_932 ();
 DECAPx10_ASAP7_75t_R FILLER_170_2 ();
 DECAPx10_ASAP7_75t_R FILLER_170_24 ();
 DECAPx10_ASAP7_75t_R FILLER_170_46 ();
 DECAPx10_ASAP7_75t_R FILLER_170_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_90 ();
 DECAPx10_ASAP7_75t_R FILLER_170_117 ();
 DECAPx10_ASAP7_75t_R FILLER_170_139 ();
 DECAPx4_ASAP7_75t_R FILLER_170_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_195 ();
 DECAPx10_ASAP7_75t_R FILLER_170_227 ();
 DECAPx1_ASAP7_75t_R FILLER_170_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_253 ();
 DECAPx10_ASAP7_75t_R FILLER_170_283 ();
 DECAPx10_ASAP7_75t_R FILLER_170_305 ();
 FILLER_ASAP7_75t_R FILLER_170_327 ();
 FILLER_ASAP7_75t_R FILLER_170_363 ();
 DECAPx10_ASAP7_75t_R FILLER_170_371 ();
 DECAPx10_ASAP7_75t_R FILLER_170_393 ();
 DECAPx1_ASAP7_75t_R FILLER_170_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_419 ();
 DECAPx6_ASAP7_75t_R FILLER_170_430 ();
 DECAPx2_ASAP7_75t_R FILLER_170_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_450 ();
 DECAPx1_ASAP7_75t_R FILLER_170_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_464 ();
 DECAPx2_ASAP7_75t_R FILLER_170_474 ();
 DECAPx10_ASAP7_75t_R FILLER_170_489 ();
 DECAPx4_ASAP7_75t_R FILLER_170_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_538 ();
 FILLER_ASAP7_75t_R FILLER_170_547 ();
 FILLER_ASAP7_75t_R FILLER_170_552 ();
 DECAPx1_ASAP7_75t_R FILLER_170_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_570 ();
 DECAPx10_ASAP7_75t_R FILLER_170_578 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_600 ();
 DECAPx1_ASAP7_75t_R FILLER_170_612 ();
 DECAPx6_ASAP7_75t_R FILLER_170_622 ();
 FILLER_ASAP7_75t_R FILLER_170_636 ();
 DECAPx2_ASAP7_75t_R FILLER_170_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_664 ();
 DECAPx10_ASAP7_75t_R FILLER_170_671 ();
 DECAPx6_ASAP7_75t_R FILLER_170_693 ();
 DECAPx2_ASAP7_75t_R FILLER_170_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_739 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_170_766 ();
 DECAPx4_ASAP7_75t_R FILLER_170_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_787 ();
 DECAPx10_ASAP7_75t_R FILLER_170_828 ();
 DECAPx4_ASAP7_75t_R FILLER_170_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_874 ();
 FILLER_ASAP7_75t_R FILLER_170_891 ();
 FILLER_ASAP7_75t_R FILLER_170_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_170_928 ();
 DECAPx10_ASAP7_75t_R FILLER_171_2 ();
 DECAPx10_ASAP7_75t_R FILLER_171_24 ();
 DECAPx10_ASAP7_75t_R FILLER_171_46 ();
 DECAPx10_ASAP7_75t_R FILLER_171_68 ();
 DECAPx6_ASAP7_75t_R FILLER_171_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_104 ();
 DECAPx2_ASAP7_75t_R FILLER_171_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_117 ();
 DECAPx2_ASAP7_75t_R FILLER_171_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_141 ();
 DECAPx2_ASAP7_75t_R FILLER_171_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_154 ();
 DECAPx10_ASAP7_75t_R FILLER_171_163 ();
 DECAPx2_ASAP7_75t_R FILLER_171_185 ();
 DECAPx2_ASAP7_75t_R FILLER_171_197 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_251 ();
 FILLER_ASAP7_75t_R FILLER_171_287 ();
 DECAPx2_ASAP7_75t_R FILLER_171_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_301 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_324 ();
 DECAPx4_ASAP7_75t_R FILLER_171_333 ();
 DECAPx10_ASAP7_75t_R FILLER_171_352 ();
 DECAPx10_ASAP7_75t_R FILLER_171_374 ();
 DECAPx10_ASAP7_75t_R FILLER_171_396 ();
 DECAPx4_ASAP7_75t_R FILLER_171_418 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_437 ();
 DECAPx1_ASAP7_75t_R FILLER_171_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_454 ();
 FILLER_ASAP7_75t_R FILLER_171_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_493 ();
 DECAPx10_ASAP7_75t_R FILLER_171_506 ();
 FILLER_ASAP7_75t_R FILLER_171_572 ();
 DECAPx6_ASAP7_75t_R FILLER_171_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_598 ();
 FILLER_ASAP7_75t_R FILLER_171_626 ();
 DECAPx6_ASAP7_75t_R FILLER_171_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_648 ();
 DECAPx2_ASAP7_75t_R FILLER_171_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_658 ();
 DECAPx4_ASAP7_75t_R FILLER_171_680 ();
 DECAPx6_ASAP7_75t_R FILLER_171_696 ();
 DECAPx2_ASAP7_75t_R FILLER_171_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_716 ();
 DECAPx1_ASAP7_75t_R FILLER_171_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_767 ();
 DECAPx10_ASAP7_75t_R FILLER_171_794 ();
 DECAPx1_ASAP7_75t_R FILLER_171_819 ();
 DECAPx6_ASAP7_75t_R FILLER_171_829 ();
 DECAPx2_ASAP7_75t_R FILLER_171_843 ();
 DECAPx4_ASAP7_75t_R FILLER_171_856 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_171_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_171_933 ();
 DECAPx10_ASAP7_75t_R FILLER_172_2 ();
 DECAPx10_ASAP7_75t_R FILLER_172_24 ();
 DECAPx10_ASAP7_75t_R FILLER_172_46 ();
 DECAPx6_ASAP7_75t_R FILLER_172_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_82 ();
 DECAPx1_ASAP7_75t_R FILLER_172_91 ();
 DECAPx4_ASAP7_75t_R FILLER_172_101 ();
 FILLER_ASAP7_75t_R FILLER_172_111 ();
 FILLER_ASAP7_75t_R FILLER_172_119 ();
 DECAPx2_ASAP7_75t_R FILLER_172_129 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_146 ();
 DECAPx2_ASAP7_75t_R FILLER_172_173 ();
 FILLER_ASAP7_75t_R FILLER_172_179 ();
 DECAPx4_ASAP7_75t_R FILLER_172_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_217 ();
 DECAPx2_ASAP7_75t_R FILLER_172_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_303 ();
 DECAPx6_ASAP7_75t_R FILLER_172_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_335 ();
 DECAPx1_ASAP7_75t_R FILLER_172_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_346 ();
 DECAPx2_ASAP7_75t_R FILLER_172_350 ();
 FILLER_ASAP7_75t_R FILLER_172_382 ();
 DECAPx2_ASAP7_75t_R FILLER_172_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_399 ();
 DECAPx2_ASAP7_75t_R FILLER_172_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_414 ();
 DECAPx6_ASAP7_75t_R FILLER_172_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_461 ();
 DECAPx1_ASAP7_75t_R FILLER_172_504 ();
 DECAPx1_ASAP7_75t_R FILLER_172_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_520 ();
 DECAPx1_ASAP7_75t_R FILLER_172_538 ();
 DECAPx2_ASAP7_75t_R FILLER_172_550 ();
 FILLER_ASAP7_75t_R FILLER_172_556 ();
 DECAPx2_ASAP7_75t_R FILLER_172_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_570 ();
 DECAPx4_ASAP7_75t_R FILLER_172_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_622 ();
 DECAPx2_ASAP7_75t_R FILLER_172_643 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_649 ();
 DECAPx1_ASAP7_75t_R FILLER_172_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_667 ();
 DECAPx4_ASAP7_75t_R FILLER_172_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_694 ();
 DECAPx4_ASAP7_75t_R FILLER_172_703 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_772 ();
 DECAPx10_ASAP7_75t_R FILLER_172_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_172_821 ();
 DECAPx1_ASAP7_75t_R FILLER_172_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_838 ();
 DECAPx6_ASAP7_75t_R FILLER_172_856 ();
 DECAPx1_ASAP7_75t_R FILLER_172_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_172_874 ();
 DECAPx10_ASAP7_75t_R FILLER_173_2 ();
 DECAPx10_ASAP7_75t_R FILLER_173_24 ();
 DECAPx10_ASAP7_75t_R FILLER_173_46 ();
 DECAPx2_ASAP7_75t_R FILLER_173_68 ();
 DECAPx6_ASAP7_75t_R FILLER_173_106 ();
 DECAPx1_ASAP7_75t_R FILLER_173_128 ();
 DECAPx6_ASAP7_75t_R FILLER_173_138 ();
 DECAPx1_ASAP7_75t_R FILLER_173_158 ();
 FILLER_ASAP7_75t_R FILLER_173_165 ();
 DECAPx1_ASAP7_75t_R FILLER_173_182 ();
 DECAPx1_ASAP7_75t_R FILLER_173_192 ();
 DECAPx10_ASAP7_75t_R FILLER_173_199 ();
 DECAPx4_ASAP7_75t_R FILLER_173_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_231 ();
 FILLER_ASAP7_75t_R FILLER_173_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_243 ();
 DECAPx4_ASAP7_75t_R FILLER_173_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_353 ();
 FILLER_ASAP7_75t_R FILLER_173_408 ();
 FILLER_ASAP7_75t_R FILLER_173_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_443 ();
 DECAPx2_ASAP7_75t_R FILLER_173_472 ();
 DECAPx2_ASAP7_75t_R FILLER_173_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_503 ();
 DECAPx1_ASAP7_75t_R FILLER_173_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_518 ();
 DECAPx10_ASAP7_75t_R FILLER_173_526 ();
 DECAPx10_ASAP7_75t_R FILLER_173_548 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_173_570 ();
 DECAPx1_ASAP7_75t_R FILLER_173_600 ();
 DECAPx10_ASAP7_75t_R FILLER_173_619 ();
 DECAPx10_ASAP7_75t_R FILLER_173_641 ();
 DECAPx2_ASAP7_75t_R FILLER_173_663 ();
 FILLER_ASAP7_75t_R FILLER_173_669 ();
 DECAPx2_ASAP7_75t_R FILLER_173_679 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_693 ();
 DECAPx1_ASAP7_75t_R FILLER_173_715 ();
 DECAPx6_ASAP7_75t_R FILLER_173_745 ();
 FILLER_ASAP7_75t_R FILLER_173_759 ();
 DECAPx1_ASAP7_75t_R FILLER_173_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_796 ();
 DECAPx6_ASAP7_75t_R FILLER_173_803 ();
 DECAPx1_ASAP7_75t_R FILLER_173_817 ();
 FILLER_ASAP7_75t_R FILLER_173_847 ();
 DECAPx6_ASAP7_75t_R FILLER_173_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_173_933 ();
 DECAPx10_ASAP7_75t_R FILLER_174_2 ();
 DECAPx10_ASAP7_75t_R FILLER_174_24 ();
 DECAPx10_ASAP7_75t_R FILLER_174_46 ();
 DECAPx4_ASAP7_75t_R FILLER_174_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_78 ();
 FILLER_ASAP7_75t_R FILLER_174_87 ();
 DECAPx2_ASAP7_75t_R FILLER_174_92 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_98 ();
 DECAPx6_ASAP7_75t_R FILLER_174_109 ();
 DECAPx2_ASAP7_75t_R FILLER_174_129 ();
 DECAPx4_ASAP7_75t_R FILLER_174_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_151 ();
 FILLER_ASAP7_75t_R FILLER_174_158 ();
 DECAPx4_ASAP7_75t_R FILLER_174_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_176 ();
 DECAPx4_ASAP7_75t_R FILLER_174_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_229 ();
 DECAPx10_ASAP7_75t_R FILLER_174_236 ();
 DECAPx2_ASAP7_75t_R FILLER_174_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_264 ();
 DECAPx6_ASAP7_75t_R FILLER_174_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_291 ();
 DECAPx6_ASAP7_75t_R FILLER_174_295 ();
 DECAPx2_ASAP7_75t_R FILLER_174_309 ();
 DECAPx6_ASAP7_75t_R FILLER_174_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_338 ();
 DECAPx4_ASAP7_75t_R FILLER_174_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_374 ();
 FILLER_ASAP7_75t_R FILLER_174_381 ();
 DECAPx6_ASAP7_75t_R FILLER_174_386 ();
 DECAPx2_ASAP7_75t_R FILLER_174_409 ();
 DECAPx4_ASAP7_75t_R FILLER_174_422 ();
 FILLER_ASAP7_75t_R FILLER_174_432 ();
 DECAPx2_ASAP7_75t_R FILLER_174_443 ();
 DECAPx1_ASAP7_75t_R FILLER_174_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_461 ();
 DECAPx10_ASAP7_75t_R FILLER_174_464 ();
 DECAPx6_ASAP7_75t_R FILLER_174_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_517 ();
 DECAPx10_ASAP7_75t_R FILLER_174_526 ();
 DECAPx10_ASAP7_75t_R FILLER_174_548 ();
 DECAPx6_ASAP7_75t_R FILLER_174_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_584 ();
 DECAPx10_ASAP7_75t_R FILLER_174_593 ();
 DECAPx2_ASAP7_75t_R FILLER_174_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_621 ();
 DECAPx4_ASAP7_75t_R FILLER_174_641 ();
 DECAPx6_ASAP7_75t_R FILLER_174_657 ();
 DECAPx1_ASAP7_75t_R FILLER_174_671 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_688 ();
 DECAPx10_ASAP7_75t_R FILLER_174_705 ();
 DECAPx2_ASAP7_75t_R FILLER_174_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_733 ();
 DECAPx10_ASAP7_75t_R FILLER_174_740 ();
 FILLER_ASAP7_75t_R FILLER_174_762 ();
 DECAPx1_ASAP7_75t_R FILLER_174_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_775 ();
 DECAPx1_ASAP7_75t_R FILLER_174_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_783 ();
 FILLER_ASAP7_75t_R FILLER_174_823 ();
 FILLER_ASAP7_75t_R FILLER_174_831 ();
 DECAPx2_ASAP7_75t_R FILLER_174_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_174_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_861 ();
 FILLER_ASAP7_75t_R FILLER_174_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_174_887 ();
 FILLER_ASAP7_75t_R FILLER_174_911 ();
 FILLER_ASAP7_75t_R FILLER_174_927 ();
 DECAPx10_ASAP7_75t_R FILLER_175_2 ();
 DECAPx10_ASAP7_75t_R FILLER_175_24 ();
 DECAPx10_ASAP7_75t_R FILLER_175_46 ();
 DECAPx10_ASAP7_75t_R FILLER_175_68 ();
 DECAPx2_ASAP7_75t_R FILLER_175_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_96 ();
 DECAPx2_ASAP7_75t_R FILLER_175_107 ();
 DECAPx1_ASAP7_75t_R FILLER_175_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_123 ();
 FILLER_ASAP7_75t_R FILLER_175_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_138 ();
 FILLER_ASAP7_75t_R FILLER_175_145 ();
 DECAPx10_ASAP7_75t_R FILLER_175_173 ();
 DECAPx4_ASAP7_75t_R FILLER_175_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_205 ();
 DECAPx10_ASAP7_75t_R FILLER_175_244 ();
 DECAPx10_ASAP7_75t_R FILLER_175_266 ();
 DECAPx10_ASAP7_75t_R FILLER_175_288 ();
 DECAPx2_ASAP7_75t_R FILLER_175_310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_316 ();
 DECAPx6_ASAP7_75t_R FILLER_175_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_348 ();
 DECAPx6_ASAP7_75t_R FILLER_175_355 ();
 FILLER_ASAP7_75t_R FILLER_175_369 ();
 DECAPx10_ASAP7_75t_R FILLER_175_377 ();
 DECAPx10_ASAP7_75t_R FILLER_175_399 ();
 FILLER_ASAP7_75t_R FILLER_175_421 ();
 DECAPx2_ASAP7_75t_R FILLER_175_433 ();
 FILLER_ASAP7_75t_R FILLER_175_439 ();
 FILLER_ASAP7_75t_R FILLER_175_448 ();
 DECAPx4_ASAP7_75t_R FILLER_175_457 ();
 FILLER_ASAP7_75t_R FILLER_175_475 ();
 DECAPx10_ASAP7_75t_R FILLER_175_487 ();
 DECAPx6_ASAP7_75t_R FILLER_175_509 ();
 DECAPx1_ASAP7_75t_R FILLER_175_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_527 ();
 DECAPx1_ASAP7_75t_R FILLER_175_542 ();
 FILLER_ASAP7_75t_R FILLER_175_559 ();
 DECAPx10_ASAP7_75t_R FILLER_175_579 ();
 DECAPx4_ASAP7_75t_R FILLER_175_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_175_611 ();
 DECAPx1_ASAP7_75t_R FILLER_175_629 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_633 ();
 DECAPx1_ASAP7_75t_R FILLER_175_642 ();
 DECAPx2_ASAP7_75t_R FILLER_175_670 ();
 DECAPx4_ASAP7_75t_R FILLER_175_698 ();
 DECAPx4_ASAP7_75t_R FILLER_175_714 ();
 FILLER_ASAP7_75t_R FILLER_175_724 ();
 DECAPx10_ASAP7_75t_R FILLER_175_731 ();
 DECAPx10_ASAP7_75t_R FILLER_175_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_775 ();
 DECAPx1_ASAP7_75t_R FILLER_175_827 ();
 DECAPx2_ASAP7_75t_R FILLER_175_851 ();
 FILLER_ASAP7_75t_R FILLER_175_857 ();
 FILLER_ASAP7_75t_R FILLER_175_869 ();
 FILLER_ASAP7_75t_R FILLER_175_881 ();
 FILLER_ASAP7_75t_R FILLER_175_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_175_933 ();
 DECAPx10_ASAP7_75t_R FILLER_176_2 ();
 DECAPx10_ASAP7_75t_R FILLER_176_24 ();
 DECAPx10_ASAP7_75t_R FILLER_176_46 ();
 DECAPx4_ASAP7_75t_R FILLER_176_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_78 ();
 DECAPx2_ASAP7_75t_R FILLER_176_91 ();
 FILLER_ASAP7_75t_R FILLER_176_97 ();
 FILLER_ASAP7_75t_R FILLER_176_131 ();
 DECAPx10_ASAP7_75t_R FILLER_176_164 ();
 FILLER_ASAP7_75t_R FILLER_176_186 ();
 DECAPx10_ASAP7_75t_R FILLER_176_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_216 ();
 FILLER_ASAP7_75t_R FILLER_176_220 ();
 DECAPx1_ASAP7_75t_R FILLER_176_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_232 ();
 DECAPx2_ASAP7_75t_R FILLER_176_236 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_242 ();
 DECAPx1_ASAP7_75t_R FILLER_176_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_267 ();
 DECAPx2_ASAP7_75t_R FILLER_176_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_288 ();
 DECAPx2_ASAP7_75t_R FILLER_176_305 ();
 FILLER_ASAP7_75t_R FILLER_176_363 ();
 DECAPx4_ASAP7_75t_R FILLER_176_400 ();
 DECAPx6_ASAP7_75t_R FILLER_176_444 ();
 DECAPx1_ASAP7_75t_R FILLER_176_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_464 ();
 FILLER_ASAP7_75t_R FILLER_176_497 ();
 DECAPx6_ASAP7_75t_R FILLER_176_509 ();
 DECAPx2_ASAP7_75t_R FILLER_176_523 ();
 FILLER_ASAP7_75t_R FILLER_176_583 ();
 DECAPx2_ASAP7_75t_R FILLER_176_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_176_613 ();
 DECAPx1_ASAP7_75t_R FILLER_176_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_658 ();
 FILLER_ASAP7_75t_R FILLER_176_680 ();
 DECAPx2_ASAP7_75t_R FILLER_176_698 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_704 ();
 DECAPx1_ASAP7_75t_R FILLER_176_721 ();
 DECAPx1_ASAP7_75t_R FILLER_176_745 ();
 DECAPx6_ASAP7_75t_R FILLER_176_767 ();
 FILLER_ASAP7_75t_R FILLER_176_781 ();
 DECAPx1_ASAP7_75t_R FILLER_176_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_812 ();
 DECAPx4_ASAP7_75t_R FILLER_176_822 ();
 FILLER_ASAP7_75t_R FILLER_176_832 ();
 DECAPx10_ASAP7_75t_R FILLER_176_845 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_176_907 ();
 DECAPx10_ASAP7_75t_R FILLER_177_2 ();
 DECAPx10_ASAP7_75t_R FILLER_177_24 ();
 DECAPx10_ASAP7_75t_R FILLER_177_46 ();
 DECAPx1_ASAP7_75t_R FILLER_177_68 ();
 DECAPx2_ASAP7_75t_R FILLER_177_101 ();
 FILLER_ASAP7_75t_R FILLER_177_107 ();
 DECAPx1_ASAP7_75t_R FILLER_177_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_123 ();
 DECAPx2_ASAP7_75t_R FILLER_177_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_133 ();
 DECAPx2_ASAP7_75t_R FILLER_177_160 ();
 FILLER_ASAP7_75t_R FILLER_177_166 ();
 DECAPx2_ASAP7_75t_R FILLER_177_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_202 ();
 DECAPx6_ASAP7_75t_R FILLER_177_209 ();
 DECAPx2_ASAP7_75t_R FILLER_177_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_229 ();
 FILLER_ASAP7_75t_R FILLER_177_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_264 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_177_313 ();
 DECAPx1_ASAP7_75t_R FILLER_177_322 ();
 DECAPx10_ASAP7_75t_R FILLER_177_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_351 ();
 DECAPx1_ASAP7_75t_R FILLER_177_355 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_359 ();
 DECAPx1_ASAP7_75t_R FILLER_177_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_376 ();
 DECAPx4_ASAP7_75t_R FILLER_177_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_423 ();
 DECAPx10_ASAP7_75t_R FILLER_177_427 ();
 DECAPx10_ASAP7_75t_R FILLER_177_449 ();
 FILLER_ASAP7_75t_R FILLER_177_471 ();
 DECAPx1_ASAP7_75t_R FILLER_177_481 ();
 DECAPx4_ASAP7_75t_R FILLER_177_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_498 ();
 DECAPx4_ASAP7_75t_R FILLER_177_505 ();
 FILLER_ASAP7_75t_R FILLER_177_515 ();
 DECAPx1_ASAP7_75t_R FILLER_177_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_567 ();
 DECAPx2_ASAP7_75t_R FILLER_177_578 ();
 FILLER_ASAP7_75t_R FILLER_177_584 ();
 DECAPx1_ASAP7_75t_R FILLER_177_595 ();
 DECAPx10_ASAP7_75t_R FILLER_177_619 ();
 DECAPx1_ASAP7_75t_R FILLER_177_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_645 ();
 DECAPx2_ASAP7_75t_R FILLER_177_656 ();
 FILLER_ASAP7_75t_R FILLER_177_662 ();
 DECAPx2_ASAP7_75t_R FILLER_177_671 ();
 FILLER_ASAP7_75t_R FILLER_177_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_775 ();
 DECAPx6_ASAP7_75t_R FILLER_177_786 ();
 DECAPx2_ASAP7_75t_R FILLER_177_800 ();
 DECAPx10_ASAP7_75t_R FILLER_177_811 ();
 DECAPx6_ASAP7_75t_R FILLER_177_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_177_924 ();
 FILLER_ASAP7_75t_R FILLER_177_927 ();
 DECAPx10_ASAP7_75t_R FILLER_178_2 ();
 DECAPx10_ASAP7_75t_R FILLER_178_24 ();
 DECAPx10_ASAP7_75t_R FILLER_178_46 ();
 DECAPx6_ASAP7_75t_R FILLER_178_68 ();
 DECAPx1_ASAP7_75t_R FILLER_178_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_86 ();
 DECAPx2_ASAP7_75t_R FILLER_178_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_96 ();
 DECAPx10_ASAP7_75t_R FILLER_178_105 ();
 DECAPx6_ASAP7_75t_R FILLER_178_127 ();
 DECAPx2_ASAP7_75t_R FILLER_178_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_147 ();
 DECAPx2_ASAP7_75t_R FILLER_178_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_211 ();
 DECAPx2_ASAP7_75t_R FILLER_178_218 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_293 ();
 FILLER_ASAP7_75t_R FILLER_178_308 ();
 DECAPx6_ASAP7_75t_R FILLER_178_316 ();
 DECAPx2_ASAP7_75t_R FILLER_178_330 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_351 ();
 FILLER_ASAP7_75t_R FILLER_178_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_378 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_382 ();
 DECAPx1_ASAP7_75t_R FILLER_178_389 ();
 DECAPx2_ASAP7_75t_R FILLER_178_424 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_430 ();
 FILLER_ASAP7_75t_R FILLER_178_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_461 ();
 DECAPx4_ASAP7_75t_R FILLER_178_464 ();
 FILLER_ASAP7_75t_R FILLER_178_474 ();
 DECAPx2_ASAP7_75t_R FILLER_178_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_508 ();
 DECAPx2_ASAP7_75t_R FILLER_178_527 ();
 DECAPx1_ASAP7_75t_R FILLER_178_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_543 ();
 DECAPx10_ASAP7_75t_R FILLER_178_550 ();
 DECAPx2_ASAP7_75t_R FILLER_178_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_585 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_597 ();
 DECAPx10_ASAP7_75t_R FILLER_178_623 ();
 DECAPx6_ASAP7_75t_R FILLER_178_645 ();
 DECAPx1_ASAP7_75t_R FILLER_178_659 ();
 DECAPx4_ASAP7_75t_R FILLER_178_679 ();
 FILLER_ASAP7_75t_R FILLER_178_689 ();
 DECAPx6_ASAP7_75t_R FILLER_178_697 ();
 DECAPx2_ASAP7_75t_R FILLER_178_711 ();
 DECAPx2_ASAP7_75t_R FILLER_178_756 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_762 ();
 DECAPx10_ASAP7_75t_R FILLER_178_785 ();
 DECAPx6_ASAP7_75t_R FILLER_178_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_178_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_178_933 ();
 DECAPx10_ASAP7_75t_R FILLER_179_7 ();
 DECAPx10_ASAP7_75t_R FILLER_179_29 ();
 DECAPx10_ASAP7_75t_R FILLER_179_51 ();
 DECAPx1_ASAP7_75t_R FILLER_179_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_77 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_90 ();
 DECAPx10_ASAP7_75t_R FILLER_179_105 ();
 DECAPx10_ASAP7_75t_R FILLER_179_127 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_149 ();
 DECAPx2_ASAP7_75t_R FILLER_179_184 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_207 ();
 DECAPx1_ASAP7_75t_R FILLER_179_230 ();
 FILLER_ASAP7_75t_R FILLER_179_240 ();
 DECAPx2_ASAP7_75t_R FILLER_179_245 ();
 DECAPx10_ASAP7_75t_R FILLER_179_257 ();
 DECAPx10_ASAP7_75t_R FILLER_179_279 ();
 DECAPx1_ASAP7_75t_R FILLER_179_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_305 ();
 DECAPx1_ASAP7_75t_R FILLER_179_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_370 ();
 DECAPx2_ASAP7_75t_R FILLER_179_378 ();
 DECAPx4_ASAP7_75t_R FILLER_179_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_426 ();
 DECAPx2_ASAP7_75t_R FILLER_179_453 ();
 FILLER_ASAP7_75t_R FILLER_179_459 ();
 DECAPx6_ASAP7_75t_R FILLER_179_467 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_481 ();
 DECAPx10_ASAP7_75t_R FILLER_179_512 ();
 DECAPx10_ASAP7_75t_R FILLER_179_534 ();
 DECAPx10_ASAP7_75t_R FILLER_179_556 ();
 DECAPx10_ASAP7_75t_R FILLER_179_578 ();
 DECAPx2_ASAP7_75t_R FILLER_179_600 ();
 FILLER_ASAP7_75t_R FILLER_179_606 ();
 DECAPx10_ASAP7_75t_R FILLER_179_613 ();
 DECAPx10_ASAP7_75t_R FILLER_179_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_657 ();
 DECAPx10_ASAP7_75t_R FILLER_179_667 ();
 DECAPx2_ASAP7_75t_R FILLER_179_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_695 ();
 DECAPx10_ASAP7_75t_R FILLER_179_706 ();
 DECAPx4_ASAP7_75t_R FILLER_179_728 ();
 FILLER_ASAP7_75t_R FILLER_179_738 ();
 DECAPx10_ASAP7_75t_R FILLER_179_748 ();
 DECAPx4_ASAP7_75t_R FILLER_179_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_795 ();
 FILLER_ASAP7_75t_R FILLER_179_808 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_852 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_179_879 ();
 FILLER_ASAP7_75t_R FILLER_179_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_179_921 ();
 DECAPx10_ASAP7_75t_R FILLER_180_7 ();
 DECAPx10_ASAP7_75t_R FILLER_180_29 ();
 DECAPx10_ASAP7_75t_R FILLER_180_51 ();
 DECAPx1_ASAP7_75t_R FILLER_180_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_111 ();
 FILLER_ASAP7_75t_R FILLER_180_118 ();
 DECAPx10_ASAP7_75t_R FILLER_180_129 ();
 DECAPx1_ASAP7_75t_R FILLER_180_151 ();
 DECAPx1_ASAP7_75t_R FILLER_180_161 ();
 DECAPx1_ASAP7_75t_R FILLER_180_168 ();
 DECAPx10_ASAP7_75t_R FILLER_180_175 ();
 DECAPx10_ASAP7_75t_R FILLER_180_197 ();
 DECAPx10_ASAP7_75t_R FILLER_180_219 ();
 DECAPx10_ASAP7_75t_R FILLER_180_241 ();
 DECAPx10_ASAP7_75t_R FILLER_180_263 ();
 DECAPx10_ASAP7_75t_R FILLER_180_285 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_336 ();
 DECAPx4_ASAP7_75t_R FILLER_180_386 ();
 FILLER_ASAP7_75t_R FILLER_180_396 ();
 DECAPx6_ASAP7_75t_R FILLER_180_404 ();
 DECAPx1_ASAP7_75t_R FILLER_180_418 ();
 FILLER_ASAP7_75t_R FILLER_180_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_464 ();
 DECAPx6_ASAP7_75t_R FILLER_180_471 ();
 DECAPx2_ASAP7_75t_R FILLER_180_485 ();
 DECAPx6_ASAP7_75t_R FILLER_180_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_508 ();
 DECAPx4_ASAP7_75t_R FILLER_180_517 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_527 ();
 DECAPx2_ASAP7_75t_R FILLER_180_536 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_542 ();
 DECAPx2_ASAP7_75t_R FILLER_180_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_559 ();
 DECAPx2_ASAP7_75t_R FILLER_180_567 ();
 DECAPx10_ASAP7_75t_R FILLER_180_580 ();
 DECAPx6_ASAP7_75t_R FILLER_180_602 ();
 DECAPx2_ASAP7_75t_R FILLER_180_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_622 ();
 FILLER_ASAP7_75t_R FILLER_180_634 ();
 DECAPx1_ASAP7_75t_R FILLER_180_653 ();
 DECAPx4_ASAP7_75t_R FILLER_180_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_180_673 ();
 FILLER_ASAP7_75t_R FILLER_180_694 ();
 DECAPx10_ASAP7_75t_R FILLER_180_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_738 ();
 DECAPx4_ASAP7_75t_R FILLER_180_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_775 ();
 FILLER_ASAP7_75t_R FILLER_180_802 ();
 FILLER_ASAP7_75t_R FILLER_180_833 ();
 DECAPx6_ASAP7_75t_R FILLER_180_841 ();
 DECAPx1_ASAP7_75t_R FILLER_180_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_180_902 ();
 DECAPx10_ASAP7_75t_R FILLER_181_2 ();
 DECAPx10_ASAP7_75t_R FILLER_181_24 ();
 DECAPx10_ASAP7_75t_R FILLER_181_46 ();
 DECAPx6_ASAP7_75t_R FILLER_181_68 ();
 DECAPx2_ASAP7_75t_R FILLER_181_82 ();
 DECAPx6_ASAP7_75t_R FILLER_181_91 ();
 DECAPx2_ASAP7_75t_R FILLER_181_137 ();
 DECAPx10_ASAP7_75t_R FILLER_181_155 ();
 DECAPx10_ASAP7_75t_R FILLER_181_177 ();
 DECAPx10_ASAP7_75t_R FILLER_181_199 ();
 DECAPx2_ASAP7_75t_R FILLER_181_221 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_227 ();
 DECAPx10_ASAP7_75t_R FILLER_181_236 ();
 DECAPx6_ASAP7_75t_R FILLER_181_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_302 ();
 DECAPx4_ASAP7_75t_R FILLER_181_309 ();
 FILLER_ASAP7_75t_R FILLER_181_319 ();
 DECAPx1_ASAP7_75t_R FILLER_181_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_346 ();
 DECAPx6_ASAP7_75t_R FILLER_181_391 ();
 FILLER_ASAP7_75t_R FILLER_181_405 ();
 DECAPx1_ASAP7_75t_R FILLER_181_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_431 ();
 FILLER_ASAP7_75t_R FILLER_181_445 ();
 DECAPx1_ASAP7_75t_R FILLER_181_454 ();
 DECAPx2_ASAP7_75t_R FILLER_181_466 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_472 ();
 DECAPx6_ASAP7_75t_R FILLER_181_487 ();
 DECAPx1_ASAP7_75t_R FILLER_181_501 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_505 ();
 DECAPx4_ASAP7_75t_R FILLER_181_513 ();
 DECAPx1_ASAP7_75t_R FILLER_181_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_555 ();
 DECAPx1_ASAP7_75t_R FILLER_181_574 ();
 DECAPx6_ASAP7_75t_R FILLER_181_586 ();
 DECAPx2_ASAP7_75t_R FILLER_181_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_606 ();
 DECAPx2_ASAP7_75t_R FILLER_181_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_619 ();
 FILLER_ASAP7_75t_R FILLER_181_636 ();
 FILLER_ASAP7_75t_R FILLER_181_669 ();
 DECAPx1_ASAP7_75t_R FILLER_181_679 ();
 DECAPx4_ASAP7_75t_R FILLER_181_699 ();
 DECAPx1_ASAP7_75t_R FILLER_181_716 ();
 FILLER_ASAP7_75t_R FILLER_181_734 ();
 DECAPx2_ASAP7_75t_R FILLER_181_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_749 ();
 DECAPx1_ASAP7_75t_R FILLER_181_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_780 ();
 DECAPx2_ASAP7_75t_R FILLER_181_804 ();
 FILLER_ASAP7_75t_R FILLER_181_824 ();
 DECAPx6_ASAP7_75t_R FILLER_181_833 ();
 FILLER_ASAP7_75t_R FILLER_181_847 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_181_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_181_933 ();
 DECAPx10_ASAP7_75t_R FILLER_182_7 ();
 DECAPx10_ASAP7_75t_R FILLER_182_29 ();
 DECAPx10_ASAP7_75t_R FILLER_182_51 ();
 DECAPx10_ASAP7_75t_R FILLER_182_73 ();
 DECAPx4_ASAP7_75t_R FILLER_182_95 ();
 DECAPx1_ASAP7_75t_R FILLER_182_111 ();
 FILLER_ASAP7_75t_R FILLER_182_121 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_129 ();
 DECAPx6_ASAP7_75t_R FILLER_182_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_198 ();
 FILLER_ASAP7_75t_R FILLER_182_205 ();
 DECAPx2_ASAP7_75t_R FILLER_182_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_225 ();
 DECAPx4_ASAP7_75t_R FILLER_182_252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_268 ();
 DECAPx1_ASAP7_75t_R FILLER_182_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_297 ();
 DECAPx4_ASAP7_75t_R FILLER_182_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_356 ();
 DECAPx1_ASAP7_75t_R FILLER_182_388 ();
 DECAPx6_ASAP7_75t_R FILLER_182_431 ();
 FILLER_ASAP7_75t_R FILLER_182_445 ();
 DECAPx2_ASAP7_75t_R FILLER_182_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_459 ();
 DECAPx2_ASAP7_75t_R FILLER_182_464 ();
 FILLER_ASAP7_75t_R FILLER_182_470 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_501 ();
 DECAPx10_ASAP7_75t_R FILLER_182_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_538 ();
 DECAPx1_ASAP7_75t_R FILLER_182_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_624 ();
 DECAPx4_ASAP7_75t_R FILLER_182_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_671 ();
 DECAPx2_ASAP7_75t_R FILLER_182_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_694 ();
 DECAPx2_ASAP7_75t_R FILLER_182_702 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_732 ();
 DECAPx1_ASAP7_75t_R FILLER_182_788 ();
 DECAPx10_ASAP7_75t_R FILLER_182_797 ();
 DECAPx10_ASAP7_75t_R FILLER_182_819 ();
 DECAPx4_ASAP7_75t_R FILLER_182_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_182_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_182_897 ();
 FILLER_ASAP7_75t_R FILLER_182_917 ();
 DECAPx10_ASAP7_75t_R FILLER_183_7 ();
 DECAPx10_ASAP7_75t_R FILLER_183_29 ();
 DECAPx10_ASAP7_75t_R FILLER_183_51 ();
 DECAPx1_ASAP7_75t_R FILLER_183_73 ();
 DECAPx10_ASAP7_75t_R FILLER_183_89 ();
 DECAPx4_ASAP7_75t_R FILLER_183_111 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_156 ();
 DECAPx2_ASAP7_75t_R FILLER_183_165 ();
 FILLER_ASAP7_75t_R FILLER_183_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_216 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_229 ();
 DECAPx2_ASAP7_75t_R FILLER_183_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_280 ();
 DECAPx1_ASAP7_75t_R FILLER_183_287 ();
 DECAPx6_ASAP7_75t_R FILLER_183_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_308 ();
 DECAPx6_ASAP7_75t_R FILLER_183_315 ();
 DECAPx2_ASAP7_75t_R FILLER_183_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_335 ();
 FILLER_ASAP7_75t_R FILLER_183_345 ();
 DECAPx2_ASAP7_75t_R FILLER_183_350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_356 ();
 DECAPx4_ASAP7_75t_R FILLER_183_365 ();
 FILLER_ASAP7_75t_R FILLER_183_375 ();
 DECAPx4_ASAP7_75t_R FILLER_183_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_404 ();
 DECAPx4_ASAP7_75t_R FILLER_183_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_434 ();
 DECAPx2_ASAP7_75t_R FILLER_183_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_493 ();
 DECAPx2_ASAP7_75t_R FILLER_183_504 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_510 ();
 DECAPx10_ASAP7_75t_R FILLER_183_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_541 ();
 DECAPx1_ASAP7_75t_R FILLER_183_550 ();
 DECAPx4_ASAP7_75t_R FILLER_183_557 ();
 FILLER_ASAP7_75t_R FILLER_183_567 ();
 DECAPx2_ASAP7_75t_R FILLER_183_575 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_615 ();
 DECAPx10_ASAP7_75t_R FILLER_183_638 ();
 DECAPx2_ASAP7_75t_R FILLER_183_660 ();
 FILLER_ASAP7_75t_R FILLER_183_666 ();
 DECAPx2_ASAP7_75t_R FILLER_183_681 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_183_687 ();
 DECAPx4_ASAP7_75t_R FILLER_183_696 ();
 FILLER_ASAP7_75t_R FILLER_183_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_714 ();
 DECAPx2_ASAP7_75t_R FILLER_183_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_727 ();
 DECAPx2_ASAP7_75t_R FILLER_183_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_750 ();
 DECAPx10_ASAP7_75t_R FILLER_183_779 ();
 DECAPx10_ASAP7_75t_R FILLER_183_801 ();
 DECAPx4_ASAP7_75t_R FILLER_183_823 ();
 DECAPx10_ASAP7_75t_R FILLER_183_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_183_919 ();
 FILLER_ASAP7_75t_R FILLER_183_927 ();
 DECAPx10_ASAP7_75t_R FILLER_184_7 ();
 DECAPx10_ASAP7_75t_R FILLER_184_29 ();
 DECAPx6_ASAP7_75t_R FILLER_184_51 ();
 DECAPx2_ASAP7_75t_R FILLER_184_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_71 ();
 DECAPx1_ASAP7_75t_R FILLER_184_98 ();
 DECAPx6_ASAP7_75t_R FILLER_184_110 ();
 DECAPx1_ASAP7_75t_R FILLER_184_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_128 ();
 DECAPx4_ASAP7_75t_R FILLER_184_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_145 ();
 DECAPx1_ASAP7_75t_R FILLER_184_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_193 ();
 DECAPx10_ASAP7_75t_R FILLER_184_199 ();
 DECAPx4_ASAP7_75t_R FILLER_184_221 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_237 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_246 ();
 DECAPx6_ASAP7_75t_R FILLER_184_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_291 ();
 DECAPx2_ASAP7_75t_R FILLER_184_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_329 ();
 DECAPx2_ASAP7_75t_R FILLER_184_342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_348 ();
 FILLER_ASAP7_75t_R FILLER_184_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_383 ();
 DECAPx2_ASAP7_75t_R FILLER_184_403 ();
 DECAPx1_ASAP7_75t_R FILLER_184_423 ();
 DECAPx1_ASAP7_75t_R FILLER_184_441 ();
 DECAPx2_ASAP7_75t_R FILLER_184_454 ();
 FILLER_ASAP7_75t_R FILLER_184_460 ();
 DECAPx4_ASAP7_75t_R FILLER_184_464 ();
 DECAPx2_ASAP7_75t_R FILLER_184_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_483 ();
 DECAPx1_ASAP7_75t_R FILLER_184_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_498 ();
 DECAPx2_ASAP7_75t_R FILLER_184_506 ();
 DECAPx10_ASAP7_75t_R FILLER_184_521 ();
 DECAPx10_ASAP7_75t_R FILLER_184_543 ();
 DECAPx10_ASAP7_75t_R FILLER_184_565 ();
 FILLER_ASAP7_75t_R FILLER_184_590 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_621 ();
 DECAPx10_ASAP7_75t_R FILLER_184_629 ();
 DECAPx6_ASAP7_75t_R FILLER_184_651 ();
 DECAPx10_ASAP7_75t_R FILLER_184_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_696 ();
 DECAPx1_ASAP7_75t_R FILLER_184_717 ();
 FILLER_ASAP7_75t_R FILLER_184_735 ();
 DECAPx4_ASAP7_75t_R FILLER_184_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_759 ();
 DECAPx6_ASAP7_75t_R FILLER_184_768 ();
 DECAPx2_ASAP7_75t_R FILLER_184_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_788 ();
 DECAPx1_ASAP7_75t_R FILLER_184_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_799 ();
 FILLER_ASAP7_75t_R FILLER_184_806 ();
 DECAPx1_ASAP7_75t_R FILLER_184_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_184_860 ();
 DECAPx1_ASAP7_75t_R FILLER_184_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_184_909 ();
 DECAPx10_ASAP7_75t_R FILLER_185_2 ();
 DECAPx10_ASAP7_75t_R FILLER_185_24 ();
 DECAPx10_ASAP7_75t_R FILLER_185_46 ();
 DECAPx4_ASAP7_75t_R FILLER_185_68 ();
 FILLER_ASAP7_75t_R FILLER_185_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_89 ();
 DECAPx10_ASAP7_75t_R FILLER_185_113 ();
 DECAPx6_ASAP7_75t_R FILLER_185_135 ();
 DECAPx1_ASAP7_75t_R FILLER_185_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_160 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_166 ();
 DECAPx10_ASAP7_75t_R FILLER_185_175 ();
 DECAPx4_ASAP7_75t_R FILLER_185_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_207 ();
 FILLER_ASAP7_75t_R FILLER_185_214 ();
 DECAPx1_ASAP7_75t_R FILLER_185_242 ();
 DECAPx1_ASAP7_75t_R FILLER_185_254 ();
 DECAPx1_ASAP7_75t_R FILLER_185_272 ();
 DECAPx10_ASAP7_75t_R FILLER_185_282 ();
 DECAPx6_ASAP7_75t_R FILLER_185_304 ();
 DECAPx2_ASAP7_75t_R FILLER_185_318 ();
 FILLER_ASAP7_75t_R FILLER_185_350 ();
 DECAPx1_ASAP7_75t_R FILLER_185_360 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_413 ();
 DECAPx1_ASAP7_75t_R FILLER_185_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_437 ();
 DECAPx6_ASAP7_75t_R FILLER_185_446 ();
 FILLER_ASAP7_75t_R FILLER_185_460 ();
 DECAPx10_ASAP7_75t_R FILLER_185_468 ();
 DECAPx6_ASAP7_75t_R FILLER_185_490 ();
 DECAPx1_ASAP7_75t_R FILLER_185_504 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_514 ();
 DECAPx10_ASAP7_75t_R FILLER_185_544 ();
 DECAPx10_ASAP7_75t_R FILLER_185_566 ();
 DECAPx6_ASAP7_75t_R FILLER_185_588 ();
 DECAPx1_ASAP7_75t_R FILLER_185_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_606 ();
 DECAPx10_ASAP7_75t_R FILLER_185_613 ();
 DECAPx2_ASAP7_75t_R FILLER_185_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_641 ();
 FILLER_ASAP7_75t_R FILLER_185_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_664 ();
 DECAPx6_ASAP7_75t_R FILLER_185_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_691 ();
 DECAPx4_ASAP7_75t_R FILLER_185_698 ();
 DECAPx10_ASAP7_75t_R FILLER_185_714 ();
 DECAPx6_ASAP7_75t_R FILLER_185_736 ();
 DECAPx6_ASAP7_75t_R FILLER_185_765 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_185_785 ();
 DECAPx1_ASAP7_75t_R FILLER_185_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_836 ();
 DECAPx1_ASAP7_75t_R FILLER_185_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_185_867 ();
 FILLER_ASAP7_75t_R FILLER_185_878 ();
 DECAPx10_ASAP7_75t_R FILLER_186_2 ();
 DECAPx10_ASAP7_75t_R FILLER_186_24 ();
 DECAPx10_ASAP7_75t_R FILLER_186_46 ();
 DECAPx4_ASAP7_75t_R FILLER_186_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_78 ();
 DECAPx6_ASAP7_75t_R FILLER_186_105 ();
 FILLER_ASAP7_75t_R FILLER_186_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_127 ();
 DECAPx2_ASAP7_75t_R FILLER_186_131 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_137 ();
 DECAPx1_ASAP7_75t_R FILLER_186_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_186_165 ();
 DECAPx6_ASAP7_75t_R FILLER_186_182 ();
 FILLER_ASAP7_75t_R FILLER_186_196 ();
 FILLER_ASAP7_75t_R FILLER_186_224 ();
 DECAPx10_ASAP7_75t_R FILLER_186_235 ();
 DECAPx1_ASAP7_75t_R FILLER_186_257 ();
 DECAPx4_ASAP7_75t_R FILLER_186_287 ();
 DECAPx4_ASAP7_75t_R FILLER_186_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_315 ();
 DECAPx2_ASAP7_75t_R FILLER_186_331 ();
 FILLER_ASAP7_75t_R FILLER_186_337 ();
 DECAPx1_ASAP7_75t_R FILLER_186_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_346 ();
 DECAPx4_ASAP7_75t_R FILLER_186_401 ();
 FILLER_ASAP7_75t_R FILLER_186_411 ();
 DECAPx1_ASAP7_75t_R FILLER_186_439 ();
 FILLER_ASAP7_75t_R FILLER_186_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_461 ();
 FILLER_ASAP7_75t_R FILLER_186_464 ();
 DECAPx10_ASAP7_75t_R FILLER_186_474 ();
 DECAPx10_ASAP7_75t_R FILLER_186_496 ();
 DECAPx2_ASAP7_75t_R FILLER_186_518 ();
 DECAPx2_ASAP7_75t_R FILLER_186_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_551 ();
 DECAPx6_ASAP7_75t_R FILLER_186_562 ();
 DECAPx10_ASAP7_75t_R FILLER_186_584 ();
 DECAPx6_ASAP7_75t_R FILLER_186_606 ();
 DECAPx2_ASAP7_75t_R FILLER_186_625 ();
 FILLER_ASAP7_75t_R FILLER_186_631 ();
 DECAPx1_ASAP7_75t_R FILLER_186_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_648 ();
 DECAPx2_ASAP7_75t_R FILLER_186_670 ();
 FILLER_ASAP7_75t_R FILLER_186_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_699 ();
 DECAPx6_ASAP7_75t_R FILLER_186_710 ();
 DECAPx1_ASAP7_75t_R FILLER_186_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_728 ();
 DECAPx1_ASAP7_75t_R FILLER_186_735 ();
 DECAPx10_ASAP7_75t_R FILLER_186_745 ();
 DECAPx2_ASAP7_75t_R FILLER_186_767 ();
 FILLER_ASAP7_75t_R FILLER_186_811 ();
 FILLER_ASAP7_75t_R FILLER_186_842 ();
 FILLERxp5_ASAP7_75t_R FILLER_186_902 ();
 DECAPx10_ASAP7_75t_R FILLER_187_7 ();
 DECAPx10_ASAP7_75t_R FILLER_187_29 ();
 DECAPx10_ASAP7_75t_R FILLER_187_51 ();
 DECAPx6_ASAP7_75t_R FILLER_187_73 ();
 FILLER_ASAP7_75t_R FILLER_187_87 ();
 DECAPx4_ASAP7_75t_R FILLER_187_98 ();
 DECAPx1_ASAP7_75t_R FILLER_187_143 ();
 DECAPx6_ASAP7_75t_R FILLER_187_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_212 ();
 FILLER_ASAP7_75t_R FILLER_187_216 ();
 DECAPx10_ASAP7_75t_R FILLER_187_221 ();
 DECAPx1_ASAP7_75t_R FILLER_187_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_247 ();
 DECAPx2_ASAP7_75t_R FILLER_187_272 ();
 DECAPx10_ASAP7_75t_R FILLER_187_316 ();
 DECAPx10_ASAP7_75t_R FILLER_187_338 ();
 DECAPx6_ASAP7_75t_R FILLER_187_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_374 ();
 DECAPx1_ASAP7_75t_R FILLER_187_383 ();
 FILLER_ASAP7_75t_R FILLER_187_393 ();
 DECAPx10_ASAP7_75t_R FILLER_187_401 ();
 DECAPx1_ASAP7_75t_R FILLER_187_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_457 ();
 DECAPx1_ASAP7_75t_R FILLER_187_484 ();
 DECAPx10_ASAP7_75t_R FILLER_187_500 ();
 FILLER_ASAP7_75t_R FILLER_187_522 ();
 DECAPx2_ASAP7_75t_R FILLER_187_530 ();
 DECAPx1_ASAP7_75t_R FILLER_187_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_566 ();
 DECAPx6_ASAP7_75t_R FILLER_187_592 ();
 DECAPx1_ASAP7_75t_R FILLER_187_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_633 ();
 FILLER_ASAP7_75t_R FILLER_187_642 ();
 DECAPx6_ASAP7_75t_R FILLER_187_661 ();
 FILLER_ASAP7_75t_R FILLER_187_675 ();
 DECAPx6_ASAP7_75t_R FILLER_187_699 ();
 DECAPx1_ASAP7_75t_R FILLER_187_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_717 ();
 DECAPx2_ASAP7_75t_R FILLER_187_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_763 ();
 DECAPx1_ASAP7_75t_R FILLER_187_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_187_796 ();
 DECAPx2_ASAP7_75t_R FILLER_187_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_842 ();
 FILLER_ASAP7_75t_R FILLER_187_856 ();
 DECAPx4_ASAP7_75t_R FILLER_187_861 ();
 DECAPx6_ASAP7_75t_R FILLER_187_876 ();
 FILLER_ASAP7_75t_R FILLER_187_893 ();
 FILLERxp5_ASAP7_75t_R FILLER_187_933 ();
 DECAPx10_ASAP7_75t_R FILLER_188_2 ();
 DECAPx10_ASAP7_75t_R FILLER_188_24 ();
 DECAPx10_ASAP7_75t_R FILLER_188_46 ();
 DECAPx10_ASAP7_75t_R FILLER_188_68 ();
 DECAPx10_ASAP7_75t_R FILLER_188_90 ();
 DECAPx2_ASAP7_75t_R FILLER_188_112 ();
 DECAPx2_ASAP7_75t_R FILLER_188_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_130 ();
 DECAPx10_ASAP7_75t_R FILLER_188_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_161 ();
 DECAPx6_ASAP7_75t_R FILLER_188_165 ();
 DECAPx1_ASAP7_75t_R FILLER_188_179 ();
 DECAPx10_ASAP7_75t_R FILLER_188_195 ();
 DECAPx2_ASAP7_75t_R FILLER_188_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_223 ();
 FILLER_ASAP7_75t_R FILLER_188_233 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_238 ();
 DECAPx10_ASAP7_75t_R FILLER_188_247 ();
 DECAPx2_ASAP7_75t_R FILLER_188_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_275 ();
 DECAPx1_ASAP7_75t_R FILLER_188_308 ();
 DECAPx2_ASAP7_75t_R FILLER_188_322 ();
 FILLER_ASAP7_75t_R FILLER_188_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_336 ();
 DECAPx1_ASAP7_75t_R FILLER_188_343 ();
 DECAPx10_ASAP7_75t_R FILLER_188_350 ();
 DECAPx4_ASAP7_75t_R FILLER_188_372 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_382 ();
 DECAPx10_ASAP7_75t_R FILLER_188_409 ();
 DECAPx6_ASAP7_75t_R FILLER_188_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_449 ();
 DECAPx1_ASAP7_75t_R FILLER_188_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_472 ();
 DECAPx2_ASAP7_75t_R FILLER_188_476 ();
 FILLER_ASAP7_75t_R FILLER_188_508 ();
 DECAPx10_ASAP7_75t_R FILLER_188_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_556 ();
 DECAPx6_ASAP7_75t_R FILLER_188_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_579 ();
 DECAPx6_ASAP7_75t_R FILLER_188_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_627 ();
 DECAPx2_ASAP7_75t_R FILLER_188_634 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_188_640 ();
 DECAPx6_ASAP7_75t_R FILLER_188_650 ();
 DECAPx2_ASAP7_75t_R FILLER_188_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_670 ();
 DECAPx6_ASAP7_75t_R FILLER_188_689 ();
 FILLER_ASAP7_75t_R FILLER_188_703 ();
 DECAPx10_ASAP7_75t_R FILLER_188_710 ();
 FILLER_ASAP7_75t_R FILLER_188_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_760 ();
 DECAPx10_ASAP7_75t_R FILLER_188_791 ();
 DECAPx6_ASAP7_75t_R FILLER_188_813 ();
 DECAPx1_ASAP7_75t_R FILLER_188_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_831 ();
 DECAPx10_ASAP7_75t_R FILLER_188_835 ();
 DECAPx10_ASAP7_75t_R FILLER_188_857 ();
 DECAPx10_ASAP7_75t_R FILLER_188_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_907 ();
 FILLERxp5_ASAP7_75t_R FILLER_188_933 ();
 DECAPx10_ASAP7_75t_R FILLER_189_2 ();
 DECAPx10_ASAP7_75t_R FILLER_189_24 ();
 DECAPx10_ASAP7_75t_R FILLER_189_46 ();
 DECAPx6_ASAP7_75t_R FILLER_189_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_82 ();
 FILLER_ASAP7_75t_R FILLER_189_97 ();
 FILLER_ASAP7_75t_R FILLER_189_105 ();
 DECAPx10_ASAP7_75t_R FILLER_189_115 ();
 DECAPx4_ASAP7_75t_R FILLER_189_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_153 ();
 DECAPx6_ASAP7_75t_R FILLER_189_162 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_176 ();
 DECAPx10_ASAP7_75t_R FILLER_189_187 ();
 DECAPx4_ASAP7_75t_R FILLER_189_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_252 ();
 FILLER_ASAP7_75t_R FILLER_189_265 ();
 DECAPx4_ASAP7_75t_R FILLER_189_274 ();
 FILLER_ASAP7_75t_R FILLER_189_284 ();
 DECAPx6_ASAP7_75t_R FILLER_189_310 ();
 FILLER_ASAP7_75t_R FILLER_189_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_360 ();
 DECAPx4_ASAP7_75t_R FILLER_189_367 ();
 DECAPx2_ASAP7_75t_R FILLER_189_389 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_395 ();
 DECAPx2_ASAP7_75t_R FILLER_189_401 ();
 FILLER_ASAP7_75t_R FILLER_189_407 ();
 DECAPx10_ASAP7_75t_R FILLER_189_432 ();
 DECAPx6_ASAP7_75t_R FILLER_189_454 ();
 FILLER_ASAP7_75t_R FILLER_189_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_493 ();
 DECAPx2_ASAP7_75t_R FILLER_189_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_506 ();
 FILLER_ASAP7_75t_R FILLER_189_513 ();
 DECAPx10_ASAP7_75t_R FILLER_189_522 ();
 DECAPx10_ASAP7_75t_R FILLER_189_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_566 ();
 DECAPx2_ASAP7_75t_R FILLER_189_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_613 ();
 DECAPx10_ASAP7_75t_R FILLER_189_625 ();
 DECAPx6_ASAP7_75t_R FILLER_189_647 ();
 FILLER_ASAP7_75t_R FILLER_189_661 ();
 DECAPx10_ASAP7_75t_R FILLER_189_672 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_703 ();
 DECAPx4_ASAP7_75t_R FILLER_189_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_746 ();
 DECAPx2_ASAP7_75t_R FILLER_189_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_189_763 ();
 DECAPx10_ASAP7_75t_R FILLER_189_779 ();
 DECAPx10_ASAP7_75t_R FILLER_189_801 ();
 DECAPx10_ASAP7_75t_R FILLER_189_835 ();
 DECAPx4_ASAP7_75t_R FILLER_189_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_867 ();
 DECAPx10_ASAP7_75t_R FILLER_189_878 ();
 DECAPx1_ASAP7_75t_R FILLER_189_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_189_927 ();
 DECAPx10_ASAP7_75t_R FILLER_190_2 ();
 DECAPx10_ASAP7_75t_R FILLER_190_24 ();
 DECAPx10_ASAP7_75t_R FILLER_190_46 ();
 DECAPx6_ASAP7_75t_R FILLER_190_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_116 ();
 DECAPx2_ASAP7_75t_R FILLER_190_123 ();
 DECAPx4_ASAP7_75t_R FILLER_190_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_169 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_173 ();
 DECAPx1_ASAP7_75t_R FILLER_190_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_194 ();
 DECAPx6_ASAP7_75t_R FILLER_190_215 ();
 FILLER_ASAP7_75t_R FILLER_190_229 ();
 DECAPx2_ASAP7_75t_R FILLER_190_237 ();
 FILLER_ASAP7_75t_R FILLER_190_243 ();
 FILLER_ASAP7_75t_R FILLER_190_261 ();
 DECAPx4_ASAP7_75t_R FILLER_190_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_295 ();
 DECAPx4_ASAP7_75t_R FILLER_190_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_309 ();
 DECAPx4_ASAP7_75t_R FILLER_190_318 ();
 DECAPx2_ASAP7_75t_R FILLER_190_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_338 ();
 DECAPx2_ASAP7_75t_R FILLER_190_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_362 ();
 DECAPx6_ASAP7_75t_R FILLER_190_394 ();
 DECAPx1_ASAP7_75t_R FILLER_190_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_438 ();
 DECAPx6_ASAP7_75t_R FILLER_190_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_461 ();
 DECAPx4_ASAP7_75t_R FILLER_190_464 ();
 FILLER_ASAP7_75t_R FILLER_190_474 ();
 DECAPx2_ASAP7_75t_R FILLER_190_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_489 ();
 DECAPx10_ASAP7_75t_R FILLER_190_496 ();
 DECAPx10_ASAP7_75t_R FILLER_190_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_559 ();
 DECAPx6_ASAP7_75t_R FILLER_190_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_611 ();
 FILLER_ASAP7_75t_R FILLER_190_626 ();
 DECAPx6_ASAP7_75t_R FILLER_190_642 ();
 FILLER_ASAP7_75t_R FILLER_190_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_661 ();
 DECAPx6_ASAP7_75t_R FILLER_190_682 ();
 FILLERxp5_ASAP7_75t_R FILLER_190_696 ();
 DECAPx10_ASAP7_75t_R FILLER_190_726 ();
 DECAPx10_ASAP7_75t_R FILLER_190_748 ();
 DECAPx4_ASAP7_75t_R FILLER_190_770 ();
 FILLER_ASAP7_75t_R FILLER_190_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_796 ();
 FILLER_ASAP7_75t_R FILLER_190_820 ();
 FILLER_ASAP7_75t_R FILLER_190_825 ();
 DECAPx2_ASAP7_75t_R FILLER_190_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_190_905 ();
 DECAPx10_ASAP7_75t_R FILLER_191_7 ();
 DECAPx10_ASAP7_75t_R FILLER_191_29 ();
 DECAPx10_ASAP7_75t_R FILLER_191_51 ();
 DECAPx10_ASAP7_75t_R FILLER_191_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_95 ();
 DECAPx1_ASAP7_75t_R FILLER_191_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_103 ();
 DECAPx1_ASAP7_75t_R FILLER_191_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_114 ();
 DECAPx2_ASAP7_75t_R FILLER_191_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_147 ();
 DECAPx1_ASAP7_75t_R FILLER_191_154 ();
 DECAPx4_ASAP7_75t_R FILLER_191_161 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_186 ();
 DECAPx10_ASAP7_75t_R FILLER_191_223 ();
 DECAPx10_ASAP7_75t_R FILLER_191_245 ();
 DECAPx1_ASAP7_75t_R FILLER_191_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_271 ();
 DECAPx1_ASAP7_75t_R FILLER_191_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_289 ();
 DECAPx6_ASAP7_75t_R FILLER_191_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_318 ();
 DECAPx6_ASAP7_75t_R FILLER_191_325 ();
 DECAPx1_ASAP7_75t_R FILLER_191_345 ();
 DECAPx1_ASAP7_75t_R FILLER_191_355 ();
 DECAPx1_ASAP7_75t_R FILLER_191_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_383 ();
 FILLER_ASAP7_75t_R FILLER_191_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_447 ();
 DECAPx2_ASAP7_75t_R FILLER_191_458 ();
 DECAPx6_ASAP7_75t_R FILLER_191_480 ();
 DECAPx1_ASAP7_75t_R FILLER_191_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_511 ();
 DECAPx1_ASAP7_75t_R FILLER_191_528 ();
 DECAPx10_ASAP7_75t_R FILLER_191_553 ();
 DECAPx2_ASAP7_75t_R FILLER_191_575 ();
 DECAPx1_ASAP7_75t_R FILLER_191_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_612 ();
 DECAPx10_ASAP7_75t_R FILLER_191_628 ();
 DECAPx4_ASAP7_75t_R FILLER_191_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_732 ();
 DECAPx6_ASAP7_75t_R FILLER_191_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_755 ();
 DECAPx6_ASAP7_75t_R FILLER_191_763 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_793 ();
 DECAPx1_ASAP7_75t_R FILLER_191_803 ();
 FILLER_ASAP7_75t_R FILLER_191_856 ();
 DECAPx2_ASAP7_75t_R FILLER_191_874 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_191_880 ();
 FILLER_ASAP7_75t_R FILLER_191_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_191_933 ();
 DECAPx10_ASAP7_75t_R FILLER_192_2 ();
 DECAPx10_ASAP7_75t_R FILLER_192_24 ();
 DECAPx10_ASAP7_75t_R FILLER_192_46 ();
 DECAPx10_ASAP7_75t_R FILLER_192_68 ();
 DECAPx6_ASAP7_75t_R FILLER_192_90 ();
 DECAPx2_ASAP7_75t_R FILLER_192_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_110 ();
 FILLER_ASAP7_75t_R FILLER_192_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_228 ();
 DECAPx10_ASAP7_75t_R FILLER_192_237 ();
 DECAPx6_ASAP7_75t_R FILLER_192_259 ();
 DECAPx1_ASAP7_75t_R FILLER_192_273 ();
 DECAPx1_ASAP7_75t_R FILLER_192_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_328 ();
 DECAPx6_ASAP7_75t_R FILLER_192_355 ();
 FILLER_ASAP7_75t_R FILLER_192_369 ();
 DECAPx6_ASAP7_75t_R FILLER_192_377 ();
 DECAPx1_ASAP7_75t_R FILLER_192_391 ();
 DECAPx6_ASAP7_75t_R FILLER_192_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_417 ();
 DECAPx1_ASAP7_75t_R FILLER_192_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_461 ();
 DECAPx4_ASAP7_75t_R FILLER_192_464 ();
 FILLER_ASAP7_75t_R FILLER_192_474 ();
 DECAPx10_ASAP7_75t_R FILLER_192_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_510 ();
 DECAPx2_ASAP7_75t_R FILLER_192_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_533 ();
 DECAPx1_ASAP7_75t_R FILLER_192_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_570 ();
 DECAPx10_ASAP7_75t_R FILLER_192_592 ();
 DECAPx10_ASAP7_75t_R FILLER_192_614 ();
 DECAPx2_ASAP7_75t_R FILLER_192_636 ();
 FILLER_ASAP7_75t_R FILLER_192_642 ();
 DECAPx10_ASAP7_75t_R FILLER_192_652 ();
 DECAPx4_ASAP7_75t_R FILLER_192_674 ();
 DECAPx10_ASAP7_75t_R FILLER_192_691 ();
 DECAPx1_ASAP7_75t_R FILLER_192_713 ();
 DECAPx1_ASAP7_75t_R FILLER_192_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_779 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_787 ();
 DECAPx4_ASAP7_75t_R FILLER_192_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_192_835 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_869 ();
 DECAPx2_ASAP7_75t_R FILLER_192_878 ();
 FILLER_ASAP7_75t_R FILLER_192_884 ();
 FILLER_ASAP7_75t_R FILLER_192_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_192_933 ();
 DECAPx10_ASAP7_75t_R FILLER_193_7 ();
 DECAPx10_ASAP7_75t_R FILLER_193_29 ();
 DECAPx10_ASAP7_75t_R FILLER_193_51 ();
 DECAPx6_ASAP7_75t_R FILLER_193_73 ();
 DECAPx2_ASAP7_75t_R FILLER_193_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_99 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_103 ();
 DECAPx2_ASAP7_75t_R FILLER_193_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_134 ();
 FILLER_ASAP7_75t_R FILLER_193_141 ();
 DECAPx1_ASAP7_75t_R FILLER_193_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_153 ();
 DECAPx4_ASAP7_75t_R FILLER_193_157 ();
 DECAPx4_ASAP7_75t_R FILLER_193_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_219 ();
 DECAPx10_ASAP7_75t_R FILLER_193_249 ();
 DECAPx2_ASAP7_75t_R FILLER_193_271 ();
 FILLER_ASAP7_75t_R FILLER_193_277 ();
 DECAPx2_ASAP7_75t_R FILLER_193_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_333 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_340 ();
 DECAPx10_ASAP7_75t_R FILLER_193_346 ();
 DECAPx10_ASAP7_75t_R FILLER_193_368 ();
 DECAPx2_ASAP7_75t_R FILLER_193_390 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_396 ();
 DECAPx6_ASAP7_75t_R FILLER_193_407 ();
 DECAPx2_ASAP7_75t_R FILLER_193_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_427 ();
 DECAPx6_ASAP7_75t_R FILLER_193_431 ();
 DECAPx2_ASAP7_75t_R FILLER_193_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_460 ();
 DECAPx6_ASAP7_75t_R FILLER_193_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_483 ();
 DECAPx10_ASAP7_75t_R FILLER_193_498 ();
 DECAPx10_ASAP7_75t_R FILLER_193_520 ();
 FILLER_ASAP7_75t_R FILLER_193_550 ();
 DECAPx2_ASAP7_75t_R FILLER_193_555 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_561 ();
 DECAPx10_ASAP7_75t_R FILLER_193_578 ();
 DECAPx10_ASAP7_75t_R FILLER_193_600 ();
 DECAPx1_ASAP7_75t_R FILLER_193_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_626 ();
 FILLER_ASAP7_75t_R FILLER_193_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_641 ();
 DECAPx6_ASAP7_75t_R FILLER_193_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_674 ();
 DECAPx4_ASAP7_75t_R FILLER_193_687 ();
 FILLER_ASAP7_75t_R FILLER_193_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_713 ();
 DECAPx1_ASAP7_75t_R FILLER_193_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_760 ();
 FILLER_ASAP7_75t_R FILLER_193_768 ();
 DECAPx10_ASAP7_75t_R FILLER_193_777 ();
 DECAPx2_ASAP7_75t_R FILLER_193_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_805 ();
 DECAPx10_ASAP7_75t_R FILLER_193_811 ();
 DECAPx2_ASAP7_75t_R FILLER_193_833 ();
 FILLER_ASAP7_75t_R FILLER_193_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_848 ();
 DECAPx10_ASAP7_75t_R FILLER_193_865 ();
 DECAPx4_ASAP7_75t_R FILLER_193_887 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_897 ();
 DECAPx2_ASAP7_75t_R FILLER_193_903 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_193_909 ();
 FILLERxp5_ASAP7_75t_R FILLER_193_933 ();
 DECAPx10_ASAP7_75t_R FILLER_194_2 ();
 DECAPx10_ASAP7_75t_R FILLER_194_24 ();
 DECAPx10_ASAP7_75t_R FILLER_194_46 ();
 DECAPx6_ASAP7_75t_R FILLER_194_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_82 ();
 DECAPx10_ASAP7_75t_R FILLER_194_111 ();
 DECAPx10_ASAP7_75t_R FILLER_194_133 ();
 DECAPx10_ASAP7_75t_R FILLER_194_155 ();
 DECAPx6_ASAP7_75t_R FILLER_194_177 ();
 DECAPx2_ASAP7_75t_R FILLER_194_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_197 ();
 DECAPx10_ASAP7_75t_R FILLER_194_201 ();
 DECAPx1_ASAP7_75t_R FILLER_194_223 ();
 FILLER_ASAP7_75t_R FILLER_194_233 ();
 DECAPx1_ASAP7_75t_R FILLER_194_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_242 ();
 DECAPx1_ASAP7_75t_R FILLER_194_255 ();
 DECAPx6_ASAP7_75t_R FILLER_194_273 ();
 DECAPx1_ASAP7_75t_R FILLER_194_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_291 ();
 DECAPx2_ASAP7_75t_R FILLER_194_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_301 ();
 DECAPx10_ASAP7_75t_R FILLER_194_310 ();
 DECAPx10_ASAP7_75t_R FILLER_194_332 ();
 DECAPx2_ASAP7_75t_R FILLER_194_354 ();
 FILLER_ASAP7_75t_R FILLER_194_360 ();
 DECAPx2_ASAP7_75t_R FILLER_194_394 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_400 ();
 FILLER_ASAP7_75t_R FILLER_194_419 ();
 DECAPx6_ASAP7_75t_R FILLER_194_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_194_442 ();
 DECAPx2_ASAP7_75t_R FILLER_194_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_461 ();
 DECAPx10_ASAP7_75t_R FILLER_194_464 ();
 FILLER_ASAP7_75t_R FILLER_194_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_517 ();
 DECAPx4_ASAP7_75t_R FILLER_194_525 ();
 FILLER_ASAP7_75t_R FILLER_194_535 ();
 DECAPx4_ASAP7_75t_R FILLER_194_563 ();
 DECAPx4_ASAP7_75t_R FILLER_194_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_591 ();
 DECAPx2_ASAP7_75t_R FILLER_194_596 ();
 DECAPx1_ASAP7_75t_R FILLER_194_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_615 ();
 DECAPx10_ASAP7_75t_R FILLER_194_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_725 ();
 FILLER_ASAP7_75t_R FILLER_194_735 ();
 DECAPx1_ASAP7_75t_R FILLER_194_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_783 ();
 DECAPx10_ASAP7_75t_R FILLER_194_792 ();
 DECAPx2_ASAP7_75t_R FILLER_194_814 ();
 FILLER_ASAP7_75t_R FILLER_194_820 ();
 DECAPx4_ASAP7_75t_R FILLER_194_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_846 ();
 DECAPx2_ASAP7_75t_R FILLER_194_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_860 ();
 DECAPx1_ASAP7_75t_R FILLER_194_866 ();
 DECAPx2_ASAP7_75t_R FILLER_194_886 ();
 FILLER_ASAP7_75t_R FILLER_194_892 ();
 DECAPx1_ASAP7_75t_R FILLER_194_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_905 ();
 DECAPx2_ASAP7_75t_R FILLER_194_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_194_933 ();
 DECAPx10_ASAP7_75t_R FILLER_195_7 ();
 DECAPx10_ASAP7_75t_R FILLER_195_29 ();
 DECAPx10_ASAP7_75t_R FILLER_195_51 ();
 DECAPx6_ASAP7_75t_R FILLER_195_73 ();
 FILLER_ASAP7_75t_R FILLER_195_87 ();
 DECAPx10_ASAP7_75t_R FILLER_195_95 ();
 DECAPx10_ASAP7_75t_R FILLER_195_117 ();
 DECAPx10_ASAP7_75t_R FILLER_195_139 ();
 DECAPx10_ASAP7_75t_R FILLER_195_161 ();
 DECAPx10_ASAP7_75t_R FILLER_195_183 ();
 DECAPx10_ASAP7_75t_R FILLER_195_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_227 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_234 ();
 DECAPx2_ASAP7_75t_R FILLER_195_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_291 ();
 DECAPx10_ASAP7_75t_R FILLER_195_308 ();
 DECAPx4_ASAP7_75t_R FILLER_195_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_352 ();
 DECAPx2_ASAP7_75t_R FILLER_195_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_410 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_433 ();
 DECAPx4_ASAP7_75t_R FILLER_195_462 ();
 DECAPx6_ASAP7_75t_R FILLER_195_478 ();
 FILLER_ASAP7_75t_R FILLER_195_492 ();
 FILLER_ASAP7_75t_R FILLER_195_500 ();
 FILLER_ASAP7_75t_R FILLER_195_505 ();
 DECAPx2_ASAP7_75t_R FILLER_195_519 ();
 DECAPx4_ASAP7_75t_R FILLER_195_531 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_552 ();
 DECAPx6_ASAP7_75t_R FILLER_195_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_596 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_195_605 ();
 DECAPx2_ASAP7_75t_R FILLER_195_626 ();
 DECAPx2_ASAP7_75t_R FILLER_195_638 ();
 FILLER_ASAP7_75t_R FILLER_195_644 ();
 DECAPx2_ASAP7_75t_R FILLER_195_652 ();
 FILLER_ASAP7_75t_R FILLER_195_658 ();
 DECAPx6_ASAP7_75t_R FILLER_195_672 ();
 DECAPx1_ASAP7_75t_R FILLER_195_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_690 ();
 DECAPx10_ASAP7_75t_R FILLER_195_700 ();
 DECAPx10_ASAP7_75t_R FILLER_195_722 ();
 DECAPx6_ASAP7_75t_R FILLER_195_744 ();
 DECAPx2_ASAP7_75t_R FILLER_195_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_764 ();
 DECAPx2_ASAP7_75t_R FILLER_195_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_195_777 ();
 DECAPx2_ASAP7_75t_R FILLER_195_809 ();
 DECAPx2_ASAP7_75t_R FILLER_195_841 ();
 FILLER_ASAP7_75t_R FILLER_195_932 ();
 DECAPx10_ASAP7_75t_R FILLER_196_7 ();
 DECAPx10_ASAP7_75t_R FILLER_196_29 ();
 DECAPx10_ASAP7_75t_R FILLER_196_51 ();
 DECAPx10_ASAP7_75t_R FILLER_196_73 ();
 DECAPx1_ASAP7_75t_R FILLER_196_101 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_105 ();
 DECAPx6_ASAP7_75t_R FILLER_196_112 ();
 DECAPx2_ASAP7_75t_R FILLER_196_126 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_138 ();
 DECAPx2_ASAP7_75t_R FILLER_196_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_180 ();
 DECAPx2_ASAP7_75t_R FILLER_196_209 ();
 FILLER_ASAP7_75t_R FILLER_196_215 ();
 FILLER_ASAP7_75t_R FILLER_196_223 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_254 ();
 DECAPx1_ASAP7_75t_R FILLER_196_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_273 ();
 DECAPx4_ASAP7_75t_R FILLER_196_300 ();
 FILLER_ASAP7_75t_R FILLER_196_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_318 ();
 FILLER_ASAP7_75t_R FILLER_196_331 ();
 DECAPx1_ASAP7_75t_R FILLER_196_373 ();
 DECAPx1_ASAP7_75t_R FILLER_196_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_384 ();
 DECAPx1_ASAP7_75t_R FILLER_196_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_395 ();
 DECAPx6_ASAP7_75t_R FILLER_196_399 ();
 FILLER_ASAP7_75t_R FILLER_196_413 ();
 FILLER_ASAP7_75t_R FILLER_196_435 ();
 DECAPx1_ASAP7_75t_R FILLER_196_445 ();
 FILLER_ASAP7_75t_R FILLER_196_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_464 ();
 DECAPx10_ASAP7_75t_R FILLER_196_491 ();
 DECAPx10_ASAP7_75t_R FILLER_196_513 ();
 DECAPx2_ASAP7_75t_R FILLER_196_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_547 ();
 DECAPx1_ASAP7_75t_R FILLER_196_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_559 ();
 FILLER_ASAP7_75t_R FILLER_196_570 ();
 DECAPx2_ASAP7_75t_R FILLER_196_600 ();
 FILLER_ASAP7_75t_R FILLER_196_606 ();
 DECAPx6_ASAP7_75t_R FILLER_196_614 ();
 FILLERxp5_ASAP7_75t_R FILLER_196_628 ();
 DECAPx10_ASAP7_75t_R FILLER_196_638 ();
 FILLER_ASAP7_75t_R FILLER_196_660 ();
 DECAPx10_ASAP7_75t_R FILLER_196_677 ();
 DECAPx10_ASAP7_75t_R FILLER_196_699 ();
 DECAPx10_ASAP7_75t_R FILLER_196_721 ();
 DECAPx10_ASAP7_75t_R FILLER_196_743 ();
 DECAPx10_ASAP7_75t_R FILLER_196_765 ();
 DECAPx2_ASAP7_75t_R FILLER_196_787 ();
 DECAPx6_ASAP7_75t_R FILLER_196_796 ();
 DECAPx1_ASAP7_75t_R FILLER_196_810 ();
 FILLER_ASAP7_75t_R FILLER_196_835 ();
 DECAPx2_ASAP7_75t_R FILLER_196_843 ();
 DECAPx2_ASAP7_75t_R FILLER_196_855 ();
 DECAPx2_ASAP7_75t_R FILLER_196_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_870 ();
 FILLER_ASAP7_75t_R FILLER_196_883 ();
 DECAPx2_ASAP7_75t_R FILLER_196_890 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_196_896 ();
 DECAPx10_ASAP7_75t_R FILLER_197_2 ();
 DECAPx10_ASAP7_75t_R FILLER_197_24 ();
 DECAPx10_ASAP7_75t_R FILLER_197_46 ();
 DECAPx10_ASAP7_75t_R FILLER_197_68 ();
 FILLER_ASAP7_75t_R FILLER_197_90 ();
 FILLER_ASAP7_75t_R FILLER_197_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_192 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_238 ();
 DECAPx10_ASAP7_75t_R FILLER_197_242 ();
 DECAPx4_ASAP7_75t_R FILLER_197_264 ();
 DECAPx6_ASAP7_75t_R FILLER_197_282 ();
 DECAPx1_ASAP7_75t_R FILLER_197_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_300 ();
 DECAPx2_ASAP7_75t_R FILLER_197_339 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_345 ();
 DECAPx10_ASAP7_75t_R FILLER_197_382 ();
 DECAPx2_ASAP7_75t_R FILLER_197_404 ();
 FILLER_ASAP7_75t_R FILLER_197_410 ();
 DECAPx10_ASAP7_75t_R FILLER_197_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_460 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_467 ();
 DECAPx2_ASAP7_75t_R FILLER_197_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_486 ();
 DECAPx10_ASAP7_75t_R FILLER_197_500 ();
 DECAPx2_ASAP7_75t_R FILLER_197_522 ();
 FILLER_ASAP7_75t_R FILLER_197_528 ();
 DECAPx10_ASAP7_75t_R FILLER_197_538 ();
 DECAPx4_ASAP7_75t_R FILLER_197_570 ();
 FILLER_ASAP7_75t_R FILLER_197_580 ();
 DECAPx10_ASAP7_75t_R FILLER_197_610 ();
 DECAPx6_ASAP7_75t_R FILLER_197_632 ();
 DECAPx1_ASAP7_75t_R FILLER_197_646 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_650 ();
 DECAPx4_ASAP7_75t_R FILLER_197_660 ();
 DECAPx10_ASAP7_75t_R FILLER_197_686 ();
 DECAPx1_ASAP7_75t_R FILLER_197_708 ();
 DECAPx4_ASAP7_75t_R FILLER_197_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_728 ();
 DECAPx2_ASAP7_75t_R FILLER_197_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_197_754 ();
 DECAPx6_ASAP7_75t_R FILLER_197_762 ();
 DECAPx1_ASAP7_75t_R FILLER_197_776 ();
 DECAPx2_ASAP7_75t_R FILLER_197_792 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_197_798 ();
 DECAPx2_ASAP7_75t_R FILLER_197_826 ();
 DECAPx10_ASAP7_75t_R FILLER_197_847 ();
 DECAPx10_ASAP7_75t_R FILLER_197_869 ();
 DECAPx6_ASAP7_75t_R FILLER_197_891 ();
 DECAPx1_ASAP7_75t_R FILLER_197_905 ();
 FILLER_ASAP7_75t_R FILLER_197_927 ();
 DECAPx10_ASAP7_75t_R FILLER_198_2 ();
 DECAPx10_ASAP7_75t_R FILLER_198_24 ();
 DECAPx10_ASAP7_75t_R FILLER_198_46 ();
 DECAPx10_ASAP7_75t_R FILLER_198_68 ();
 DECAPx2_ASAP7_75t_R FILLER_198_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_96 ();
 FILLER_ASAP7_75t_R FILLER_198_131 ();
 DECAPx1_ASAP7_75t_R FILLER_198_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_145 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_166 ();
 DECAPx2_ASAP7_75t_R FILLER_198_175 ();
 DECAPx1_ASAP7_75t_R FILLER_198_184 ();
 DECAPx4_ASAP7_75t_R FILLER_198_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_204 ();
 FILLER_ASAP7_75t_R FILLER_198_211 ();
 DECAPx10_ASAP7_75t_R FILLER_198_225 ();
 DECAPx10_ASAP7_75t_R FILLER_198_247 ();
 DECAPx10_ASAP7_75t_R FILLER_198_269 ();
 DECAPx6_ASAP7_75t_R FILLER_198_291 ();
 FILLER_ASAP7_75t_R FILLER_198_305 ();
 FILLER_ASAP7_75t_R FILLER_198_313 ();
 FILLER_ASAP7_75t_R FILLER_198_318 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_323 ();
 DECAPx2_ASAP7_75t_R FILLER_198_330 ();
 DECAPx2_ASAP7_75t_R FILLER_198_348 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_354 ();
 DECAPx1_ASAP7_75t_R FILLER_198_361 ();
 DECAPx2_ASAP7_75t_R FILLER_198_391 ();
 DECAPx10_ASAP7_75t_R FILLER_198_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_425 ();
 DECAPx2_ASAP7_75t_R FILLER_198_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_435 ();
 DECAPx4_ASAP7_75t_R FILLER_198_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_461 ();
 DECAPx10_ASAP7_75t_R FILLER_198_464 ();
 FILLER_ASAP7_75t_R FILLER_198_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_494 ();
 DECAPx4_ASAP7_75t_R FILLER_198_510 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_520 ();
 DECAPx2_ASAP7_75t_R FILLER_198_541 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_198_555 ();
 DECAPx2_ASAP7_75t_R FILLER_198_565 ();
 FILLER_ASAP7_75t_R FILLER_198_571 ();
 DECAPx6_ASAP7_75t_R FILLER_198_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_608 ();
 DECAPx10_ASAP7_75t_R FILLER_198_615 ();
 DECAPx6_ASAP7_75t_R FILLER_198_664 ();
 FILLER_ASAP7_75t_R FILLER_198_678 ();
 FILLER_ASAP7_75t_R FILLER_198_690 ();
 DECAPx1_ASAP7_75t_R FILLER_198_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_726 ();
 DECAPx4_ASAP7_75t_R FILLER_198_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_198_774 ();
 DECAPx2_ASAP7_75t_R FILLER_198_876 ();
 FILLER_ASAP7_75t_R FILLER_198_882 ();
 DECAPx10_ASAP7_75t_R FILLER_199_7 ();
 DECAPx10_ASAP7_75t_R FILLER_199_29 ();
 DECAPx10_ASAP7_75t_R FILLER_199_51 ();
 DECAPx10_ASAP7_75t_R FILLER_199_73 ();
 DECAPx1_ASAP7_75t_R FILLER_199_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_113 ();
 DECAPx10_ASAP7_75t_R FILLER_199_143 ();
 DECAPx2_ASAP7_75t_R FILLER_199_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_171 ();
 DECAPx6_ASAP7_75t_R FILLER_199_180 ();
 FILLER_ASAP7_75t_R FILLER_199_194 ();
 DECAPx4_ASAP7_75t_R FILLER_199_222 ();
 FILLER_ASAP7_75t_R FILLER_199_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_240 ();
 DECAPx10_ASAP7_75t_R FILLER_199_244 ();
 DECAPx4_ASAP7_75t_R FILLER_199_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_295 ();
 DECAPx6_ASAP7_75t_R FILLER_199_306 ();
 DECAPx2_ASAP7_75t_R FILLER_199_320 ();
 DECAPx6_ASAP7_75t_R FILLER_199_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_371 ();
 FILLER_ASAP7_75t_R FILLER_199_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_411 ();
 DECAPx6_ASAP7_75t_R FILLER_199_417 ();
 DECAPx6_ASAP7_75t_R FILLER_199_477 ();
 DECAPx1_ASAP7_75t_R FILLER_199_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_502 ();
 DECAPx1_ASAP7_75t_R FILLER_199_509 ();
 FILLER_ASAP7_75t_R FILLER_199_527 ();
 DECAPx1_ASAP7_75t_R FILLER_199_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_583 ();
 FILLER_ASAP7_75t_R FILLER_199_599 ();
 DECAPx6_ASAP7_75t_R FILLER_199_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_644 ();
 DECAPx10_ASAP7_75t_R FILLER_199_651 ();
 DECAPx6_ASAP7_75t_R FILLER_199_673 ();
 DECAPx1_ASAP7_75t_R FILLER_199_687 ();
 FILLER_ASAP7_75t_R FILLER_199_713 ();
 DECAPx1_ASAP7_75t_R FILLER_199_723 ();
 DECAPx1_ASAP7_75t_R FILLER_199_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_747 ();
 DECAPx1_ASAP7_75t_R FILLER_199_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_777 ();
 DECAPx4_ASAP7_75t_R FILLER_199_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_199_804 ();
 DECAPx4_ASAP7_75t_R FILLER_199_818 ();
 DECAPx2_ASAP7_75t_R FILLER_199_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_199_839 ();
 DECAPx4_ASAP7_75t_R FILLER_199_845 ();
 FILLER_ASAP7_75t_R FILLER_199_927 ();
 DECAPx10_ASAP7_75t_R FILLER_200_2 ();
 DECAPx10_ASAP7_75t_R FILLER_200_24 ();
 DECAPx10_ASAP7_75t_R FILLER_200_46 ();
 DECAPx10_ASAP7_75t_R FILLER_200_68 ();
 DECAPx6_ASAP7_75t_R FILLER_200_90 ();
 FILLER_ASAP7_75t_R FILLER_200_104 ();
 FILLER_ASAP7_75t_R FILLER_200_109 ();
 DECAPx10_ASAP7_75t_R FILLER_200_114 ();
 DECAPx10_ASAP7_75t_R FILLER_200_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_158 ();
 DECAPx1_ASAP7_75t_R FILLER_200_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_166 ();
 DECAPx2_ASAP7_75t_R FILLER_200_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_199 ();
 DECAPx1_ASAP7_75t_R FILLER_200_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_210 ();
 DECAPx4_ASAP7_75t_R FILLER_200_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_253 ();
 FILLER_ASAP7_75t_R FILLER_200_287 ();
 DECAPx4_ASAP7_75t_R FILLER_200_315 ();
 FILLER_ASAP7_75t_R FILLER_200_325 ();
 DECAPx2_ASAP7_75t_R FILLER_200_337 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_343 ();
 DECAPx10_ASAP7_75t_R FILLER_200_349 ();
 DECAPx4_ASAP7_75t_R FILLER_200_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_381 ();
 FILLER_ASAP7_75t_R FILLER_200_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_424 ();
 FILLER_ASAP7_75t_R FILLER_200_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_442 ();
 DECAPx2_ASAP7_75t_R FILLER_200_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_461 ();
 DECAPx4_ASAP7_75t_R FILLER_200_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_474 ();
 DECAPx6_ASAP7_75t_R FILLER_200_481 ();
 DECAPx1_ASAP7_75t_R FILLER_200_495 ();
 DECAPx1_ASAP7_75t_R FILLER_200_506 ();
 FILLER_ASAP7_75t_R FILLER_200_523 ();
 DECAPx6_ASAP7_75t_R FILLER_200_532 ();
 DECAPx4_ASAP7_75t_R FILLER_200_563 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_573 ();
 DECAPx6_ASAP7_75t_R FILLER_200_583 ();
 DECAPx2_ASAP7_75t_R FILLER_200_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_603 ();
 DECAPx1_ASAP7_75t_R FILLER_200_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_617 ();
 DECAPx4_ASAP7_75t_R FILLER_200_650 ();
 FILLER_ASAP7_75t_R FILLER_200_660 ();
 DECAPx2_ASAP7_75t_R FILLER_200_677 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_683 ();
 FILLER_ASAP7_75t_R FILLER_200_717 ();
 DECAPx4_ASAP7_75t_R FILLER_200_732 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_755 ();
 DECAPx1_ASAP7_75t_R FILLER_200_764 ();
 DECAPx10_ASAP7_75t_R FILLER_200_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_815 ();
 DECAPx4_ASAP7_75t_R FILLER_200_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_835 ();
 DECAPx10_ASAP7_75t_R FILLER_200_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_200_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_200_910 ();
 FILLER_ASAP7_75t_R FILLER_200_922 ();
 DECAPx10_ASAP7_75t_R FILLER_201_2 ();
 DECAPx10_ASAP7_75t_R FILLER_201_24 ();
 DECAPx10_ASAP7_75t_R FILLER_201_46 ();
 DECAPx10_ASAP7_75t_R FILLER_201_68 ();
 DECAPx10_ASAP7_75t_R FILLER_201_90 ();
 DECAPx10_ASAP7_75t_R FILLER_201_112 ();
 DECAPx4_ASAP7_75t_R FILLER_201_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_144 ();
 FILLER_ASAP7_75t_R FILLER_201_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_185 ();
 DECAPx10_ASAP7_75t_R FILLER_201_192 ();
 DECAPx6_ASAP7_75t_R FILLER_201_214 ();
 FILLER_ASAP7_75t_R FILLER_201_228 ();
 DECAPx4_ASAP7_75t_R FILLER_201_236 ();
 DECAPx2_ASAP7_75t_R FILLER_201_278 ();
 FILLER_ASAP7_75t_R FILLER_201_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_301 ();
 DECAPx10_ASAP7_75t_R FILLER_201_314 ();
 FILLER_ASAP7_75t_R FILLER_201_336 ();
 DECAPx2_ASAP7_75t_R FILLER_201_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_376 ();
 DECAPx2_ASAP7_75t_R FILLER_201_380 ();
 FILLER_ASAP7_75t_R FILLER_201_407 ();
 DECAPx2_ASAP7_75t_R FILLER_201_435 ();
 DECAPx2_ASAP7_75t_R FILLER_201_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_483 ();
 DECAPx4_ASAP7_75t_R FILLER_201_492 ();
 DECAPx1_ASAP7_75t_R FILLER_201_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_519 ();
 DECAPx10_ASAP7_75t_R FILLER_201_530 ();
 DECAPx10_ASAP7_75t_R FILLER_201_552 ();
 DECAPx4_ASAP7_75t_R FILLER_201_574 ();
 DECAPx6_ASAP7_75t_R FILLER_201_592 ();
 FILLER_ASAP7_75t_R FILLER_201_606 ();
 DECAPx2_ASAP7_75t_R FILLER_201_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_619 ();
 DECAPx6_ASAP7_75t_R FILLER_201_641 ();
 DECAPx2_ASAP7_75t_R FILLER_201_655 ();
 DECAPx4_ASAP7_75t_R FILLER_201_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_694 ();
 DECAPx1_ASAP7_75t_R FILLER_201_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_703 ();
 DECAPx4_ASAP7_75t_R FILLER_201_710 ();
 DECAPx6_ASAP7_75t_R FILLER_201_726 ();
 DECAPx1_ASAP7_75t_R FILLER_201_740 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_744 ();
 DECAPx6_ASAP7_75t_R FILLER_201_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_201_771 ();
 DECAPx10_ASAP7_75t_R FILLER_201_788 ();
 DECAPx1_ASAP7_75t_R FILLER_201_810 ();
 DECAPx10_ASAP7_75t_R FILLER_201_840 ();
 DECAPx6_ASAP7_75t_R FILLER_201_862 ();
 DECAPx1_ASAP7_75t_R FILLER_201_907 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_201_922 ();
 FILLER_ASAP7_75t_R FILLER_201_932 ();
 DECAPx10_ASAP7_75t_R FILLER_202_7 ();
 DECAPx10_ASAP7_75t_R FILLER_202_29 ();
 DECAPx10_ASAP7_75t_R FILLER_202_51 ();
 DECAPx10_ASAP7_75t_R FILLER_202_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_95 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_104 ();
 DECAPx10_ASAP7_75t_R FILLER_202_113 ();
 DECAPx2_ASAP7_75t_R FILLER_202_135 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_141 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_183 ();
 DECAPx2_ASAP7_75t_R FILLER_202_192 ();
 FILLER_ASAP7_75t_R FILLER_202_198 ();
 DECAPx6_ASAP7_75t_R FILLER_202_216 ();
 DECAPx2_ASAP7_75t_R FILLER_202_236 ();
 DECAPx2_ASAP7_75t_R FILLER_202_245 ();
 DECAPx1_ASAP7_75t_R FILLER_202_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_271 ();
 DECAPx2_ASAP7_75t_R FILLER_202_279 ();
 FILLER_ASAP7_75t_R FILLER_202_285 ();
 DECAPx6_ASAP7_75t_R FILLER_202_293 ();
 DECAPx2_ASAP7_75t_R FILLER_202_307 ();
 DECAPx6_ASAP7_75t_R FILLER_202_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_341 ();
 DECAPx2_ASAP7_75t_R FILLER_202_357 ();
 DECAPx10_ASAP7_75t_R FILLER_202_389 ();
 DECAPx1_ASAP7_75t_R FILLER_202_411 ();
 FILLER_ASAP7_75t_R FILLER_202_422 ();
 DECAPx1_ASAP7_75t_R FILLER_202_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_431 ();
 DECAPx1_ASAP7_75t_R FILLER_202_458 ();
 DECAPx4_ASAP7_75t_R FILLER_202_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_481 ();
 DECAPx4_ASAP7_75t_R FILLER_202_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_508 ();
 DECAPx4_ASAP7_75t_R FILLER_202_517 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_202_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_536 ();
 DECAPx4_ASAP7_75t_R FILLER_202_551 ();
 FILLER_ASAP7_75t_R FILLER_202_561 ();
 DECAPx4_ASAP7_75t_R FILLER_202_570 ();
 DECAPx4_ASAP7_75t_R FILLER_202_587 ();
 FILLER_ASAP7_75t_R FILLER_202_597 ();
 DECAPx6_ASAP7_75t_R FILLER_202_606 ();
 DECAPx1_ASAP7_75t_R FILLER_202_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_624 ();
 FILLER_ASAP7_75t_R FILLER_202_628 ();
 DECAPx10_ASAP7_75t_R FILLER_202_648 ();
 DECAPx10_ASAP7_75t_R FILLER_202_676 ();
 DECAPx10_ASAP7_75t_R FILLER_202_698 ();
 DECAPx10_ASAP7_75t_R FILLER_202_720 ();
 DECAPx10_ASAP7_75t_R FILLER_202_760 ();
 DECAPx2_ASAP7_75t_R FILLER_202_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_202_788 ();
 FILLER_ASAP7_75t_R FILLER_202_802 ();
 DECAPx6_ASAP7_75t_R FILLER_202_807 ();
 FILLER_ASAP7_75t_R FILLER_202_827 ();
 DECAPx2_ASAP7_75t_R FILLER_202_832 ();
 FILLER_ASAP7_75t_R FILLER_202_838 ();
 FILLER_ASAP7_75t_R FILLER_202_853 ();
 FILLER_ASAP7_75t_R FILLER_202_880 ();
 FILLER_ASAP7_75t_R FILLER_202_892 ();
 DECAPx10_ASAP7_75t_R FILLER_203_12 ();
 DECAPx10_ASAP7_75t_R FILLER_203_34 ();
 DECAPx10_ASAP7_75t_R FILLER_203_56 ();
 DECAPx6_ASAP7_75t_R FILLER_203_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_92 ();
 DECAPx1_ASAP7_75t_R FILLER_203_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_137 ();
 DECAPx1_ASAP7_75t_R FILLER_203_146 ();
 DECAPx6_ASAP7_75t_R FILLER_203_173 ();
 DECAPx2_ASAP7_75t_R FILLER_203_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_193 ();
 DECAPx6_ASAP7_75t_R FILLER_203_254 ();
 DECAPx2_ASAP7_75t_R FILLER_203_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_274 ();
 DECAPx6_ASAP7_75t_R FILLER_203_290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_304 ();
 DECAPx1_ASAP7_75t_R FILLER_203_322 ();
 DECAPx10_ASAP7_75t_R FILLER_203_336 ();
 DECAPx2_ASAP7_75t_R FILLER_203_358 ();
 FILLER_ASAP7_75t_R FILLER_203_364 ();
 DECAPx1_ASAP7_75t_R FILLER_203_372 ();
 DECAPx2_ASAP7_75t_R FILLER_203_382 ();
 FILLER_ASAP7_75t_R FILLER_203_388 ();
 DECAPx2_ASAP7_75t_R FILLER_203_414 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_420 ();
 DECAPx6_ASAP7_75t_R FILLER_203_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_443 ();
 DECAPx6_ASAP7_75t_R FILLER_203_449 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_463 ();
 DECAPx4_ASAP7_75t_R FILLER_203_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_484 ();
 DECAPx10_ASAP7_75t_R FILLER_203_491 ();
 DECAPx6_ASAP7_75t_R FILLER_203_513 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_203_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_556 ();
 DECAPx4_ASAP7_75t_R FILLER_203_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_585 ();
 DECAPx10_ASAP7_75t_R FILLER_203_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_629 ();
 DECAPx4_ASAP7_75t_R FILLER_203_639 ();
 FILLER_ASAP7_75t_R FILLER_203_649 ();
 DECAPx2_ASAP7_75t_R FILLER_203_667 ();
 FILLER_ASAP7_75t_R FILLER_203_673 ();
 DECAPx10_ASAP7_75t_R FILLER_203_690 ();
 DECAPx4_ASAP7_75t_R FILLER_203_720 ();
 DECAPx6_ASAP7_75t_R FILLER_203_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_760 ();
 DECAPx4_ASAP7_75t_R FILLER_203_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_788 ();
 DECAPx6_ASAP7_75t_R FILLER_203_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_855 ();
 FILLER_ASAP7_75t_R FILLER_203_890 ();
 FILLER_ASAP7_75t_R FILLER_203_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_203_933 ();
 DECAPx10_ASAP7_75t_R FILLER_204_2 ();
 DECAPx10_ASAP7_75t_R FILLER_204_24 ();
 DECAPx10_ASAP7_75t_R FILLER_204_46 ();
 DECAPx6_ASAP7_75t_R FILLER_204_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_82 ();
 FILLER_ASAP7_75t_R FILLER_204_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_159 ();
 DECAPx1_ASAP7_75t_R FILLER_204_172 ();
 DECAPx4_ASAP7_75t_R FILLER_204_184 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_194 ();
 FILLER_ASAP7_75t_R FILLER_204_224 ();
 FILLER_ASAP7_75t_R FILLER_204_232 ();
 FILLER_ASAP7_75t_R FILLER_204_237 ();
 DECAPx10_ASAP7_75t_R FILLER_204_245 ();
 DECAPx2_ASAP7_75t_R FILLER_204_267 ();
 DECAPx10_ASAP7_75t_R FILLER_204_287 ();
 DECAPx2_ASAP7_75t_R FILLER_204_309 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_350 ();
 DECAPx1_ASAP7_75t_R FILLER_204_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_367 ();
 DECAPx6_ASAP7_75t_R FILLER_204_394 ();
 DECAPx1_ASAP7_75t_R FILLER_204_408 ();
 FILLER_ASAP7_75t_R FILLER_204_424 ();
 DECAPx10_ASAP7_75t_R FILLER_204_433 ();
 DECAPx2_ASAP7_75t_R FILLER_204_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_500 ();
 DECAPx6_ASAP7_75t_R FILLER_204_515 ();
 FILLER_ASAP7_75t_R FILLER_204_529 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_561 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_571 ();
 DECAPx2_ASAP7_75t_R FILLER_204_580 ();
 FILLER_ASAP7_75t_R FILLER_204_586 ();
 DECAPx2_ASAP7_75t_R FILLER_204_595 ();
 DECAPx1_ASAP7_75t_R FILLER_204_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_619 ();
 DECAPx4_ASAP7_75t_R FILLER_204_629 ();
 FILLER_ASAP7_75t_R FILLER_204_639 ();
 DECAPx1_ASAP7_75t_R FILLER_204_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_675 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_204_688 ();
 DECAPx1_ASAP7_75t_R FILLER_204_704 ();
 DECAPx4_ASAP7_75t_R FILLER_204_715 ();
 DECAPx4_ASAP7_75t_R FILLER_204_731 ();
 FILLER_ASAP7_75t_R FILLER_204_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_751 ();
 DECAPx2_ASAP7_75t_R FILLER_204_774 ();
 DECAPx10_ASAP7_75t_R FILLER_204_806 ();
 DECAPx4_ASAP7_75t_R FILLER_204_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_877 ();
 DECAPx1_ASAP7_75t_R FILLER_204_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_204_892 ();
 DECAPx10_ASAP7_75t_R FILLER_205_2 ();
 DECAPx10_ASAP7_75t_R FILLER_205_24 ();
 DECAPx10_ASAP7_75t_R FILLER_205_46 ();
 DECAPx10_ASAP7_75t_R FILLER_205_68 ();
 DECAPx2_ASAP7_75t_R FILLER_205_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_105 ();
 DECAPx1_ASAP7_75t_R FILLER_205_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_130 ();
 DECAPx2_ASAP7_75t_R FILLER_205_146 ();
 DECAPx2_ASAP7_75t_R FILLER_205_168 ();
 DECAPx2_ASAP7_75t_R FILLER_205_194 ();
 DECAPx1_ASAP7_75t_R FILLER_205_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_253 ();
 DECAPx10_ASAP7_75t_R FILLER_205_262 ();
 DECAPx2_ASAP7_75t_R FILLER_205_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_303 ();
 DECAPx2_ASAP7_75t_R FILLER_205_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_317 ();
 FILLER_ASAP7_75t_R FILLER_205_356 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_380 ();
 DECAPx2_ASAP7_75t_R FILLER_205_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_398 ();
 DECAPx1_ASAP7_75t_R FILLER_205_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_412 ();
 DECAPx10_ASAP7_75t_R FILLER_205_419 ();
 DECAPx1_ASAP7_75t_R FILLER_205_441 ();
 DECAPx6_ASAP7_75t_R FILLER_205_455 ();
 FILLER_ASAP7_75t_R FILLER_205_469 ();
 DECAPx6_ASAP7_75t_R FILLER_205_474 ();
 DECAPx1_ASAP7_75t_R FILLER_205_488 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_502 ();
 DECAPx1_ASAP7_75t_R FILLER_205_511 ();
 DECAPx10_ASAP7_75t_R FILLER_205_529 ();
 DECAPx10_ASAP7_75t_R FILLER_205_551 ();
 DECAPx1_ASAP7_75t_R FILLER_205_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_577 ();
 DECAPx6_ASAP7_75t_R FILLER_205_586 ();
 DECAPx1_ASAP7_75t_R FILLER_205_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_604 ();
 DECAPx1_ASAP7_75t_R FILLER_205_613 ();
 DECAPx10_ASAP7_75t_R FILLER_205_625 ();
 DECAPx1_ASAP7_75t_R FILLER_205_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_651 ();
 DECAPx2_ASAP7_75t_R FILLER_205_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_667 ();
 DECAPx1_ASAP7_75t_R FILLER_205_672 ();
 DECAPx1_ASAP7_75t_R FILLER_205_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_689 ();
 FILLER_ASAP7_75t_R FILLER_205_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_728 ();
 DECAPx2_ASAP7_75t_R FILLER_205_738 ();
 FILLER_ASAP7_75t_R FILLER_205_744 ();
 DECAPx1_ASAP7_75t_R FILLER_205_752 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_764 ();
 DECAPx2_ASAP7_75t_R FILLER_205_788 ();
 DECAPx6_ASAP7_75t_R FILLER_205_797 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_811 ();
 DECAPx2_ASAP7_75t_R FILLER_205_820 ();
 DECAPx2_ASAP7_75t_R FILLER_205_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_842 ();
 FILLER_ASAP7_75t_R FILLER_205_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_855 ();
 DECAPx10_ASAP7_75t_R FILLER_205_861 ();
 DECAPx4_ASAP7_75t_R FILLER_205_883 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_205_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_205_933 ();
 DECAPx10_ASAP7_75t_R FILLER_206_2 ();
 DECAPx10_ASAP7_75t_R FILLER_206_24 ();
 DECAPx10_ASAP7_75t_R FILLER_206_46 ();
 DECAPx10_ASAP7_75t_R FILLER_206_68 ();
 DECAPx6_ASAP7_75t_R FILLER_206_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_104 ();
 DECAPx10_ASAP7_75t_R FILLER_206_108 ();
 DECAPx10_ASAP7_75t_R FILLER_206_130 ();
 DECAPx2_ASAP7_75t_R FILLER_206_152 ();
 DECAPx6_ASAP7_75t_R FILLER_206_164 ();
 DECAPx1_ASAP7_75t_R FILLER_206_178 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_188 ();
 DECAPx1_ASAP7_75t_R FILLER_206_203 ();
 DECAPx2_ASAP7_75t_R FILLER_206_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_228 ();
 DECAPx10_ASAP7_75t_R FILLER_206_237 ();
 FILLER_ASAP7_75t_R FILLER_206_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_267 ();
 DECAPx4_ASAP7_75t_R FILLER_206_274 ();
 DECAPx4_ASAP7_75t_R FILLER_206_328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_338 ();
 FILLER_ASAP7_75t_R FILLER_206_350 ();
 DECAPx10_ASAP7_75t_R FILLER_206_355 ();
 DECAPx2_ASAP7_75t_R FILLER_206_377 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_383 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_419 ();
 DECAPx1_ASAP7_75t_R FILLER_206_432 ();
 DECAPx10_ASAP7_75t_R FILLER_206_472 ();
 DECAPx1_ASAP7_75t_R FILLER_206_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_504 ();
 DECAPx1_ASAP7_75t_R FILLER_206_515 ();
 DECAPx10_ASAP7_75t_R FILLER_206_525 ();
 DECAPx10_ASAP7_75t_R FILLER_206_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_569 ();
 DECAPx1_ASAP7_75t_R FILLER_206_596 ();
 DECAPx1_ASAP7_75t_R FILLER_206_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_627 ();
 FILLER_ASAP7_75t_R FILLER_206_636 ();
 DECAPx10_ASAP7_75t_R FILLER_206_649 ();
 DECAPx2_ASAP7_75t_R FILLER_206_671 ();
 DECAPx6_ASAP7_75t_R FILLER_206_683 ();
 DECAPx2_ASAP7_75t_R FILLER_206_697 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_206_716 ();
 DECAPx1_ASAP7_75t_R FILLER_206_750 ();
 DECAPx1_ASAP7_75t_R FILLER_206_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_765 ();
 DECAPx4_ASAP7_75t_R FILLER_206_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_796 ();
 FILLER_ASAP7_75t_R FILLER_206_815 ();
 DECAPx2_ASAP7_75t_R FILLER_206_843 ();
 DECAPx6_ASAP7_75t_R FILLER_206_862 ();
 DECAPx2_ASAP7_75t_R FILLER_206_876 ();
 DECAPx1_ASAP7_75t_R FILLER_206_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_206_928 ();
 DECAPx10_ASAP7_75t_R FILLER_207_7 ();
 DECAPx10_ASAP7_75t_R FILLER_207_29 ();
 DECAPx10_ASAP7_75t_R FILLER_207_51 ();
 DECAPx10_ASAP7_75t_R FILLER_207_73 ();
 DECAPx10_ASAP7_75t_R FILLER_207_95 ();
 DECAPx2_ASAP7_75t_R FILLER_207_117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_123 ();
 FILLER_ASAP7_75t_R FILLER_207_132 ();
 DECAPx6_ASAP7_75t_R FILLER_207_146 ();
 FILLER_ASAP7_75t_R FILLER_207_160 ();
 DECAPx1_ASAP7_75t_R FILLER_207_168 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_178 ();
 FILLER_ASAP7_75t_R FILLER_207_203 ();
 DECAPx4_ASAP7_75t_R FILLER_207_247 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_264 ();
 DECAPx1_ASAP7_75t_R FILLER_207_277 ();
 DECAPx10_ASAP7_75t_R FILLER_207_299 ();
 DECAPx10_ASAP7_75t_R FILLER_207_321 ();
 DECAPx10_ASAP7_75t_R FILLER_207_343 ();
 DECAPx2_ASAP7_75t_R FILLER_207_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_371 ();
 DECAPx10_ASAP7_75t_R FILLER_207_378 ();
 DECAPx2_ASAP7_75t_R FILLER_207_403 ();
 FILLER_ASAP7_75t_R FILLER_207_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_437 ();
 DECAPx2_ASAP7_75t_R FILLER_207_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_451 ();
 DECAPx6_ASAP7_75t_R FILLER_207_463 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_477 ();
 FILLER_ASAP7_75t_R FILLER_207_485 ();
 DECAPx10_ASAP7_75t_R FILLER_207_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_515 ();
 DECAPx1_ASAP7_75t_R FILLER_207_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_529 ();
 DECAPx2_ASAP7_75t_R FILLER_207_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_543 ();
 DECAPx10_ASAP7_75t_R FILLER_207_565 ();
 DECAPx1_ASAP7_75t_R FILLER_207_587 ();
 DECAPx1_ASAP7_75t_R FILLER_207_600 ();
 DECAPx4_ASAP7_75t_R FILLER_207_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_625 ();
 DECAPx10_ASAP7_75t_R FILLER_207_632 ();
 DECAPx4_ASAP7_75t_R FILLER_207_654 ();
 FILLER_ASAP7_75t_R FILLER_207_664 ();
 FILLER_ASAP7_75t_R FILLER_207_672 ();
 DECAPx1_ASAP7_75t_R FILLER_207_686 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_694 ();
 FILLER_ASAP7_75t_R FILLER_207_707 ();
 DECAPx6_ASAP7_75t_R FILLER_207_727 ();
 FILLER_ASAP7_75t_R FILLER_207_741 ();
 DECAPx2_ASAP7_75t_R FILLER_207_765 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_771 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_207_818 ();
 DECAPx2_ASAP7_75t_R FILLER_207_837 ();
 FILLER_ASAP7_75t_R FILLER_207_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_871 ();
 DECAPx1_ASAP7_75t_R FILLER_207_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_912 ();
 FILLER_ASAP7_75t_R FILLER_207_923 ();
 DECAPx2_ASAP7_75t_R FILLER_207_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_207_933 ();
 DECAPx10_ASAP7_75t_R FILLER_208_12 ();
 DECAPx10_ASAP7_75t_R FILLER_208_34 ();
 DECAPx10_ASAP7_75t_R FILLER_208_56 ();
 FILLER_ASAP7_75t_R FILLER_208_78 ();
 DECAPx1_ASAP7_75t_R FILLER_208_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_128 ();
 DECAPx4_ASAP7_75t_R FILLER_208_157 ();
 FILLER_ASAP7_75t_R FILLER_208_167 ();
 DECAPx10_ASAP7_75t_R FILLER_208_195 ();
 DECAPx2_ASAP7_75t_R FILLER_208_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_223 ();
 DECAPx1_ASAP7_75t_R FILLER_208_232 ();
 DECAPx1_ASAP7_75t_R FILLER_208_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_243 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_266 ();
 FILLER_ASAP7_75t_R FILLER_208_274 ();
 DECAPx10_ASAP7_75t_R FILLER_208_288 ();
 DECAPx10_ASAP7_75t_R FILLER_208_310 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_332 ();
 DECAPx10_ASAP7_75t_R FILLER_208_341 ();
 DECAPx10_ASAP7_75t_R FILLER_208_389 ();
 DECAPx6_ASAP7_75t_R FILLER_208_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_425 ();
 DECAPx6_ASAP7_75t_R FILLER_208_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_443 ();
 DECAPx2_ASAP7_75t_R FILLER_208_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_459 ();
 DECAPx1_ASAP7_75t_R FILLER_208_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_487 ();
 DECAPx6_ASAP7_75t_R FILLER_208_500 ();
 DECAPx2_ASAP7_75t_R FILLER_208_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_520 ();
 FILLER_ASAP7_75t_R FILLER_208_586 ();
 DECAPx10_ASAP7_75t_R FILLER_208_596 ();
 DECAPx10_ASAP7_75t_R FILLER_208_618 ();
 DECAPx1_ASAP7_75t_R FILLER_208_640 ();
 FILLER_ASAP7_75t_R FILLER_208_654 ();
 DECAPx1_ASAP7_75t_R FILLER_208_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_678 ();
 DECAPx10_ASAP7_75t_R FILLER_208_689 ();
 DECAPx10_ASAP7_75t_R FILLER_208_711 ();
 DECAPx6_ASAP7_75t_R FILLER_208_733 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_747 ();
 DECAPx6_ASAP7_75t_R FILLER_208_761 ();
 DECAPx2_ASAP7_75t_R FILLER_208_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_781 ();
 DECAPx2_ASAP7_75t_R FILLER_208_788 ();
 FILLER_ASAP7_75t_R FILLER_208_794 ();
 DECAPx6_ASAP7_75t_R FILLER_208_812 ();
 DECAPx2_ASAP7_75t_R FILLER_208_826 ();
 DECAPx2_ASAP7_75t_R FILLER_208_847 ();
 DECAPx4_ASAP7_75t_R FILLER_208_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_208_884 ();
 DECAPx6_ASAP7_75t_R FILLER_208_894 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_208_931 ();
 DECAPx10_ASAP7_75t_R FILLER_209_7 ();
 DECAPx10_ASAP7_75t_R FILLER_209_29 ();
 DECAPx10_ASAP7_75t_R FILLER_209_51 ();
 DECAPx6_ASAP7_75t_R FILLER_209_73 ();
 DECAPx1_ASAP7_75t_R FILLER_209_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_91 ();
 DECAPx4_ASAP7_75t_R FILLER_209_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_145 ();
 DECAPx10_ASAP7_75t_R FILLER_209_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_183 ();
 DECAPx2_ASAP7_75t_R FILLER_209_187 ();
 FILLER_ASAP7_75t_R FILLER_209_193 ();
 DECAPx10_ASAP7_75t_R FILLER_209_201 ();
 DECAPx4_ASAP7_75t_R FILLER_209_223 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_233 ();
 DECAPx2_ASAP7_75t_R FILLER_209_242 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_248 ();
 DECAPx10_ASAP7_75t_R FILLER_209_255 ();
 DECAPx10_ASAP7_75t_R FILLER_209_277 ();
 DECAPx6_ASAP7_75t_R FILLER_209_299 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_313 ();
 DECAPx1_ASAP7_75t_R FILLER_209_319 ();
 DECAPx4_ASAP7_75t_R FILLER_209_355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_384 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_393 ();
 FILLER_ASAP7_75t_R FILLER_209_420 ();
 DECAPx2_ASAP7_75t_R FILLER_209_432 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_450 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_459 ();
 DECAPx1_ASAP7_75t_R FILLER_209_492 ();
 DECAPx6_ASAP7_75t_R FILLER_209_503 ();
 DECAPx2_ASAP7_75t_R FILLER_209_517 ();
 DECAPx6_ASAP7_75t_R FILLER_209_529 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_543 ();
 FILLER_ASAP7_75t_R FILLER_209_557 ();
 DECAPx2_ASAP7_75t_R FILLER_209_574 ();
 DECAPx10_ASAP7_75t_R FILLER_209_603 ();
 DECAPx1_ASAP7_75t_R FILLER_209_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_629 ();
 DECAPx1_ASAP7_75t_R FILLER_209_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_661 ();
 DECAPx4_ASAP7_75t_R FILLER_209_680 ();
 DECAPx1_ASAP7_75t_R FILLER_209_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_700 ();
 DECAPx10_ASAP7_75t_R FILLER_209_707 ();
 DECAPx6_ASAP7_75t_R FILLER_209_729 ();
 DECAPx2_ASAP7_75t_R FILLER_209_743 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_749 ();
 DECAPx10_ASAP7_75t_R FILLER_209_766 ();
 DECAPx10_ASAP7_75t_R FILLER_209_788 ();
 DECAPx4_ASAP7_75t_R FILLER_209_810 ();
 FILLER_ASAP7_75t_R FILLER_209_820 ();
 DECAPx2_ASAP7_75t_R FILLER_209_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_836 ();
 DECAPx6_ASAP7_75t_R FILLER_209_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_862 ();
 DECAPx10_ASAP7_75t_R FILLER_209_877 ();
 DECAPx2_ASAP7_75t_R FILLER_209_899 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_209_905 ();
 DECAPx2_ASAP7_75t_R FILLER_209_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_209_924 ();
 FILLER_ASAP7_75t_R FILLER_209_932 ();
 DECAPx10_ASAP7_75t_R FILLER_210_2 ();
 DECAPx10_ASAP7_75t_R FILLER_210_24 ();
 DECAPx10_ASAP7_75t_R FILLER_210_46 ();
 DECAPx6_ASAP7_75t_R FILLER_210_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_82 ();
 DECAPx2_ASAP7_75t_R FILLER_210_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_101 ();
 DECAPx1_ASAP7_75t_R FILLER_210_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_116 ();
 FILLER_ASAP7_75t_R FILLER_210_125 ();
 DECAPx2_ASAP7_75t_R FILLER_210_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_162 ();
 DECAPx1_ASAP7_75t_R FILLER_210_169 ();
 DECAPx4_ASAP7_75t_R FILLER_210_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_193 ();
 DECAPx2_ASAP7_75t_R FILLER_210_209 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_215 ();
 FILLER_ASAP7_75t_R FILLER_210_224 ();
 DECAPx2_ASAP7_75t_R FILLER_210_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_263 ();
 DECAPx6_ASAP7_75t_R FILLER_210_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_286 ();
 DECAPx2_ASAP7_75t_R FILLER_210_293 ();
 FILLER_ASAP7_75t_R FILLER_210_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_326 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_461 ();
 DECAPx2_ASAP7_75t_R FILLER_210_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_470 ();
 DECAPx10_ASAP7_75t_R FILLER_210_479 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_501 ();
 DECAPx6_ASAP7_75t_R FILLER_210_510 ();
 DECAPx1_ASAP7_75t_R FILLER_210_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_528 ();
 DECAPx10_ASAP7_75t_R FILLER_210_537 ();
 DECAPx1_ASAP7_75t_R FILLER_210_559 ();
 FILLER_ASAP7_75t_R FILLER_210_571 ();
 DECAPx10_ASAP7_75t_R FILLER_210_580 ();
 DECAPx1_ASAP7_75t_R FILLER_210_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_606 ();
 DECAPx2_ASAP7_75t_R FILLER_210_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_640 ();
 DECAPx2_ASAP7_75t_R FILLER_210_655 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_661 ();
 DECAPx6_ASAP7_75t_R FILLER_210_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_684 ();
 FILLER_ASAP7_75t_R FILLER_210_701 ();
 DECAPx1_ASAP7_75t_R FILLER_210_711 ();
 FILLER_ASAP7_75t_R FILLER_210_722 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_210_740 ();
 DECAPx1_ASAP7_75t_R FILLER_210_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_772 ();
 DECAPx6_ASAP7_75t_R FILLER_210_783 ();
 DECAPx4_ASAP7_75t_R FILLER_210_802 ();
 FILLER_ASAP7_75t_R FILLER_210_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_840 ();
 DECAPx4_ASAP7_75t_R FILLER_210_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_210_876 ();
 DECAPx6_ASAP7_75t_R FILLER_210_883 ();
 FILLER_ASAP7_75t_R FILLER_210_897 ();
 DECAPx1_ASAP7_75t_R FILLER_210_911 ();
 DECAPx1_ASAP7_75t_R FILLER_210_920 ();
 DECAPx10_ASAP7_75t_R FILLER_211_2 ();
 DECAPx10_ASAP7_75t_R FILLER_211_24 ();
 DECAPx10_ASAP7_75t_R FILLER_211_46 ();
 DECAPx6_ASAP7_75t_R FILLER_211_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_82 ();
 DECAPx2_ASAP7_75t_R FILLER_211_91 ();
 FILLER_ASAP7_75t_R FILLER_211_97 ();
 DECAPx6_ASAP7_75t_R FILLER_211_111 ();
 FILLER_ASAP7_75t_R FILLER_211_125 ();
 DECAPx4_ASAP7_75t_R FILLER_211_133 ();
 FILLER_ASAP7_75t_R FILLER_211_143 ();
 DECAPx2_ASAP7_75t_R FILLER_211_151 ();
 FILLER_ASAP7_75t_R FILLER_211_157 ();
 DECAPx6_ASAP7_75t_R FILLER_211_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_207 ();
 DECAPx4_ASAP7_75t_R FILLER_211_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_224 ();
 DECAPx4_ASAP7_75t_R FILLER_211_253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_263 ();
 DECAPx1_ASAP7_75t_R FILLER_211_306 ();
 DECAPx1_ASAP7_75t_R FILLER_211_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_362 ();
 DECAPx2_ASAP7_75t_R FILLER_211_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_375 ();
 DECAPx6_ASAP7_75t_R FILLER_211_386 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_400 ();
 DECAPx1_ASAP7_75t_R FILLER_211_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_435 ();
 DECAPx2_ASAP7_75t_R FILLER_211_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_460 ();
 DECAPx10_ASAP7_75t_R FILLER_211_467 ();
 DECAPx4_ASAP7_75t_R FILLER_211_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_499 ();
 FILLER_ASAP7_75t_R FILLER_211_503 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_513 ();
 DECAPx1_ASAP7_75t_R FILLER_211_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_527 ();
 DECAPx10_ASAP7_75t_R FILLER_211_540 ();
 DECAPx4_ASAP7_75t_R FILLER_211_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_572 ();
 DECAPx6_ASAP7_75t_R FILLER_211_581 ();
 DECAPx2_ASAP7_75t_R FILLER_211_606 ();
 FILLER_ASAP7_75t_R FILLER_211_612 ();
 DECAPx10_ASAP7_75t_R FILLER_211_626 ();
 DECAPx10_ASAP7_75t_R FILLER_211_648 ();
 DECAPx6_ASAP7_75t_R FILLER_211_670 ();
 FILLER_ASAP7_75t_R FILLER_211_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_692 ();
 DECAPx4_ASAP7_75t_R FILLER_211_699 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_211_716 ();
 DECAPx1_ASAP7_75t_R FILLER_211_727 ();
 DECAPx1_ASAP7_75t_R FILLER_211_741 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_745 ();
 DECAPx1_ASAP7_75t_R FILLER_211_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_766 ();
 FILLER_ASAP7_75t_R FILLER_211_793 ();
 DECAPx2_ASAP7_75t_R FILLER_211_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_827 ();
 DECAPx2_ASAP7_75t_R FILLER_211_854 ();
 DECAPx1_ASAP7_75t_R FILLER_211_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_211_933 ();
 DECAPx10_ASAP7_75t_R FILLER_212_2 ();
 DECAPx10_ASAP7_75t_R FILLER_212_24 ();
 DECAPx10_ASAP7_75t_R FILLER_212_46 ();
 DECAPx2_ASAP7_75t_R FILLER_212_68 ();
 FILLER_ASAP7_75t_R FILLER_212_100 ();
 DECAPx10_ASAP7_75t_R FILLER_212_110 ();
 DECAPx4_ASAP7_75t_R FILLER_212_132 ();
 FILLER_ASAP7_75t_R FILLER_212_142 ();
 DECAPx1_ASAP7_75t_R FILLER_212_156 ();
 DECAPx6_ASAP7_75t_R FILLER_212_166 ();
 DECAPx2_ASAP7_75t_R FILLER_212_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_186 ();
 DECAPx2_ASAP7_75t_R FILLER_212_199 ();
 FILLER_ASAP7_75t_R FILLER_212_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_215 ();
 DECAPx1_ASAP7_75t_R FILLER_212_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_240 ();
 DECAPx2_ASAP7_75t_R FILLER_212_250 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_256 ();
 DECAPx4_ASAP7_75t_R FILLER_212_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_276 ();
 FILLER_ASAP7_75t_R FILLER_212_291 ();
 DECAPx2_ASAP7_75t_R FILLER_212_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_306 ();
 FILLER_ASAP7_75t_R FILLER_212_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_390 ();
 DECAPx10_ASAP7_75t_R FILLER_212_413 ();
 DECAPx10_ASAP7_75t_R FILLER_212_435 ();
 DECAPx1_ASAP7_75t_R FILLER_212_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_461 ();
 DECAPx4_ASAP7_75t_R FILLER_212_464 ();
 FILLER_ASAP7_75t_R FILLER_212_488 ();
 DECAPx6_ASAP7_75t_R FILLER_212_496 ();
 FILLER_ASAP7_75t_R FILLER_212_510 ();
 DECAPx2_ASAP7_75t_R FILLER_212_526 ();
 DECAPx1_ASAP7_75t_R FILLER_212_538 ();
 DECAPx10_ASAP7_75t_R FILLER_212_556 ();
 DECAPx6_ASAP7_75t_R FILLER_212_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_592 ();
 DECAPx2_ASAP7_75t_R FILLER_212_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_632 ();
 DECAPx10_ASAP7_75t_R FILLER_212_639 ();
 DECAPx6_ASAP7_75t_R FILLER_212_661 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_675 ();
 DECAPx10_ASAP7_75t_R FILLER_212_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_212_705 ();
 FILLER_ASAP7_75t_R FILLER_212_714 ();
 DECAPx2_ASAP7_75t_R FILLER_212_722 ();
 FILLER_ASAP7_75t_R FILLER_212_728 ();
 DECAPx6_ASAP7_75t_R FILLER_212_749 ();
 DECAPx1_ASAP7_75t_R FILLER_212_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_767 ();
 FILLER_ASAP7_75t_R FILLER_212_781 ();
 DECAPx6_ASAP7_75t_R FILLER_212_825 ();
 DECAPx1_ASAP7_75t_R FILLER_212_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_843 ();
 DECAPx6_ASAP7_75t_R FILLER_212_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_212_918 ();
 DECAPx10_ASAP7_75t_R FILLER_213_7 ();
 DECAPx10_ASAP7_75t_R FILLER_213_29 ();
 DECAPx10_ASAP7_75t_R FILLER_213_51 ();
 DECAPx2_ASAP7_75t_R FILLER_213_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_79 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_86 ();
 DECAPx4_ASAP7_75t_R FILLER_213_92 ();
 DECAPx6_ASAP7_75t_R FILLER_213_136 ();
 DECAPx2_ASAP7_75t_R FILLER_213_150 ();
 DECAPx6_ASAP7_75t_R FILLER_213_182 ();
 DECAPx1_ASAP7_75t_R FILLER_213_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_206 ();
 DECAPx2_ASAP7_75t_R FILLER_213_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_219 ();
 FILLER_ASAP7_75t_R FILLER_213_256 ();
 DECAPx4_ASAP7_75t_R FILLER_213_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_275 ();
 DECAPx2_ASAP7_75t_R FILLER_213_282 ();
 FILLER_ASAP7_75t_R FILLER_213_288 ();
 DECAPx10_ASAP7_75t_R FILLER_213_295 ();
 DECAPx6_ASAP7_75t_R FILLER_213_317 ();
 DECAPx2_ASAP7_75t_R FILLER_213_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_350 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_354 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_370 ();
 FILLER_ASAP7_75t_R FILLER_213_383 ();
 DECAPx1_ASAP7_75t_R FILLER_213_420 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_443 ();
 DECAPx1_ASAP7_75t_R FILLER_213_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_456 ();
 FILLER_ASAP7_75t_R FILLER_213_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_502 ();
 DECAPx2_ASAP7_75t_R FILLER_213_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_532 ();
 DECAPx6_ASAP7_75t_R FILLER_213_559 ();
 FILLER_ASAP7_75t_R FILLER_213_573 ();
 FILLER_ASAP7_75t_R FILLER_213_582 ();
 DECAPx1_ASAP7_75t_R FILLER_213_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_595 ();
 DECAPx6_ASAP7_75t_R FILLER_213_612 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_641 ();
 DECAPx2_ASAP7_75t_R FILLER_213_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_663 ();
 DECAPx4_ASAP7_75t_R FILLER_213_680 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_690 ();
 DECAPx2_ASAP7_75t_R FILLER_213_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_714 ();
 DECAPx10_ASAP7_75t_R FILLER_213_723 ();
 DECAPx2_ASAP7_75t_R FILLER_213_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_751 ();
 DECAPx4_ASAP7_75t_R FILLER_213_768 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_213_778 ();
 DECAPx1_ASAP7_75t_R FILLER_213_784 ();
 DECAPx2_ASAP7_75t_R FILLER_213_804 ();
 FILLER_ASAP7_75t_R FILLER_213_810 ();
 FILLER_ASAP7_75t_R FILLER_213_819 ();
 DECAPx10_ASAP7_75t_R FILLER_213_824 ();
 DECAPx1_ASAP7_75t_R FILLER_213_846 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_850 ();
 DECAPx6_ASAP7_75t_R FILLER_213_870 ();
 DECAPx2_ASAP7_75t_R FILLER_213_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_213_933 ();
 DECAPx10_ASAP7_75t_R FILLER_214_12 ();
 DECAPx10_ASAP7_75t_R FILLER_214_34 ();
 DECAPx10_ASAP7_75t_R FILLER_214_56 ();
 DECAPx10_ASAP7_75t_R FILLER_214_84 ();
 DECAPx2_ASAP7_75t_R FILLER_214_106 ();
 DECAPx4_ASAP7_75t_R FILLER_214_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_160 ();
 DECAPx2_ASAP7_75t_R FILLER_214_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_173 ();
 DECAPx1_ASAP7_75t_R FILLER_214_190 ();
 DECAPx1_ASAP7_75t_R FILLER_214_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_224 ();
 DECAPx6_ASAP7_75t_R FILLER_214_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_244 ();
 FILLER_ASAP7_75t_R FILLER_214_248 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_278 ();
 DECAPx10_ASAP7_75t_R FILLER_214_291 ();
 DECAPx10_ASAP7_75t_R FILLER_214_313 ();
 DECAPx10_ASAP7_75t_R FILLER_214_335 ();
 FILLER_ASAP7_75t_R FILLER_214_357 ();
 DECAPx2_ASAP7_75t_R FILLER_214_365 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_384 ();
 FILLER_ASAP7_75t_R FILLER_214_388 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_402 ();
 DECAPx4_ASAP7_75t_R FILLER_214_408 ();
 FILLER_ASAP7_75t_R FILLER_214_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_471 ();
 FILLER_ASAP7_75t_R FILLER_214_494 ();
 DECAPx1_ASAP7_75t_R FILLER_214_505 ();
 DECAPx10_ASAP7_75t_R FILLER_214_514 ();
 DECAPx2_ASAP7_75t_R FILLER_214_536 ();
 FILLER_ASAP7_75t_R FILLER_214_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_552 ();
 DECAPx6_ASAP7_75t_R FILLER_214_599 ();
 DECAPx2_ASAP7_75t_R FILLER_214_613 ();
 DECAPx1_ASAP7_75t_R FILLER_214_684 ();
 FILLERxp5_ASAP7_75t_R FILLER_214_688 ();
 DECAPx4_ASAP7_75t_R FILLER_214_709 ();
 FILLER_ASAP7_75t_R FILLER_214_719 ();
 DECAPx6_ASAP7_75t_R FILLER_214_728 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_742 ();
 DECAPx10_ASAP7_75t_R FILLER_214_751 ();
 DECAPx10_ASAP7_75t_R FILLER_214_781 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_803 ();
 DECAPx4_ASAP7_75t_R FILLER_214_832 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_842 ();
 DECAPx10_ASAP7_75t_R FILLER_214_871 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_214_893 ();
 FILLER_ASAP7_75t_R FILLER_214_932 ();
 DECAPx10_ASAP7_75t_R FILLER_215_12 ();
 DECAPx10_ASAP7_75t_R FILLER_215_34 ();
 DECAPx6_ASAP7_75t_R FILLER_215_56 ();
 DECAPx10_ASAP7_75t_R FILLER_215_96 ();
 DECAPx1_ASAP7_75t_R FILLER_215_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_122 ();
 FILLER_ASAP7_75t_R FILLER_215_132 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_143 ();
 DECAPx6_ASAP7_75t_R FILLER_215_152 ();
 FILLER_ASAP7_75t_R FILLER_215_166 ();
 DECAPx6_ASAP7_75t_R FILLER_215_174 ();
 DECAPx2_ASAP7_75t_R FILLER_215_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_194 ();
 DECAPx2_ASAP7_75t_R FILLER_215_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_207 ();
 DECAPx10_ASAP7_75t_R FILLER_215_211 ();
 DECAPx10_ASAP7_75t_R FILLER_215_233 ();
 DECAPx1_ASAP7_75t_R FILLER_215_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_294 ();
 DECAPx2_ASAP7_75t_R FILLER_215_305 ();
 FILLER_ASAP7_75t_R FILLER_215_311 ();
 FILLER_ASAP7_75t_R FILLER_215_319 ();
 DECAPx2_ASAP7_75t_R FILLER_215_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_341 ();
 DECAPx10_ASAP7_75t_R FILLER_215_348 ();
 DECAPx1_ASAP7_75t_R FILLER_215_370 ();
 DECAPx1_ASAP7_75t_R FILLER_215_383 ();
 DECAPx1_ASAP7_75t_R FILLER_215_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_412 ();
 DECAPx1_ASAP7_75t_R FILLER_215_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_456 ();
 DECAPx10_ASAP7_75t_R FILLER_215_483 ();
 DECAPx1_ASAP7_75t_R FILLER_215_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_509 ();
 DECAPx1_ASAP7_75t_R FILLER_215_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_521 ();
 DECAPx6_ASAP7_75t_R FILLER_215_529 ();
 DECAPx1_ASAP7_75t_R FILLER_215_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_547 ();
 DECAPx2_ASAP7_75t_R FILLER_215_551 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_557 ();
 FILLER_ASAP7_75t_R FILLER_215_564 ();
 DECAPx10_ASAP7_75t_R FILLER_215_587 ();
 DECAPx6_ASAP7_75t_R FILLER_215_609 ();
 DECAPx1_ASAP7_75t_R FILLER_215_623 ();
 DECAPx2_ASAP7_75t_R FILLER_215_633 ();
 FILLER_ASAP7_75t_R FILLER_215_639 ();
 DECAPx2_ASAP7_75t_R FILLER_215_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_680 ();
 DECAPx2_ASAP7_75t_R FILLER_215_719 ();
 FILLER_ASAP7_75t_R FILLER_215_725 ();
 DECAPx2_ASAP7_75t_R FILLER_215_732 ();
 DECAPx1_ASAP7_75t_R FILLER_215_744 ();
 DECAPx1_ASAP7_75t_R FILLER_215_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_759 ();
 DECAPx1_ASAP7_75t_R FILLER_215_769 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_773 ();
 DECAPx1_ASAP7_75t_R FILLER_215_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_788 ();
 DECAPx6_ASAP7_75t_R FILLER_215_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_813 ();
 DECAPx1_ASAP7_75t_R FILLER_215_822 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_841 ();
 DECAPx2_ASAP7_75t_R FILLER_215_848 ();
 DECAPx2_ASAP7_75t_R FILLER_215_869 ();
 FILLER_ASAP7_75t_R FILLER_215_875 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_215_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_215_927 ();
 DECAPx10_ASAP7_75t_R FILLER_216_2 ();
 DECAPx10_ASAP7_75t_R FILLER_216_24 ();
 DECAPx10_ASAP7_75t_R FILLER_216_46 ();
 DECAPx4_ASAP7_75t_R FILLER_216_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_78 ();
 FILLER_ASAP7_75t_R FILLER_216_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_109 ();
 DECAPx10_ASAP7_75t_R FILLER_216_122 ();
 DECAPx2_ASAP7_75t_R FILLER_216_144 ();
 DECAPx10_ASAP7_75t_R FILLER_216_158 ();
 DECAPx10_ASAP7_75t_R FILLER_216_180 ();
 DECAPx1_ASAP7_75t_R FILLER_216_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_206 ();
 DECAPx1_ASAP7_75t_R FILLER_216_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_221 ();
 DECAPx6_ASAP7_75t_R FILLER_216_225 ();
 DECAPx1_ASAP7_75t_R FILLER_216_239 ();
 DECAPx6_ASAP7_75t_R FILLER_216_246 ();
 DECAPx1_ASAP7_75t_R FILLER_216_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_264 ();
 DECAPx2_ASAP7_75t_R FILLER_216_281 ();
 FILLER_ASAP7_75t_R FILLER_216_287 ();
 DECAPx4_ASAP7_75t_R FILLER_216_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_369 ();
 DECAPx1_ASAP7_75t_R FILLER_216_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_396 ();
 DECAPx1_ASAP7_75t_R FILLER_216_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_417 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_431 ();
 DECAPx2_ASAP7_75t_R FILLER_216_440 ();
 FILLER_ASAP7_75t_R FILLER_216_446 ();
 DECAPx2_ASAP7_75t_R FILLER_216_454 ();
 FILLER_ASAP7_75t_R FILLER_216_460 ();
 DECAPx2_ASAP7_75t_R FILLER_216_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_470 ();
 DECAPx10_ASAP7_75t_R FILLER_216_474 ();
 DECAPx10_ASAP7_75t_R FILLER_216_496 ();
 FILLER_ASAP7_75t_R FILLER_216_518 ();
 DECAPx1_ASAP7_75t_R FILLER_216_534 ();
 DECAPx2_ASAP7_75t_R FILLER_216_541 ();
 FILLER_ASAP7_75t_R FILLER_216_547 ();
 FILLER_ASAP7_75t_R FILLER_216_559 ();
 DECAPx10_ASAP7_75t_R FILLER_216_569 ();
 DECAPx4_ASAP7_75t_R FILLER_216_591 ();
 FILLER_ASAP7_75t_R FILLER_216_615 ();
 DECAPx10_ASAP7_75t_R FILLER_216_626 ();
 DECAPx10_ASAP7_75t_R FILLER_216_648 ();
 DECAPx2_ASAP7_75t_R FILLER_216_670 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_676 ();
 DECAPx6_ASAP7_75t_R FILLER_216_685 ();
 DECAPx4_ASAP7_75t_R FILLER_216_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_713 ();
 DECAPx1_ASAP7_75t_R FILLER_216_745 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_756 ();
 DECAPx4_ASAP7_75t_R FILLER_216_790 ();
 FILLER_ASAP7_75t_R FILLER_216_800 ();
 DECAPx6_ASAP7_75t_R FILLER_216_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_821 ();
 DECAPx6_ASAP7_75t_R FILLER_216_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_216_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_906 ();
 FILLERxp5_ASAP7_75t_R FILLER_216_920 ();
 DECAPx10_ASAP7_75t_R FILLER_217_2 ();
 DECAPx10_ASAP7_75t_R FILLER_217_24 ();
 DECAPx10_ASAP7_75t_R FILLER_217_46 ();
 DECAPx6_ASAP7_75t_R FILLER_217_68 ();
 DECAPx1_ASAP7_75t_R FILLER_217_82 ();
 DECAPx1_ASAP7_75t_R FILLER_217_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_132 ();
 FILLER_ASAP7_75t_R FILLER_217_139 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_152 ();
 DECAPx4_ASAP7_75t_R FILLER_217_161 ();
 DECAPx4_ASAP7_75t_R FILLER_217_179 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_195 ();
 FILLER_ASAP7_75t_R FILLER_217_230 ();
 DECAPx10_ASAP7_75t_R FILLER_217_258 ();
 DECAPx6_ASAP7_75t_R FILLER_217_280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_294 ();
 DECAPx1_ASAP7_75t_R FILLER_217_300 ();
 DECAPx1_ASAP7_75t_R FILLER_217_312 ();
 FILLER_ASAP7_75t_R FILLER_217_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_361 ();
 DECAPx1_ASAP7_75t_R FILLER_217_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_375 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_382 ();
 DECAPx10_ASAP7_75t_R FILLER_217_391 ();
 DECAPx10_ASAP7_75t_R FILLER_217_413 ();
 FILLER_ASAP7_75t_R FILLER_217_435 ();
 DECAPx2_ASAP7_75t_R FILLER_217_463 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_469 ();
 DECAPx1_ASAP7_75t_R FILLER_217_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_522 ();
 DECAPx10_ASAP7_75t_R FILLER_217_549 ();
 DECAPx6_ASAP7_75t_R FILLER_217_571 ();
 DECAPx2_ASAP7_75t_R FILLER_217_585 ();
 DECAPx1_ASAP7_75t_R FILLER_217_599 ();
 DECAPx10_ASAP7_75t_R FILLER_217_610 ();
 DECAPx10_ASAP7_75t_R FILLER_217_632 ();
 DECAPx2_ASAP7_75t_R FILLER_217_654 ();
 DECAPx10_ASAP7_75t_R FILLER_217_672 ();
 DECAPx4_ASAP7_75t_R FILLER_217_694 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_704 ();
 DECAPx1_ASAP7_75t_R FILLER_217_728 ();
 DECAPx2_ASAP7_75t_R FILLER_217_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_217_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_217_804 ();
 DECAPx4_ASAP7_75t_R FILLER_217_811 ();
 DECAPx2_ASAP7_75t_R FILLER_217_824 ();
 FILLER_ASAP7_75t_R FILLER_217_830 ();
 DECAPx6_ASAP7_75t_R FILLER_217_850 ();
 DECAPx1_ASAP7_75t_R FILLER_217_864 ();
 DECAPx1_ASAP7_75t_R FILLER_217_886 ();
 FILLER_ASAP7_75t_R FILLER_217_927 ();
 DECAPx10_ASAP7_75t_R FILLER_218_7 ();
 DECAPx10_ASAP7_75t_R FILLER_218_29 ();
 DECAPx10_ASAP7_75t_R FILLER_218_51 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_100 ();
 FILLER_ASAP7_75t_R FILLER_218_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_164 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_179 ();
 DECAPx2_ASAP7_75t_R FILLER_218_208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_214 ();
 FILLER_ASAP7_75t_R FILLER_218_243 ();
 DECAPx4_ASAP7_75t_R FILLER_218_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_275 ();
 DECAPx2_ASAP7_75t_R FILLER_218_288 ();
 DECAPx10_ASAP7_75t_R FILLER_218_301 ();
 DECAPx10_ASAP7_75t_R FILLER_218_323 ();
 FILLER_ASAP7_75t_R FILLER_218_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_352 ();
 DECAPx2_ASAP7_75t_R FILLER_218_359 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_365 ();
 DECAPx4_ASAP7_75t_R FILLER_218_374 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_384 ();
 DECAPx10_ASAP7_75t_R FILLER_218_399 ();
 DECAPx10_ASAP7_75t_R FILLER_218_421 ();
 DECAPx2_ASAP7_75t_R FILLER_218_443 ();
 FILLER_ASAP7_75t_R FILLER_218_449 ();
 DECAPx2_ASAP7_75t_R FILLER_218_454 ();
 FILLER_ASAP7_75t_R FILLER_218_460 ();
 DECAPx2_ASAP7_75t_R FILLER_218_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_470 ();
 DECAPx1_ASAP7_75t_R FILLER_218_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_487 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_504 ();
 DECAPx6_ASAP7_75t_R FILLER_218_510 ();
 DECAPx2_ASAP7_75t_R FILLER_218_524 ();
 DECAPx10_ASAP7_75t_R FILLER_218_538 ();
 DECAPx10_ASAP7_75t_R FILLER_218_560 ();
 FILLER_ASAP7_75t_R FILLER_218_582 ();
 FILLER_ASAP7_75t_R FILLER_218_590 ();
 FILLER_ASAP7_75t_R FILLER_218_601 ();
 DECAPx6_ASAP7_75t_R FILLER_218_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_631 ();
 DECAPx6_ASAP7_75t_R FILLER_218_643 ();
 DECAPx1_ASAP7_75t_R FILLER_218_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_661 ();
 DECAPx10_ASAP7_75t_R FILLER_218_669 ();
 DECAPx1_ASAP7_75t_R FILLER_218_691 ();
 DECAPx2_ASAP7_75t_R FILLER_218_707 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_719 ();
 FILLER_ASAP7_75t_R FILLER_218_728 ();
 DECAPx4_ASAP7_75t_R FILLER_218_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_748 ();
 FILLER_ASAP7_75t_R FILLER_218_761 ();
 DECAPx1_ASAP7_75t_R FILLER_218_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_777 ();
 DECAPx1_ASAP7_75t_R FILLER_218_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_792 ();
 DECAPx4_ASAP7_75t_R FILLER_218_836 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_218_846 ();
 DECAPx2_ASAP7_75t_R FILLER_218_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_860 ();
 DECAPx1_ASAP7_75t_R FILLER_218_875 ();
 FILLER_ASAP7_75t_R FILLER_218_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_218_933 ();
 DECAPx10_ASAP7_75t_R FILLER_219_7 ();
 DECAPx10_ASAP7_75t_R FILLER_219_29 ();
 DECAPx10_ASAP7_75t_R FILLER_219_51 ();
 DECAPx2_ASAP7_75t_R FILLER_219_73 ();
 FILLER_ASAP7_75t_R FILLER_219_79 ();
 FILLER_ASAP7_75t_R FILLER_219_87 ();
 DECAPx10_ASAP7_75t_R FILLER_219_92 ();
 DECAPx2_ASAP7_75t_R FILLER_219_114 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_126 ();
 DECAPx2_ASAP7_75t_R FILLER_219_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_146 ();
 DECAPx2_ASAP7_75t_R FILLER_219_150 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_156 ();
 DECAPx1_ASAP7_75t_R FILLER_219_171 ();
 DECAPx2_ASAP7_75t_R FILLER_219_190 ();
 DECAPx6_ASAP7_75t_R FILLER_219_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_248 ();
 DECAPx1_ASAP7_75t_R FILLER_219_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_261 ();
 FILLER_ASAP7_75t_R FILLER_219_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_307 ();
 DECAPx10_ASAP7_75t_R FILLER_219_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_336 ();
 DECAPx2_ASAP7_75t_R FILLER_219_343 ();
 FILLER_ASAP7_75t_R FILLER_219_356 ();
 FILLER_ASAP7_75t_R FILLER_219_413 ();
 DECAPx6_ASAP7_75t_R FILLER_219_420 ();
 FILLER_ASAP7_75t_R FILLER_219_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_441 ();
 FILLER_ASAP7_75t_R FILLER_219_474 ();
 FILLER_ASAP7_75t_R FILLER_219_502 ();
 DECAPx6_ASAP7_75t_R FILLER_219_524 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_538 ();
 FILLER_ASAP7_75t_R FILLER_219_553 ();
 FILLER_ASAP7_75t_R FILLER_219_575 ();
 DECAPx2_ASAP7_75t_R FILLER_219_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_627 ();
 DECAPx1_ASAP7_75t_R FILLER_219_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_646 ();
 DECAPx4_ASAP7_75t_R FILLER_219_657 ();
 FILLER_ASAP7_75t_R FILLER_219_667 ();
 DECAPx2_ASAP7_75t_R FILLER_219_675 ();
 DECAPx6_ASAP7_75t_R FILLER_219_708 ();
 FILLER_ASAP7_75t_R FILLER_219_722 ();
 DECAPx4_ASAP7_75t_R FILLER_219_730 ();
 DECAPx10_ASAP7_75t_R FILLER_219_745 ();
 DECAPx10_ASAP7_75t_R FILLER_219_767 ();
 DECAPx2_ASAP7_75t_R FILLER_219_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_795 ();
 DECAPx1_ASAP7_75t_R FILLER_219_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_817 ();
 DECAPx10_ASAP7_75t_R FILLER_219_821 ();
 DECAPx1_ASAP7_75t_R FILLER_219_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_847 ();
 DECAPx4_ASAP7_75t_R FILLER_219_872 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_882 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_219_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_219_897 ();
 FILLER_ASAP7_75t_R FILLER_219_927 ();
 DECAPx10_ASAP7_75t_R FILLER_220_7 ();
 DECAPx10_ASAP7_75t_R FILLER_220_29 ();
 DECAPx10_ASAP7_75t_R FILLER_220_51 ();
 DECAPx10_ASAP7_75t_R FILLER_220_73 ();
 DECAPx4_ASAP7_75t_R FILLER_220_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_105 ();
 DECAPx6_ASAP7_75t_R FILLER_220_141 ();
 DECAPx1_ASAP7_75t_R FILLER_220_155 ();
 DECAPx4_ASAP7_75t_R FILLER_220_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_245 ();
 DECAPx2_ASAP7_75t_R FILLER_220_249 ();
 FILLER_ASAP7_75t_R FILLER_220_255 ();
 DECAPx1_ASAP7_75t_R FILLER_220_271 ();
 DECAPx1_ASAP7_75t_R FILLER_220_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_291 ();
 DECAPx2_ASAP7_75t_R FILLER_220_318 ();
 FILLER_ASAP7_75t_R FILLER_220_324 ();
 FILLER_ASAP7_75t_R FILLER_220_363 ();
 DECAPx2_ASAP7_75t_R FILLER_220_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_377 ();
 DECAPx6_ASAP7_75t_R FILLER_220_381 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_395 ();
 FILLER_ASAP7_75t_R FILLER_220_401 ();
 DECAPx1_ASAP7_75t_R FILLER_220_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_425 ();
 DECAPx4_ASAP7_75t_R FILLER_220_445 ();
 FILLER_ASAP7_75t_R FILLER_220_455 ();
 FILLER_ASAP7_75t_R FILLER_220_460 ();
 DECAPx6_ASAP7_75t_R FILLER_220_471 ();
 DECAPx2_ASAP7_75t_R FILLER_220_485 ();
 DECAPx2_ASAP7_75t_R FILLER_220_494 ();
 FILLER_ASAP7_75t_R FILLER_220_500 ();
 DECAPx2_ASAP7_75t_R FILLER_220_528 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_534 ();
 FILLER_ASAP7_75t_R FILLER_220_564 ();
 DECAPx4_ASAP7_75t_R FILLER_220_593 ();
 FILLER_ASAP7_75t_R FILLER_220_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_611 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_663 ();
 DECAPx1_ASAP7_75t_R FILLER_220_707 ();
 DECAPx2_ASAP7_75t_R FILLER_220_717 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_723 ();
 DECAPx2_ASAP7_75t_R FILLER_220_732 ();
 FILLER_ASAP7_75t_R FILLER_220_738 ();
 DECAPx10_ASAP7_75t_R FILLER_220_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_220_767 ();
 DECAPx6_ASAP7_75t_R FILLER_220_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_789 ();
 DECAPx6_ASAP7_75t_R FILLER_220_821 ();
 DECAPx10_ASAP7_75t_R FILLER_220_843 ();
 DECAPx2_ASAP7_75t_R FILLER_220_865 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_871 ();
 DECAPx4_ASAP7_75t_R FILLER_220_879 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_889 ();
 DECAPx2_ASAP7_75t_R FILLER_220_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_220_901 ();
 DECAPx10_ASAP7_75t_R FILLER_221_7 ();
 DECAPx10_ASAP7_75t_R FILLER_221_29 ();
 DECAPx10_ASAP7_75t_R FILLER_221_51 ();
 DECAPx10_ASAP7_75t_R FILLER_221_73 ();
 DECAPx1_ASAP7_75t_R FILLER_221_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_99 ();
 DECAPx10_ASAP7_75t_R FILLER_221_135 ();
 DECAPx6_ASAP7_75t_R FILLER_221_157 ();
 FILLER_ASAP7_75t_R FILLER_221_171 ();
 DECAPx4_ASAP7_75t_R FILLER_221_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_224 ();
 DECAPx10_ASAP7_75t_R FILLER_221_244 ();
 DECAPx10_ASAP7_75t_R FILLER_221_266 ();
 DECAPx6_ASAP7_75t_R FILLER_221_288 ();
 DECAPx1_ASAP7_75t_R FILLER_221_302 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_306 ();
 DECAPx1_ASAP7_75t_R FILLER_221_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_339 ();
 DECAPx1_ASAP7_75t_R FILLER_221_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_353 ();
 DECAPx10_ASAP7_75t_R FILLER_221_362 ();
 DECAPx6_ASAP7_75t_R FILLER_221_384 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_398 ();
 DECAPx1_ASAP7_75t_R FILLER_221_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_441 ();
 DECAPx10_ASAP7_75t_R FILLER_221_470 ();
 DECAPx2_ASAP7_75t_R FILLER_221_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_498 ();
 DECAPx2_ASAP7_75t_R FILLER_221_509 ();
 FILLER_ASAP7_75t_R FILLER_221_515 ();
 DECAPx1_ASAP7_75t_R FILLER_221_520 ();
 DECAPx1_ASAP7_75t_R FILLER_221_532 ();
 DECAPx6_ASAP7_75t_R FILLER_221_539 ();
 DECAPx2_ASAP7_75t_R FILLER_221_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_559 ();
 DECAPx1_ASAP7_75t_R FILLER_221_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_572 ();
 DECAPx2_ASAP7_75t_R FILLER_221_581 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_628 ();
 DECAPx6_ASAP7_75t_R FILLER_221_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_646 ();
 DECAPx2_ASAP7_75t_R FILLER_221_664 ();
 FILLER_ASAP7_75t_R FILLER_221_670 ();
 DECAPx1_ASAP7_75t_R FILLER_221_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_691 ();
 DECAPx6_ASAP7_75t_R FILLER_221_710 ();
 DECAPx2_ASAP7_75t_R FILLER_221_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_730 ();
 DECAPx2_ASAP7_75t_R FILLER_221_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_757 ();
 FILLER_ASAP7_75t_R FILLER_221_776 ();
 DECAPx6_ASAP7_75t_R FILLER_221_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_807 ();
 DECAPx4_ASAP7_75t_R FILLER_221_814 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_221_824 ();
 DECAPx1_ASAP7_75t_R FILLER_221_851 ();
 DECAPx2_ASAP7_75t_R FILLER_221_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_867 ();
 DECAPx1_ASAP7_75t_R FILLER_221_874 ();
 DECAPx10_ASAP7_75t_R FILLER_221_883 ();
 DECAPx2_ASAP7_75t_R FILLER_221_905 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_221_919 ();
 DECAPx10_ASAP7_75t_R FILLER_222_7 ();
 DECAPx10_ASAP7_75t_R FILLER_222_29 ();
 DECAPx10_ASAP7_75t_R FILLER_222_51 ();
 DECAPx1_ASAP7_75t_R FILLER_222_73 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_77 ();
 DECAPx2_ASAP7_75t_R FILLER_222_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_99 ();
 DECAPx6_ASAP7_75t_R FILLER_222_130 ();
 FILLER_ASAP7_75t_R FILLER_222_144 ();
 DECAPx10_ASAP7_75t_R FILLER_222_161 ();
 DECAPx2_ASAP7_75t_R FILLER_222_183 ();
 DECAPx6_ASAP7_75t_R FILLER_222_203 ();
 FILLER_ASAP7_75t_R FILLER_222_217 ();
 DECAPx10_ASAP7_75t_R FILLER_222_222 ();
 DECAPx4_ASAP7_75t_R FILLER_222_247 ();
 FILLER_ASAP7_75t_R FILLER_222_263 ();
 DECAPx4_ASAP7_75t_R FILLER_222_271 ();
 FILLER_ASAP7_75t_R FILLER_222_281 ();
 DECAPx2_ASAP7_75t_R FILLER_222_289 ();
 FILLER_ASAP7_75t_R FILLER_222_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_303 ();
 DECAPx1_ASAP7_75t_R FILLER_222_314 ();
 DECAPx6_ASAP7_75t_R FILLER_222_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_338 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_370 ();
 DECAPx4_ASAP7_75t_R FILLER_222_385 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_395 ();
 FILLER_ASAP7_75t_R FILLER_222_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_424 ();
 DECAPx6_ASAP7_75t_R FILLER_222_438 ();
 DECAPx2_ASAP7_75t_R FILLER_222_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_464 ();
 DECAPx2_ASAP7_75t_R FILLER_222_471 ();
 DECAPx10_ASAP7_75t_R FILLER_222_483 ();
 DECAPx2_ASAP7_75t_R FILLER_222_505 ();
 FILLER_ASAP7_75t_R FILLER_222_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_521 ();
 DECAPx10_ASAP7_75t_R FILLER_222_548 ();
 FILLER_ASAP7_75t_R FILLER_222_570 ();
 DECAPx10_ASAP7_75t_R FILLER_222_578 ();
 DECAPx6_ASAP7_75t_R FILLER_222_600 ();
 DECAPx10_ASAP7_75t_R FILLER_222_629 ();
 DECAPx10_ASAP7_75t_R FILLER_222_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_673 ();
 DECAPx4_ASAP7_75t_R FILLER_222_692 ();
 FILLER_ASAP7_75t_R FILLER_222_702 ();
 DECAPx1_ASAP7_75t_R FILLER_222_732 ();
 DECAPx2_ASAP7_75t_R FILLER_222_758 ();
 DECAPx1_ASAP7_75t_R FILLER_222_770 ();
 DECAPx2_ASAP7_75t_R FILLER_222_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_809 ();
 DECAPx4_ASAP7_75t_R FILLER_222_813 ();
 DECAPx2_ASAP7_75t_R FILLER_222_833 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_859 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_222_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_878 ();
 DECAPx1_ASAP7_75t_R FILLER_222_908 ();
 FILLERxp5_ASAP7_75t_R FILLER_222_912 ();
 DECAPx10_ASAP7_75t_R FILLER_223_2 ();
 DECAPx10_ASAP7_75t_R FILLER_223_24 ();
 DECAPx10_ASAP7_75t_R FILLER_223_46 ();
 DECAPx2_ASAP7_75t_R FILLER_223_68 ();
 DECAPx2_ASAP7_75t_R FILLER_223_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_106 ();
 DECAPx4_ASAP7_75t_R FILLER_223_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_170 ();
 FILLER_ASAP7_75t_R FILLER_223_177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_185 ();
 DECAPx10_ASAP7_75t_R FILLER_223_191 ();
 DECAPx4_ASAP7_75t_R FILLER_223_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_223 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_280 ();
 DECAPx2_ASAP7_75t_R FILLER_223_314 ();
 FILLER_ASAP7_75t_R FILLER_223_320 ();
 DECAPx1_ASAP7_75t_R FILLER_223_328 ();
 DECAPx2_ASAP7_75t_R FILLER_223_358 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_364 ();
 DECAPx10_ASAP7_75t_R FILLER_223_396 ();
 DECAPx2_ASAP7_75t_R FILLER_223_418 ();
 DECAPx2_ASAP7_75t_R FILLER_223_431 ();
 DECAPx2_ASAP7_75t_R FILLER_223_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_463 ();
 DECAPx1_ASAP7_75t_R FILLER_223_470 ();
 FILLER_ASAP7_75t_R FILLER_223_482 ();
 DECAPx10_ASAP7_75t_R FILLER_223_499 ();
 FILLER_ASAP7_75t_R FILLER_223_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_537 ();
 DECAPx10_ASAP7_75t_R FILLER_223_548 ();
 DECAPx10_ASAP7_75t_R FILLER_223_570 ();
 DECAPx6_ASAP7_75t_R FILLER_223_592 ();
 DECAPx2_ASAP7_75t_R FILLER_223_606 ();
 DECAPx10_ASAP7_75t_R FILLER_223_617 ();
 DECAPx6_ASAP7_75t_R FILLER_223_639 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_653 ();
 DECAPx10_ASAP7_75t_R FILLER_223_659 ();
 DECAPx6_ASAP7_75t_R FILLER_223_681 ();
 FILLER_ASAP7_75t_R FILLER_223_695 ();
 DECAPx6_ASAP7_75t_R FILLER_223_703 ();
 FILLER_ASAP7_75t_R FILLER_223_717 ();
 DECAPx4_ASAP7_75t_R FILLER_223_727 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_737 ();
 FILLER_ASAP7_75t_R FILLER_223_746 ();
 DECAPx2_ASAP7_75t_R FILLER_223_769 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_810 ();
 DECAPx2_ASAP7_75t_R FILLER_223_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_223_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_223_924 ();
 FILLER_ASAP7_75t_R FILLER_223_932 ();
 DECAPx10_ASAP7_75t_R FILLER_224_7 ();
 DECAPx10_ASAP7_75t_R FILLER_224_29 ();
 DECAPx6_ASAP7_75t_R FILLER_224_51 ();
 DECAPx2_ASAP7_75t_R FILLER_224_65 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_71 ();
 DECAPx10_ASAP7_75t_R FILLER_224_101 ();
 DECAPx2_ASAP7_75t_R FILLER_224_123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_129 ();
 DECAPx4_ASAP7_75t_R FILLER_224_158 ();
 DECAPx6_ASAP7_75t_R FILLER_224_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_215 ();
 DECAPx6_ASAP7_75t_R FILLER_224_278 ();
 DECAPx1_ASAP7_75t_R FILLER_224_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_302 ();
 DECAPx6_ASAP7_75t_R FILLER_224_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_320 ();
 DECAPx1_ASAP7_75t_R FILLER_224_341 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_345 ();
 DECAPx2_ASAP7_75t_R FILLER_224_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_355 ();
 DECAPx6_ASAP7_75t_R FILLER_224_362 ();
 DECAPx2_ASAP7_75t_R FILLER_224_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_391 ();
 DECAPx10_ASAP7_75t_R FILLER_224_399 ();
 DECAPx6_ASAP7_75t_R FILLER_224_421 ();
 FILLER_ASAP7_75t_R FILLER_224_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_444 ();
 DECAPx1_ASAP7_75t_R FILLER_224_458 ();
 FILLER_ASAP7_75t_R FILLER_224_464 ();
 FILLER_ASAP7_75t_R FILLER_224_472 ();
 DECAPx2_ASAP7_75t_R FILLER_224_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_520 ();
 DECAPx6_ASAP7_75t_R FILLER_224_524 ();
 DECAPx1_ASAP7_75t_R FILLER_224_538 ();
 DECAPx6_ASAP7_75t_R FILLER_224_558 ();
 DECAPx2_ASAP7_75t_R FILLER_224_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_578 ();
 DECAPx10_ASAP7_75t_R FILLER_224_606 ();
 DECAPx2_ASAP7_75t_R FILLER_224_628 ();
 FILLER_ASAP7_75t_R FILLER_224_634 ();
 DECAPx6_ASAP7_75t_R FILLER_224_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_705 ();
 FILLER_ASAP7_75t_R FILLER_224_718 ();
 FILLER_ASAP7_75t_R FILLER_224_743 ();
 DECAPx2_ASAP7_75t_R FILLER_224_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_757 ();
 DECAPx4_ASAP7_75t_R FILLER_224_778 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_842 ();
 DECAPx2_ASAP7_75t_R FILLER_224_887 ();
 FILLER_ASAP7_75t_R FILLER_224_893 ();
 DECAPx1_ASAP7_75t_R FILLER_224_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_906 ();
 DECAPx1_ASAP7_75t_R FILLER_224_910 ();
 FILLERxp5_ASAP7_75t_R FILLER_224_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_224_921 ();
 DECAPx10_ASAP7_75t_R FILLER_225_7 ();
 DECAPx10_ASAP7_75t_R FILLER_225_29 ();
 DECAPx10_ASAP7_75t_R FILLER_225_51 ();
 DECAPx2_ASAP7_75t_R FILLER_225_73 ();
 FILLER_ASAP7_75t_R FILLER_225_79 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_121 ();
 DECAPx2_ASAP7_75t_R FILLER_225_130 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_136 ();
 FILLER_ASAP7_75t_R FILLER_225_145 ();
 DECAPx2_ASAP7_75t_R FILLER_225_150 ();
 FILLER_ASAP7_75t_R FILLER_225_156 ();
 DECAPx2_ASAP7_75t_R FILLER_225_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_179 ();
 DECAPx6_ASAP7_75t_R FILLER_225_185 ();
 FILLER_ASAP7_75t_R FILLER_225_199 ();
 FILLER_ASAP7_75t_R FILLER_225_241 ();
 DECAPx4_ASAP7_75t_R FILLER_225_263 ();
 FILLER_ASAP7_75t_R FILLER_225_273 ();
 DECAPx10_ASAP7_75t_R FILLER_225_281 ();
 DECAPx10_ASAP7_75t_R FILLER_225_303 ();
 DECAPx10_ASAP7_75t_R FILLER_225_325 ();
 FILLER_ASAP7_75t_R FILLER_225_368 ();
 FILLER_ASAP7_75t_R FILLER_225_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_404 ();
 DECAPx10_ASAP7_75t_R FILLER_225_411 ();
 DECAPx6_ASAP7_75t_R FILLER_225_455 ();
 DECAPx2_ASAP7_75t_R FILLER_225_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_475 ();
 DECAPx2_ASAP7_75t_R FILLER_225_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_488 ();
 FILLER_ASAP7_75t_R FILLER_225_492 ();
 DECAPx4_ASAP7_75t_R FILLER_225_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_583 ();
 DECAPx10_ASAP7_75t_R FILLER_225_609 ();
 DECAPx2_ASAP7_75t_R FILLER_225_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_637 ();
 DECAPx4_ASAP7_75t_R FILLER_225_650 ();
 DECAPx1_ASAP7_75t_R FILLER_225_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_679 ();
 DECAPx1_ASAP7_75t_R FILLER_225_696 ();
 DECAPx2_ASAP7_75t_R FILLER_225_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_716 ();
 DECAPx2_ASAP7_75t_R FILLER_225_723 ();
 FILLER_ASAP7_75t_R FILLER_225_729 ();
 DECAPx10_ASAP7_75t_R FILLER_225_736 ();
 DECAPx10_ASAP7_75t_R FILLER_225_758 ();
 DECAPx10_ASAP7_75t_R FILLER_225_780 ();
 DECAPx1_ASAP7_75t_R FILLER_225_802 ();
 DECAPx10_ASAP7_75t_R FILLER_225_828 ();
 DECAPx2_ASAP7_75t_R FILLER_225_850 ();
 FILLER_ASAP7_75t_R FILLER_225_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_872 ();
 FILLER_ASAP7_75t_R FILLER_225_878 ();
 DECAPx10_ASAP7_75t_R FILLER_225_885 ();
 DECAPx4_ASAP7_75t_R FILLER_225_907 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_225_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_225_927 ();
 DECAPx10_ASAP7_75t_R FILLER_226_7 ();
 DECAPx10_ASAP7_75t_R FILLER_226_29 ();
 DECAPx10_ASAP7_75t_R FILLER_226_51 ();
 DECAPx4_ASAP7_75t_R FILLER_226_73 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_83 ();
 DECAPx2_ASAP7_75t_R FILLER_226_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_95 ();
 FILLER_ASAP7_75t_R FILLER_226_102 ();
 DECAPx4_ASAP7_75t_R FILLER_226_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_154 ();
 DECAPx10_ASAP7_75t_R FILLER_226_181 ();
 FILLER_ASAP7_75t_R FILLER_226_203 ();
 DECAPx1_ASAP7_75t_R FILLER_226_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_215 ();
 DECAPx10_ASAP7_75t_R FILLER_226_219 ();
 DECAPx6_ASAP7_75t_R FILLER_226_241 ();
 DECAPx1_ASAP7_75t_R FILLER_226_255 ();
 DECAPx2_ASAP7_75t_R FILLER_226_265 ();
 FILLER_ASAP7_75t_R FILLER_226_271 ();
 DECAPx10_ASAP7_75t_R FILLER_226_291 ();
 DECAPx1_ASAP7_75t_R FILLER_226_313 ();
 DECAPx6_ASAP7_75t_R FILLER_226_323 ();
 DECAPx2_ASAP7_75t_R FILLER_226_363 ();
 FILLER_ASAP7_75t_R FILLER_226_369 ();
 DECAPx4_ASAP7_75t_R FILLER_226_397 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_419 ();
 DECAPx2_ASAP7_75t_R FILLER_226_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_434 ();
 DECAPx6_ASAP7_75t_R FILLER_226_441 ();
 DECAPx2_ASAP7_75t_R FILLER_226_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_461 ();
 DECAPx4_ASAP7_75t_R FILLER_226_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_474 ();
 DECAPx2_ASAP7_75t_R FILLER_226_483 ();
 DECAPx10_ASAP7_75t_R FILLER_226_495 ();
 DECAPx10_ASAP7_75t_R FILLER_226_517 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_545 ();
 DECAPx2_ASAP7_75t_R FILLER_226_580 ();
 FILLER_ASAP7_75t_R FILLER_226_586 ();
 DECAPx6_ASAP7_75t_R FILLER_226_594 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_608 ();
 DECAPx2_ASAP7_75t_R FILLER_226_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_623 ();
 DECAPx6_ASAP7_75t_R FILLER_226_645 ();
 DECAPx2_ASAP7_75t_R FILLER_226_659 ();
 DECAPx10_ASAP7_75t_R FILLER_226_691 ();
 DECAPx6_ASAP7_75t_R FILLER_226_713 ();
 DECAPx1_ASAP7_75t_R FILLER_226_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_731 ();
 DECAPx10_ASAP7_75t_R FILLER_226_738 ();
 DECAPx2_ASAP7_75t_R FILLER_226_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_766 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_774 ();
 DECAPx6_ASAP7_75t_R FILLER_226_803 ();
 FILLER_ASAP7_75t_R FILLER_226_817 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_826 ();
 FILLER_ASAP7_75t_R FILLER_226_839 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_847 ();
 DECAPx2_ASAP7_75t_R FILLER_226_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_226_867 ();
 DECAPx1_ASAP7_75t_R FILLER_226_873 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_882 ();
 DECAPx4_ASAP7_75t_R FILLER_226_888 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_226_898 ();
 FILLER_ASAP7_75t_R FILLER_226_918 ();
 DECAPx10_ASAP7_75t_R FILLER_227_2 ();
 DECAPx10_ASAP7_75t_R FILLER_227_24 ();
 DECAPx10_ASAP7_75t_R FILLER_227_46 ();
 DECAPx10_ASAP7_75t_R FILLER_227_68 ();
 DECAPx10_ASAP7_75t_R FILLER_227_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_130 ();
 DECAPx10_ASAP7_75t_R FILLER_227_143 ();
 DECAPx1_ASAP7_75t_R FILLER_227_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_169 ();
 DECAPx4_ASAP7_75t_R FILLER_227_173 ();
 FILLER_ASAP7_75t_R FILLER_227_183 ();
 DECAPx1_ASAP7_75t_R FILLER_227_201 ();
 DECAPx10_ASAP7_75t_R FILLER_227_211 ();
 DECAPx10_ASAP7_75t_R FILLER_227_233 ();
 DECAPx2_ASAP7_75t_R FILLER_227_255 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_307 ();
 DECAPx2_ASAP7_75t_R FILLER_227_334 ();
 FILLER_ASAP7_75t_R FILLER_227_340 ();
 DECAPx1_ASAP7_75t_R FILLER_227_348 ();
 DECAPx6_ASAP7_75t_R FILLER_227_355 ();
 FILLER_ASAP7_75t_R FILLER_227_369 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_227_379 ();
 DECAPx2_ASAP7_75t_R FILLER_227_391 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_406 ();
 DECAPx1_ASAP7_75t_R FILLER_227_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_422 ();
 DECAPx1_ASAP7_75t_R FILLER_227_430 ();
 DECAPx2_ASAP7_75t_R FILLER_227_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_446 ();
 DECAPx1_ASAP7_75t_R FILLER_227_473 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_477 ();
 DECAPx1_ASAP7_75t_R FILLER_227_484 ();
 DECAPx6_ASAP7_75t_R FILLER_227_494 ();
 FILLER_ASAP7_75t_R FILLER_227_508 ();
 DECAPx6_ASAP7_75t_R FILLER_227_536 ();
 DECAPx2_ASAP7_75t_R FILLER_227_550 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_565 ();
 DECAPx10_ASAP7_75t_R FILLER_227_579 ();
 DECAPx10_ASAP7_75t_R FILLER_227_650 ();
 DECAPx2_ASAP7_75t_R FILLER_227_672 ();
 DECAPx10_ASAP7_75t_R FILLER_227_684 ();
 FILLER_ASAP7_75t_R FILLER_227_706 ();
 DECAPx2_ASAP7_75t_R FILLER_227_724 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_730 ();
 DECAPx6_ASAP7_75t_R FILLER_227_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_751 ();
 DECAPx1_ASAP7_75t_R FILLER_227_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_806 ();
 DECAPx1_ASAP7_75t_R FILLER_227_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_836 ();
 DECAPx1_ASAP7_75t_R FILLER_227_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_878 ();
 DECAPx1_ASAP7_75t_R FILLER_227_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_227_924 ();
 FILLER_ASAP7_75t_R FILLER_227_932 ();
 DECAPx10_ASAP7_75t_R FILLER_228_7 ();
 DECAPx10_ASAP7_75t_R FILLER_228_29 ();
 DECAPx10_ASAP7_75t_R FILLER_228_51 ();
 DECAPx1_ASAP7_75t_R FILLER_228_73 ();
 DECAPx10_ASAP7_75t_R FILLER_228_83 ();
 DECAPx10_ASAP7_75t_R FILLER_228_105 ();
 DECAPx6_ASAP7_75t_R FILLER_228_127 ();
 FILLER_ASAP7_75t_R FILLER_228_141 ();
 DECAPx6_ASAP7_75t_R FILLER_228_161 ();
 DECAPx1_ASAP7_75t_R FILLER_228_175 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_198 ();
 DECAPx2_ASAP7_75t_R FILLER_228_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_240 ();
 DECAPx2_ASAP7_75t_R FILLER_228_247 ();
 DECAPx10_ASAP7_75t_R FILLER_228_256 ();
 DECAPx1_ASAP7_75t_R FILLER_228_284 ();
 FILLER_ASAP7_75t_R FILLER_228_311 ();
 DECAPx1_ASAP7_75t_R FILLER_228_319 ();
 DECAPx10_ASAP7_75t_R FILLER_228_338 ();
 DECAPx10_ASAP7_75t_R FILLER_228_360 ();
 DECAPx6_ASAP7_75t_R FILLER_228_382 ();
 DECAPx2_ASAP7_75t_R FILLER_228_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_402 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_409 ();
 FILLER_ASAP7_75t_R FILLER_228_433 ();
 DECAPx2_ASAP7_75t_R FILLER_228_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_461 ();
 DECAPx1_ASAP7_75t_R FILLER_228_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_468 ();
 DECAPx10_ASAP7_75t_R FILLER_228_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_499 ();
 DECAPx6_ASAP7_75t_R FILLER_228_509 ();
 DECAPx2_ASAP7_75t_R FILLER_228_523 ();
 DECAPx10_ASAP7_75t_R FILLER_228_536 ();
 DECAPx10_ASAP7_75t_R FILLER_228_558 ();
 DECAPx6_ASAP7_75t_R FILLER_228_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_594 ();
 DECAPx2_ASAP7_75t_R FILLER_228_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_610 ();
 FILLER_ASAP7_75t_R FILLER_228_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_622 ();
 DECAPx2_ASAP7_75t_R FILLER_228_637 ();
 DECAPx4_ASAP7_75t_R FILLER_228_659 ();
 FILLER_ASAP7_75t_R FILLER_228_669 ();
 DECAPx2_ASAP7_75t_R FILLER_228_677 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_687 ();
 DECAPx6_ASAP7_75t_R FILLER_228_696 ();
 DECAPx2_ASAP7_75t_R FILLER_228_731 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_228_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_760 ();
 DECAPx1_ASAP7_75t_R FILLER_228_767 ();
 DECAPx1_ASAP7_75t_R FILLER_228_776 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_228_833 ();
 FILLER_ASAP7_75t_R FILLER_228_882 ();
 DECAPx10_ASAP7_75t_R FILLER_229_12 ();
 DECAPx10_ASAP7_75t_R FILLER_229_34 ();
 DECAPx4_ASAP7_75t_R FILLER_229_56 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_66 ();
 DECAPx10_ASAP7_75t_R FILLER_229_95 ();
 DECAPx4_ASAP7_75t_R FILLER_229_117 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_127 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_138 ();
 DECAPx1_ASAP7_75t_R FILLER_229_167 ();
 DECAPx1_ASAP7_75t_R FILLER_229_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_201 ();
 DECAPx2_ASAP7_75t_R FILLER_229_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_225 ();
 DECAPx10_ASAP7_75t_R FILLER_229_263 ();
 DECAPx4_ASAP7_75t_R FILLER_229_285 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_295 ();
 DECAPx2_ASAP7_75t_R FILLER_229_299 ();
 FILLER_ASAP7_75t_R FILLER_229_305 ();
 DECAPx2_ASAP7_75t_R FILLER_229_319 ();
 FILLER_ASAP7_75t_R FILLER_229_325 ();
 DECAPx2_ASAP7_75t_R FILLER_229_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_349 ();
 DECAPx2_ASAP7_75t_R FILLER_229_356 ();
 DECAPx10_ASAP7_75t_R FILLER_229_365 ();
 DECAPx10_ASAP7_75t_R FILLER_229_387 ();
 DECAPx6_ASAP7_75t_R FILLER_229_409 ();
 DECAPx4_ASAP7_75t_R FILLER_229_435 ();
 DECAPx1_ASAP7_75t_R FILLER_229_458 ();
 DECAPx2_ASAP7_75t_R FILLER_229_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_531 ();
 FILLER_ASAP7_75t_R FILLER_229_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_578 ();
 DECAPx2_ASAP7_75t_R FILLER_229_584 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_590 ();
 DECAPx10_ASAP7_75t_R FILLER_229_614 ();
 DECAPx4_ASAP7_75t_R FILLER_229_636 ();
 DECAPx2_ASAP7_75t_R FILLER_229_665 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_677 ();
 DECAPx1_ASAP7_75t_R FILLER_229_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_690 ();
 DECAPx2_ASAP7_75t_R FILLER_229_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_717 ();
 FILLER_ASAP7_75t_R FILLER_229_728 ();
 FILLER_ASAP7_75t_R FILLER_229_746 ();
 FILLER_ASAP7_75t_R FILLER_229_754 ();
 DECAPx10_ASAP7_75t_R FILLER_229_772 ();
 DECAPx4_ASAP7_75t_R FILLER_229_794 ();
 FILLER_ASAP7_75t_R FILLER_229_804 ();
 DECAPx4_ASAP7_75t_R FILLER_229_812 ();
 DECAPx6_ASAP7_75t_R FILLER_229_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_839 ();
 DECAPx6_ASAP7_75t_R FILLER_229_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_872 ();
 DECAPx2_ASAP7_75t_R FILLER_229_880 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_229_886 ();
 DECAPx2_ASAP7_75t_R FILLER_229_913 ();
 FILLERxp5_ASAP7_75t_R FILLER_229_919 ();
 FILLER_ASAP7_75t_R FILLER_229_927 ();
 DECAPx10_ASAP7_75t_R FILLER_230_7 ();
 DECAPx10_ASAP7_75t_R FILLER_230_29 ();
 DECAPx10_ASAP7_75t_R FILLER_230_51 ();
 DECAPx2_ASAP7_75t_R FILLER_230_73 ();
 FILLER_ASAP7_75t_R FILLER_230_88 ();
 DECAPx1_ASAP7_75t_R FILLER_230_113 ();
 DECAPx2_ASAP7_75t_R FILLER_230_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_143 ();
 DECAPx6_ASAP7_75t_R FILLER_230_159 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_173 ();
 DECAPx2_ASAP7_75t_R FILLER_230_180 ();
 DECAPx10_ASAP7_75t_R FILLER_230_189 ();
 DECAPx2_ASAP7_75t_R FILLER_230_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_223 ();
 FILLER_ASAP7_75t_R FILLER_230_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_244 ();
 DECAPx10_ASAP7_75t_R FILLER_230_278 ();
 DECAPx1_ASAP7_75t_R FILLER_230_300 ();
 DECAPx2_ASAP7_75t_R FILLER_230_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_320 ();
 DECAPx1_ASAP7_75t_R FILLER_230_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_339 ();
 FILLER_ASAP7_75t_R FILLER_230_366 ();
 DECAPx10_ASAP7_75t_R FILLER_230_400 ();
 DECAPx10_ASAP7_75t_R FILLER_230_422 ();
 DECAPx6_ASAP7_75t_R FILLER_230_444 ();
 DECAPx1_ASAP7_75t_R FILLER_230_458 ();
 DECAPx10_ASAP7_75t_R FILLER_230_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_486 ();
 DECAPx1_ASAP7_75t_R FILLER_230_498 ();
 DECAPx1_ASAP7_75t_R FILLER_230_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_512 ();
 DECAPx6_ASAP7_75t_R FILLER_230_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_553 ();
 DECAPx4_ASAP7_75t_R FILLER_230_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_575 ();
 DECAPx10_ASAP7_75t_R FILLER_230_594 ();
 DECAPx2_ASAP7_75t_R FILLER_230_616 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_622 ();
 DECAPx4_ASAP7_75t_R FILLER_230_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_645 ();
 FILLER_ASAP7_75t_R FILLER_230_664 ();
 FILLER_ASAP7_75t_R FILLER_230_678 ();
 DECAPx2_ASAP7_75t_R FILLER_230_692 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_698 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_716 ();
 DECAPx4_ASAP7_75t_R FILLER_230_725 ();
 DECAPx6_ASAP7_75t_R FILLER_230_741 ();
 DECAPx2_ASAP7_75t_R FILLER_230_755 ();
 DECAPx2_ASAP7_75t_R FILLER_230_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_773 ();
 DECAPx2_ASAP7_75t_R FILLER_230_785 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_791 ();
 DECAPx10_ASAP7_75t_R FILLER_230_812 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_834 ();
 DECAPx1_ASAP7_75t_R FILLER_230_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_230_844 ();
 FILLER_ASAP7_75t_R FILLER_230_852 ();
 DECAPx2_ASAP7_75t_R FILLER_230_864 ();
 DECAPx10_ASAP7_75t_R FILLER_230_875 ();
 DECAPx2_ASAP7_75t_R FILLER_230_897 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_903 ();
 FILLER_ASAP7_75t_R FILLER_230_911 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_230_931 ();
 DECAPx10_ASAP7_75t_R FILLER_231_2 ();
 DECAPx10_ASAP7_75t_R FILLER_231_24 ();
 DECAPx10_ASAP7_75t_R FILLER_231_46 ();
 DECAPx2_ASAP7_75t_R FILLER_231_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_108 ();
 DECAPx10_ASAP7_75t_R FILLER_231_141 ();
 DECAPx6_ASAP7_75t_R FILLER_231_163 ();
 FILLER_ASAP7_75t_R FILLER_231_177 ();
 FILLER_ASAP7_75t_R FILLER_231_185 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_190 ();
 DECAPx4_ASAP7_75t_R FILLER_231_196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_206 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_221 ();
 DECAPx6_ASAP7_75t_R FILLER_231_225 ();
 DECAPx2_ASAP7_75t_R FILLER_231_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_245 ();
 FILLER_ASAP7_75t_R FILLER_231_255 ();
 DECAPx6_ASAP7_75t_R FILLER_231_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_283 ();
 DECAPx2_ASAP7_75t_R FILLER_231_290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_296 ();
 DECAPx6_ASAP7_75t_R FILLER_231_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_328 ();
 DECAPx6_ASAP7_75t_R FILLER_231_332 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_352 ();
 DECAPx1_ASAP7_75t_R FILLER_231_358 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_362 ();
 DECAPx1_ASAP7_75t_R FILLER_231_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_388 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_410 ();
 DECAPx2_ASAP7_75t_R FILLER_231_422 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_428 ();
 DECAPx10_ASAP7_75t_R FILLER_231_437 ();
 FILLER_ASAP7_75t_R FILLER_231_459 ();
 DECAPx1_ASAP7_75t_R FILLER_231_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_473 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_486 ();
 DECAPx1_ASAP7_75t_R FILLER_231_515 ();
 FILLER_ASAP7_75t_R FILLER_231_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_553 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_562 ();
 DECAPx6_ASAP7_75t_R FILLER_231_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_583 ();
 DECAPx2_ASAP7_75t_R FILLER_231_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_602 ();
 DECAPx4_ASAP7_75t_R FILLER_231_619 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_629 ();
 DECAPx6_ASAP7_75t_R FILLER_231_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_652 ();
 FILLER_ASAP7_75t_R FILLER_231_666 ();
 DECAPx10_ASAP7_75t_R FILLER_231_674 ();
 DECAPx2_ASAP7_75t_R FILLER_231_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_702 ();
 DECAPx10_ASAP7_75t_R FILLER_231_709 ();
 DECAPx4_ASAP7_75t_R FILLER_231_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_741 ();
 DECAPx1_ASAP7_75t_R FILLER_231_748 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_776 ();
 FILLER_ASAP7_75t_R FILLER_231_785 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_832 ();
 DECAPx10_ASAP7_75t_R FILLER_231_846 ();
 DECAPx6_ASAP7_75t_R FILLER_231_868 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_231_882 ();
 DECAPx2_ASAP7_75t_R FILLER_231_897 ();
 FILLER_ASAP7_75t_R FILLER_231_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_231_933 ();
 DECAPx10_ASAP7_75t_R FILLER_232_2 ();
 DECAPx10_ASAP7_75t_R FILLER_232_24 ();
 DECAPx10_ASAP7_75t_R FILLER_232_46 ();
 DECAPx4_ASAP7_75t_R FILLER_232_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_78 ();
 FILLER_ASAP7_75t_R FILLER_232_94 ();
 DECAPx1_ASAP7_75t_R FILLER_232_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_118 ();
 DECAPx10_ASAP7_75t_R FILLER_232_130 ();
 FILLER_ASAP7_75t_R FILLER_232_152 ();
 DECAPx4_ASAP7_75t_R FILLER_232_198 ();
 DECAPx10_ASAP7_75t_R FILLER_232_234 ();
 DECAPx6_ASAP7_75t_R FILLER_232_256 ();
 FILLER_ASAP7_75t_R FILLER_232_270 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_298 ();
 DECAPx2_ASAP7_75t_R FILLER_232_307 ();
 FILLER_ASAP7_75t_R FILLER_232_313 ();
 DECAPx6_ASAP7_75t_R FILLER_232_341 ();
 DECAPx2_ASAP7_75t_R FILLER_232_377 ();
 DECAPx2_ASAP7_75t_R FILLER_232_394 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_426 ();
 DECAPx6_ASAP7_75t_R FILLER_232_444 ();
 DECAPx1_ASAP7_75t_R FILLER_232_458 ();
 DECAPx4_ASAP7_75t_R FILLER_232_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_474 ();
 DECAPx6_ASAP7_75t_R FILLER_232_483 ();
 DECAPx2_ASAP7_75t_R FILLER_232_497 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_503 ();
 DECAPx4_ASAP7_75t_R FILLER_232_507 ();
 FILLER_ASAP7_75t_R FILLER_232_517 ();
 DECAPx1_ASAP7_75t_R FILLER_232_525 ();
 DECAPx4_ASAP7_75t_R FILLER_232_571 ();
 DECAPx4_ASAP7_75t_R FILLER_232_596 ();
 FILLER_ASAP7_75t_R FILLER_232_606 ();
 DECAPx2_ASAP7_75t_R FILLER_232_625 ();
 FILLER_ASAP7_75t_R FILLER_232_631 ();
 DECAPx10_ASAP7_75t_R FILLER_232_647 ();
 DECAPx6_ASAP7_75t_R FILLER_232_669 ();
 DECAPx1_ASAP7_75t_R FILLER_232_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_693 ();
 DECAPx4_ASAP7_75t_R FILLER_232_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_707 ();
 DECAPx2_ASAP7_75t_R FILLER_232_719 ();
 DECAPx10_ASAP7_75t_R FILLER_232_737 ();
 DECAPx4_ASAP7_75t_R FILLER_232_759 ();
 DECAPx1_ASAP7_75t_R FILLER_232_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_788 ();
 FILLER_ASAP7_75t_R FILLER_232_796 ();
 DECAPx6_ASAP7_75t_R FILLER_232_824 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_838 ();
 DECAPx4_ASAP7_75t_R FILLER_232_852 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_232_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_232_902 ();
 FILLER_ASAP7_75t_R FILLER_232_932 ();
 DECAPx10_ASAP7_75t_R FILLER_233_2 ();
 DECAPx10_ASAP7_75t_R FILLER_233_24 ();
 DECAPx10_ASAP7_75t_R FILLER_233_46 ();
 DECAPx10_ASAP7_75t_R FILLER_233_68 ();
 DECAPx10_ASAP7_75t_R FILLER_233_90 ();
 DECAPx10_ASAP7_75t_R FILLER_233_112 ();
 DECAPx2_ASAP7_75t_R FILLER_233_134 ();
 FILLER_ASAP7_75t_R FILLER_233_181 ();
 DECAPx10_ASAP7_75t_R FILLER_233_212 ();
 DECAPx2_ASAP7_75t_R FILLER_233_234 ();
 FILLER_ASAP7_75t_R FILLER_233_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_248 ();
 DECAPx2_ASAP7_75t_R FILLER_233_255 ();
 FILLER_ASAP7_75t_R FILLER_233_261 ();
 DECAPx6_ASAP7_75t_R FILLER_233_269 ();
 FILLER_ASAP7_75t_R FILLER_233_310 ();
 DECAPx10_ASAP7_75t_R FILLER_233_324 ();
 DECAPx10_ASAP7_75t_R FILLER_233_346 ();
 DECAPx6_ASAP7_75t_R FILLER_233_368 ();
 DECAPx1_ASAP7_75t_R FILLER_233_382 ();
 DECAPx6_ASAP7_75t_R FILLER_233_392 ();
 DECAPx2_ASAP7_75t_R FILLER_233_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_412 ();
 DECAPx2_ASAP7_75t_R FILLER_233_427 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_433 ();
 DECAPx1_ASAP7_75t_R FILLER_233_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_443 ();
 DECAPx10_ASAP7_75t_R FILLER_233_453 ();
 DECAPx2_ASAP7_75t_R FILLER_233_475 ();
 DECAPx10_ASAP7_75t_R FILLER_233_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_515 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_542 ();
 DECAPx10_ASAP7_75t_R FILLER_233_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_596 ();
 DECAPx10_ASAP7_75t_R FILLER_233_603 ();
 DECAPx10_ASAP7_75t_R FILLER_233_625 ();
 DECAPx10_ASAP7_75t_R FILLER_233_647 ();
 DECAPx6_ASAP7_75t_R FILLER_233_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_689 ();
 DECAPx2_ASAP7_75t_R FILLER_233_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_706 ();
 DECAPx2_ASAP7_75t_R FILLER_233_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_733 ();
 DECAPx10_ASAP7_75t_R FILLER_233_746 ();
 DECAPx4_ASAP7_75t_R FILLER_233_768 ();
 DECAPx10_ASAP7_75t_R FILLER_233_788 ();
 FILLER_ASAP7_75t_R FILLER_233_810 ();
 DECAPx6_ASAP7_75t_R FILLER_233_815 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_845 ();
 FILLER_ASAP7_75t_R FILLER_233_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_233_867 ();
 FILLER_ASAP7_75t_R FILLER_233_876 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_233_927 ();
 DECAPx10_ASAP7_75t_R FILLER_234_2 ();
 DECAPx10_ASAP7_75t_R FILLER_234_24 ();
 DECAPx10_ASAP7_75t_R FILLER_234_46 ();
 DECAPx10_ASAP7_75t_R FILLER_234_68 ();
 DECAPx10_ASAP7_75t_R FILLER_234_90 ();
 DECAPx10_ASAP7_75t_R FILLER_234_112 ();
 DECAPx10_ASAP7_75t_R FILLER_234_163 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_185 ();
 DECAPx10_ASAP7_75t_R FILLER_234_203 ();
 DECAPx4_ASAP7_75t_R FILLER_234_225 ();
 FILLER_ASAP7_75t_R FILLER_234_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_263 ();
 DECAPx1_ASAP7_75t_R FILLER_234_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_310 ();
 DECAPx6_ASAP7_75t_R FILLER_234_337 ();
 FILLER_ASAP7_75t_R FILLER_234_351 ();
 FILLER_ASAP7_75t_R FILLER_234_359 ();
 DECAPx10_ASAP7_75t_R FILLER_234_373 ();
 DECAPx10_ASAP7_75t_R FILLER_234_395 ();
 DECAPx10_ASAP7_75t_R FILLER_234_417 ();
 DECAPx2_ASAP7_75t_R FILLER_234_439 ();
 FILLER_ASAP7_75t_R FILLER_234_445 ();
 DECAPx1_ASAP7_75t_R FILLER_234_454 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_458 ();
 DECAPx2_ASAP7_75t_R FILLER_234_476 ();
 DECAPx2_ASAP7_75t_R FILLER_234_492 ();
 FILLER_ASAP7_75t_R FILLER_234_498 ();
 DECAPx6_ASAP7_75t_R FILLER_234_508 ();
 DECAPx2_ASAP7_75t_R FILLER_234_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_528 ();
 DECAPx10_ASAP7_75t_R FILLER_234_538 ();
 DECAPx2_ASAP7_75t_R FILLER_234_560 ();
 DECAPx6_ASAP7_75t_R FILLER_234_574 ();
 DECAPx2_ASAP7_75t_R FILLER_234_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_613 ();
 DECAPx4_ASAP7_75t_R FILLER_234_626 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_234_636 ();
 DECAPx4_ASAP7_75t_R FILLER_234_648 ();
 FILLER_ASAP7_75t_R FILLER_234_658 ();
 DECAPx10_ASAP7_75t_R FILLER_234_689 ();
 DECAPx1_ASAP7_75t_R FILLER_234_711 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_715 ();
 DECAPx2_ASAP7_75t_R FILLER_234_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_747 ();
 DECAPx10_ASAP7_75t_R FILLER_234_780 ();
 DECAPx1_ASAP7_75t_R FILLER_234_802 ();
 DECAPx10_ASAP7_75t_R FILLER_234_816 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_234_933 ();
 DECAPx10_ASAP7_75t_R FILLER_235_2 ();
 DECAPx10_ASAP7_75t_R FILLER_235_24 ();
 DECAPx10_ASAP7_75t_R FILLER_235_46 ();
 DECAPx6_ASAP7_75t_R FILLER_235_68 ();
 FILLER_ASAP7_75t_R FILLER_235_82 ();
 FILLER_ASAP7_75t_R FILLER_235_90 ();
 DECAPx4_ASAP7_75t_R FILLER_235_98 ();
 FILLER_ASAP7_75t_R FILLER_235_108 ();
 FILLER_ASAP7_75t_R FILLER_235_116 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_135 ();
 DECAPx2_ASAP7_75t_R FILLER_235_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_148 ();
 DECAPx1_ASAP7_75t_R FILLER_235_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_156 ();
 DECAPx10_ASAP7_75t_R FILLER_235_163 ();
 DECAPx10_ASAP7_75t_R FILLER_235_185 ();
 DECAPx4_ASAP7_75t_R FILLER_235_207 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_246 ();
 FILLER_ASAP7_75t_R FILLER_235_288 ();
 FILLER_ASAP7_75t_R FILLER_235_293 ();
 DECAPx1_ASAP7_75t_R FILLER_235_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_302 ();
 DECAPx1_ASAP7_75t_R FILLER_235_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_313 ();
 DECAPx1_ASAP7_75t_R FILLER_235_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_328 ();
 DECAPx2_ASAP7_75t_R FILLER_235_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_338 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_371 ();
 DECAPx1_ASAP7_75t_R FILLER_235_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_387 ();
 DECAPx1_ASAP7_75t_R FILLER_235_408 ();
 DECAPx2_ASAP7_75t_R FILLER_235_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_424 ();
 FILLER_ASAP7_75t_R FILLER_235_431 ();
 FILLER_ASAP7_75t_R FILLER_235_442 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_447 ();
 DECAPx2_ASAP7_75t_R FILLER_235_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_477 ();
 DECAPx2_ASAP7_75t_R FILLER_235_486 ();
 FILLER_ASAP7_75t_R FILLER_235_492 ();
 DECAPx1_ASAP7_75t_R FILLER_235_519 ();
 DECAPx10_ASAP7_75t_R FILLER_235_526 ();
 DECAPx6_ASAP7_75t_R FILLER_235_548 ();
 DECAPx2_ASAP7_75t_R FILLER_235_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_585 ();
 FILLER_ASAP7_75t_R FILLER_235_598 ();
 DECAPx2_ASAP7_75t_R FILLER_235_616 ();
 FILLER_ASAP7_75t_R FILLER_235_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_632 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_658 ();
 DECAPx1_ASAP7_75t_R FILLER_235_670 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_674 ();
 DECAPx4_ASAP7_75t_R FILLER_235_689 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_699 ();
 DECAPx6_ASAP7_75t_R FILLER_235_706 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_235_720 ();
 DECAPx4_ASAP7_75t_R FILLER_235_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_736 ();
 DECAPx1_ASAP7_75t_R FILLER_235_761 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_765 ();
 DECAPx1_ASAP7_75t_R FILLER_235_778 ();
 DECAPx2_ASAP7_75t_R FILLER_235_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_804 ();
 DECAPx6_ASAP7_75t_R FILLER_235_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_822 ();
 DECAPx4_ASAP7_75t_R FILLER_235_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_865 ();
 FILLERxp5_ASAP7_75t_R FILLER_235_883 ();
 FILLER_ASAP7_75t_R FILLER_235_932 ();
 DECAPx10_ASAP7_75t_R FILLER_236_2 ();
 DECAPx10_ASAP7_75t_R FILLER_236_24 ();
 DECAPx10_ASAP7_75t_R FILLER_236_46 ();
 DECAPx1_ASAP7_75t_R FILLER_236_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_72 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_105 ();
 DECAPx1_ASAP7_75t_R FILLER_236_134 ();
 DECAPx2_ASAP7_75t_R FILLER_236_156 ();
 FILLER_ASAP7_75t_R FILLER_236_162 ();
 DECAPx6_ASAP7_75t_R FILLER_236_176 ();
 DECAPx1_ASAP7_75t_R FILLER_236_190 ();
 DECAPx1_ASAP7_75t_R FILLER_236_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_224 ();
 DECAPx6_ASAP7_75t_R FILLER_236_240 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_254 ();
 DECAPx2_ASAP7_75t_R FILLER_236_261 ();
 DECAPx10_ASAP7_75t_R FILLER_236_285 ();
 DECAPx10_ASAP7_75t_R FILLER_236_307 ();
 DECAPx1_ASAP7_75t_R FILLER_236_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_368 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_395 ();
 DECAPx4_ASAP7_75t_R FILLER_236_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_454 ();
 DECAPx1_ASAP7_75t_R FILLER_236_458 ();
 DECAPx1_ASAP7_75t_R FILLER_236_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_468 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_506 ();
 DECAPx2_ASAP7_75t_R FILLER_236_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_541 ();
 DECAPx2_ASAP7_75t_R FILLER_236_559 ();
 FILLER_ASAP7_75t_R FILLER_236_565 ();
 FILLER_ASAP7_75t_R FILLER_236_570 ();
 DECAPx10_ASAP7_75t_R FILLER_236_585 ();
 DECAPx2_ASAP7_75t_R FILLER_236_607 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_652 ();
 DECAPx2_ASAP7_75t_R FILLER_236_663 ();
 FILLER_ASAP7_75t_R FILLER_236_669 ();
 DECAPx1_ASAP7_75t_R FILLER_236_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_695 ();
 DECAPx10_ASAP7_75t_R FILLER_236_712 ();
 DECAPx6_ASAP7_75t_R FILLER_236_734 ();
 DECAPx1_ASAP7_75t_R FILLER_236_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_752 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_236_758 ();
 DECAPx1_ASAP7_75t_R FILLER_236_767 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_771 ();
 FILLER_ASAP7_75t_R FILLER_236_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_816 ();
 DECAPx1_ASAP7_75t_R FILLER_236_843 ();
 DECAPx1_ASAP7_75t_R FILLER_236_855 ();
 DECAPx4_ASAP7_75t_R FILLER_236_864 ();
 FILLER_ASAP7_75t_R FILLER_236_877 ();
 DECAPx1_ASAP7_75t_R FILLER_236_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_236_888 ();
 DECAPx10_ASAP7_75t_R FILLER_237_2 ();
 DECAPx10_ASAP7_75t_R FILLER_237_24 ();
 DECAPx10_ASAP7_75t_R FILLER_237_46 ();
 DECAPx4_ASAP7_75t_R FILLER_237_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_78 ();
 FILLER_ASAP7_75t_R FILLER_237_85 ();
 DECAPx2_ASAP7_75t_R FILLER_237_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_112 ();
 DECAPx1_ASAP7_75t_R FILLER_237_119 ();
 DECAPx2_ASAP7_75t_R FILLER_237_126 ();
 FILLER_ASAP7_75t_R FILLER_237_132 ();
 DECAPx6_ASAP7_75t_R FILLER_237_140 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_183 ();
 DECAPx10_ASAP7_75t_R FILLER_237_218 ();
 DECAPx10_ASAP7_75t_R FILLER_237_240 ();
 DECAPx10_ASAP7_75t_R FILLER_237_262 ();
 DECAPx6_ASAP7_75t_R FILLER_237_284 ();
 DECAPx1_ASAP7_75t_R FILLER_237_298 ();
 DECAPx4_ASAP7_75t_R FILLER_237_324 ();
 DECAPx6_ASAP7_75t_R FILLER_237_355 ();
 DECAPx1_ASAP7_75t_R FILLER_237_369 ();
 DECAPx2_ASAP7_75t_R FILLER_237_379 ();
 DECAPx1_ASAP7_75t_R FILLER_237_399 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_403 ();
 DECAPx6_ASAP7_75t_R FILLER_237_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_424 ();
 DECAPx10_ASAP7_75t_R FILLER_237_431 ();
 DECAPx6_ASAP7_75t_R FILLER_237_453 ();
 DECAPx1_ASAP7_75t_R FILLER_237_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_471 ();
 DECAPx4_ASAP7_75t_R FILLER_237_484 ();
 DECAPx2_ASAP7_75t_R FILLER_237_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_528 ();
 DECAPx1_ASAP7_75t_R FILLER_237_534 ();
 FILLER_ASAP7_75t_R FILLER_237_551 ();
 DECAPx6_ASAP7_75t_R FILLER_237_565 ();
 FILLER_ASAP7_75t_R FILLER_237_579 ();
 DECAPx4_ASAP7_75t_R FILLER_237_597 ();
 FILLER_ASAP7_75t_R FILLER_237_607 ();
 DECAPx2_ASAP7_75t_R FILLER_237_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_621 ();
 DECAPx6_ASAP7_75t_R FILLER_237_628 ();
 DECAPx1_ASAP7_75t_R FILLER_237_642 ();
 DECAPx1_ASAP7_75t_R FILLER_237_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_657 ();
 DECAPx6_ASAP7_75t_R FILLER_237_669 ();
 DECAPx2_ASAP7_75t_R FILLER_237_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_689 ();
 DECAPx10_ASAP7_75t_R FILLER_237_696 ();
 DECAPx1_ASAP7_75t_R FILLER_237_718 ();
 DECAPx1_ASAP7_75t_R FILLER_237_732 ();
 DECAPx6_ASAP7_75t_R FILLER_237_742 ();
 DECAPx2_ASAP7_75t_R FILLER_237_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_793 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_801 ();
 DECAPx1_ASAP7_75t_R FILLER_237_816 ();
 DECAPx1_ASAP7_75t_R FILLER_237_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_830 ();
 DECAPx10_ASAP7_75t_R FILLER_237_847 ();
 DECAPx6_ASAP7_75t_R FILLER_237_869 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_237_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_237_919 ();
 FILLER_ASAP7_75t_R FILLER_237_927 ();
 DECAPx10_ASAP7_75t_R FILLER_238_2 ();
 DECAPx10_ASAP7_75t_R FILLER_238_24 ();
 DECAPx10_ASAP7_75t_R FILLER_238_46 ();
 DECAPx10_ASAP7_75t_R FILLER_238_68 ();
 DECAPx6_ASAP7_75t_R FILLER_238_90 ();
 DECAPx10_ASAP7_75t_R FILLER_238_116 ();
 DECAPx10_ASAP7_75t_R FILLER_238_138 ();
 DECAPx2_ASAP7_75t_R FILLER_238_160 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_166 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_186 ();
 DECAPx2_ASAP7_75t_R FILLER_238_195 ();
 DECAPx4_ASAP7_75t_R FILLER_238_210 ();
 FILLER_ASAP7_75t_R FILLER_238_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_228 ();
 DECAPx1_ASAP7_75t_R FILLER_238_235 ();
 FILLER_ASAP7_75t_R FILLER_238_248 ();
 DECAPx10_ASAP7_75t_R FILLER_238_256 ();
 DECAPx2_ASAP7_75t_R FILLER_238_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_291 ();
 FILLER_ASAP7_75t_R FILLER_238_310 ();
 DECAPx10_ASAP7_75t_R FILLER_238_326 ();
 DECAPx10_ASAP7_75t_R FILLER_238_348 ();
 DECAPx4_ASAP7_75t_R FILLER_238_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_380 ();
 DECAPx1_ASAP7_75t_R FILLER_238_389 ();
 DECAPx10_ASAP7_75t_R FILLER_238_396 ();
 DECAPx10_ASAP7_75t_R FILLER_238_418 ();
 DECAPx6_ASAP7_75t_R FILLER_238_440 ();
 FILLER_ASAP7_75t_R FILLER_238_454 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_459 ();
 DECAPx10_ASAP7_75t_R FILLER_238_464 ();
 DECAPx10_ASAP7_75t_R FILLER_238_486 ();
 DECAPx2_ASAP7_75t_R FILLER_238_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_514 ();
 DECAPx1_ASAP7_75t_R FILLER_238_543 ();
 DECAPx2_ASAP7_75t_R FILLER_238_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_559 ();
 DECAPx2_ASAP7_75t_R FILLER_238_566 ();
 DECAPx10_ASAP7_75t_R FILLER_238_582 ();
 DECAPx10_ASAP7_75t_R FILLER_238_604 ();
 DECAPx10_ASAP7_75t_R FILLER_238_626 ();
 DECAPx4_ASAP7_75t_R FILLER_238_648 ();
 DECAPx10_ASAP7_75t_R FILLER_238_669 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_238_691 ();
 DECAPx2_ASAP7_75t_R FILLER_238_700 ();
 FILLER_ASAP7_75t_R FILLER_238_706 ();
 DECAPx4_ASAP7_75t_R FILLER_238_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_765 ();
 FILLER_ASAP7_75t_R FILLER_238_818 ();
 DECAPx6_ASAP7_75t_R FILLER_238_856 ();
 DECAPx1_ASAP7_75t_R FILLER_238_870 ();
 FILLER_ASAP7_75t_R FILLER_238_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_238_921 ();
 FILLER_ASAP7_75t_R FILLER_238_932 ();
 DECAPx10_ASAP7_75t_R FILLER_239_2 ();
 DECAPx10_ASAP7_75t_R FILLER_239_24 ();
 DECAPx10_ASAP7_75t_R FILLER_239_46 ();
 DECAPx4_ASAP7_75t_R FILLER_239_68 ();
 FILLER_ASAP7_75t_R FILLER_239_90 ();
 DECAPx10_ASAP7_75t_R FILLER_239_95 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_117 ();
 DECAPx10_ASAP7_75t_R FILLER_239_124 ();
 DECAPx10_ASAP7_75t_R FILLER_239_146 ();
 DECAPx1_ASAP7_75t_R FILLER_239_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_175 ();
 DECAPx10_ASAP7_75t_R FILLER_239_188 ();
 DECAPx2_ASAP7_75t_R FILLER_239_210 ();
 FILLER_ASAP7_75t_R FILLER_239_242 ();
 DECAPx1_ASAP7_75t_R FILLER_239_260 ();
 DECAPx4_ASAP7_75t_R FILLER_239_270 ();
 FILLER_ASAP7_75t_R FILLER_239_280 ();
 FILLER_ASAP7_75t_R FILLER_239_308 ();
 FILLER_ASAP7_75t_R FILLER_239_328 ();
 DECAPx4_ASAP7_75t_R FILLER_239_350 ();
 FILLER_ASAP7_75t_R FILLER_239_360 ();
 FILLER_ASAP7_75t_R FILLER_239_365 ();
 DECAPx2_ASAP7_75t_R FILLER_239_375 ();
 DECAPx6_ASAP7_75t_R FILLER_239_387 ();
 FILLER_ASAP7_75t_R FILLER_239_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_409 ();
 DECAPx6_ASAP7_75t_R FILLER_239_419 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_433 ();
 DECAPx10_ASAP7_75t_R FILLER_239_478 ();
 DECAPx10_ASAP7_75t_R FILLER_239_500 ();
 DECAPx1_ASAP7_75t_R FILLER_239_522 ();
 DECAPx2_ASAP7_75t_R FILLER_239_539 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_552 ();
 DECAPx2_ASAP7_75t_R FILLER_239_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_579 ();
 DECAPx4_ASAP7_75t_R FILLER_239_588 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_598 ();
 DECAPx1_ASAP7_75t_R FILLER_239_611 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_626 ();
 FILLER_ASAP7_75t_R FILLER_239_635 ();
 DECAPx10_ASAP7_75t_R FILLER_239_644 ();
 DECAPx6_ASAP7_75t_R FILLER_239_666 ();
 DECAPx6_ASAP7_75t_R FILLER_239_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_239_722 ();
 FILLER_ASAP7_75t_R FILLER_239_735 ();
 DECAPx6_ASAP7_75t_R FILLER_239_789 ();
 FILLER_ASAP7_75t_R FILLER_239_803 ();
 DECAPx10_ASAP7_75t_R FILLER_239_819 ();
 DECAPx1_ASAP7_75t_R FILLER_239_841 ();
 DECAPx1_ASAP7_75t_R FILLER_239_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_239_867 ();
 FILLER_ASAP7_75t_R FILLER_239_911 ();
 FILLER_ASAP7_75t_R FILLER_239_923 ();
 FILLER_ASAP7_75t_R FILLER_239_927 ();
 DECAPx10_ASAP7_75t_R FILLER_240_2 ();
 DECAPx10_ASAP7_75t_R FILLER_240_24 ();
 DECAPx10_ASAP7_75t_R FILLER_240_46 ();
 FILLER_ASAP7_75t_R FILLER_240_68 ();
 DECAPx4_ASAP7_75t_R FILLER_240_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_106 ();
 FILLER_ASAP7_75t_R FILLER_240_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_126 ();
 DECAPx10_ASAP7_75t_R FILLER_240_150 ();
 DECAPx6_ASAP7_75t_R FILLER_240_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_186 ();
 DECAPx10_ASAP7_75t_R FILLER_240_201 ();
 DECAPx2_ASAP7_75t_R FILLER_240_223 ();
 FILLER_ASAP7_75t_R FILLER_240_229 ();
 DECAPx2_ASAP7_75t_R FILLER_240_234 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_246 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_323 ();
 DECAPx2_ASAP7_75t_R FILLER_240_336 ();
 DECAPx4_ASAP7_75t_R FILLER_240_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_434 ();
 DECAPx1_ASAP7_75t_R FILLER_240_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_450 ();
 DECAPx2_ASAP7_75t_R FILLER_240_454 ();
 FILLER_ASAP7_75t_R FILLER_240_460 ();
 DECAPx1_ASAP7_75t_R FILLER_240_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_468 ();
 DECAPx4_ASAP7_75t_R FILLER_240_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_482 ();
 DECAPx10_ASAP7_75t_R FILLER_240_496 ();
 DECAPx2_ASAP7_75t_R FILLER_240_518 ();
 FILLER_ASAP7_75t_R FILLER_240_524 ();
 DECAPx10_ASAP7_75t_R FILLER_240_532 ();
 DECAPx6_ASAP7_75t_R FILLER_240_554 ();
 DECAPx4_ASAP7_75t_R FILLER_240_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_588 ();
 DECAPx6_ASAP7_75t_R FILLER_240_595 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_609 ();
 DECAPx1_ASAP7_75t_R FILLER_240_627 ();
 DECAPx10_ASAP7_75t_R FILLER_240_638 ();
 DECAPx4_ASAP7_75t_R FILLER_240_660 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_670 ();
 DECAPx2_ASAP7_75t_R FILLER_240_691 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_697 ();
 DECAPx4_ASAP7_75t_R FILLER_240_708 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_240_718 ();
 DECAPx1_ASAP7_75t_R FILLER_240_733 ();
 DECAPx4_ASAP7_75t_R FILLER_240_754 ();
 FILLER_ASAP7_75t_R FILLER_240_764 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_772 ();
 DECAPx10_ASAP7_75t_R FILLER_240_778 ();
 DECAPx6_ASAP7_75t_R FILLER_240_800 ();
 DECAPx1_ASAP7_75t_R FILLER_240_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_818 ();
 DECAPx6_ASAP7_75t_R FILLER_240_826 ();
 FILLER_ASAP7_75t_R FILLER_240_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_883 ();
 FILLER_ASAP7_75t_R FILLER_240_900 ();
 FILLERxp5_ASAP7_75t_R FILLER_240_927 ();
 DECAPx10_ASAP7_75t_R FILLER_241_2 ();
 DECAPx10_ASAP7_75t_R FILLER_241_24 ();
 DECAPx10_ASAP7_75t_R FILLER_241_46 ();
 DECAPx6_ASAP7_75t_R FILLER_241_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_82 ();
 DECAPx6_ASAP7_75t_R FILLER_241_88 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_102 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_129 ();
 DECAPx6_ASAP7_75t_R FILLER_241_170 ();
 FILLER_ASAP7_75t_R FILLER_241_210 ();
 DECAPx6_ASAP7_75t_R FILLER_241_226 ();
 DECAPx1_ASAP7_75t_R FILLER_241_240 ();
 DECAPx1_ASAP7_75t_R FILLER_241_292 ();
 FILLER_ASAP7_75t_R FILLER_241_302 ();
 DECAPx10_ASAP7_75t_R FILLER_241_307 ();
 DECAPx6_ASAP7_75t_R FILLER_241_329 ();
 FILLER_ASAP7_75t_R FILLER_241_343 ();
 DECAPx1_ASAP7_75t_R FILLER_241_383 ();
 DECAPx6_ASAP7_75t_R FILLER_241_390 ();
 DECAPx2_ASAP7_75t_R FILLER_241_404 ();
 DECAPx4_ASAP7_75t_R FILLER_241_413 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_423 ();
 DECAPx2_ASAP7_75t_R FILLER_241_429 ();
 FILLER_ASAP7_75t_R FILLER_241_435 ();
 DECAPx6_ASAP7_75t_R FILLER_241_459 ();
 DECAPx1_ASAP7_75t_R FILLER_241_473 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_514 ();
 DECAPx1_ASAP7_75t_R FILLER_241_528 ();
 DECAPx2_ASAP7_75t_R FILLER_241_539 ();
 DECAPx10_ASAP7_75t_R FILLER_241_555 ();
 DECAPx2_ASAP7_75t_R FILLER_241_577 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_583 ();
 DECAPx6_ASAP7_75t_R FILLER_241_614 ();
 FILLER_ASAP7_75t_R FILLER_241_628 ();
 DECAPx4_ASAP7_75t_R FILLER_241_637 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_653 ();
 DECAPx1_ASAP7_75t_R FILLER_241_662 ();
 DECAPx1_ASAP7_75t_R FILLER_241_699 ();
 DECAPx6_ASAP7_75t_R FILLER_241_709 ();
 FILLER_ASAP7_75t_R FILLER_241_735 ();
 DECAPx4_ASAP7_75t_R FILLER_241_743 ();
 DECAPx2_ASAP7_75t_R FILLER_241_765 ();
 FILLER_ASAP7_75t_R FILLER_241_771 ();
 FILLER_ASAP7_75t_R FILLER_241_780 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_798 ();
 DECAPx4_ASAP7_75t_R FILLER_241_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_819 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_241_831 ();
 DECAPx1_ASAP7_75t_R FILLER_241_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_241_914 ();
 FILLER_ASAP7_75t_R FILLER_241_927 ();
 DECAPx10_ASAP7_75t_R FILLER_242_2 ();
 DECAPx10_ASAP7_75t_R FILLER_242_24 ();
 DECAPx10_ASAP7_75t_R FILLER_242_46 ();
 DECAPx6_ASAP7_75t_R FILLER_242_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_82 ();
 DECAPx2_ASAP7_75t_R FILLER_242_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_97 ();
 FILLER_ASAP7_75t_R FILLER_242_120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_143 ();
 FILLER_ASAP7_75t_R FILLER_242_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_205 ();
 DECAPx10_ASAP7_75t_R FILLER_242_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_268 ();
 DECAPx2_ASAP7_75t_R FILLER_242_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_278 ();
 DECAPx10_ASAP7_75t_R FILLER_242_288 ();
 DECAPx10_ASAP7_75t_R FILLER_242_310 ();
 DECAPx1_ASAP7_75t_R FILLER_242_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_336 ();
 DECAPx2_ASAP7_75t_R FILLER_242_343 ();
 FILLER_ASAP7_75t_R FILLER_242_349 ();
 FILLER_ASAP7_75t_R FILLER_242_357 ();
 FILLER_ASAP7_75t_R FILLER_242_362 ();
 DECAPx10_ASAP7_75t_R FILLER_242_370 ();
 DECAPx10_ASAP7_75t_R FILLER_242_392 ();
 DECAPx2_ASAP7_75t_R FILLER_242_414 ();
 DECAPx2_ASAP7_75t_R FILLER_242_426 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_432 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_448 ();
 DECAPx2_ASAP7_75t_R FILLER_242_454 ();
 FILLER_ASAP7_75t_R FILLER_242_460 ();
 DECAPx6_ASAP7_75t_R FILLER_242_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_478 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_507 ();
 DECAPx10_ASAP7_75t_R FILLER_242_524 ();
 DECAPx6_ASAP7_75t_R FILLER_242_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_560 ();
 DECAPx1_ASAP7_75t_R FILLER_242_570 ();
 DECAPx1_ASAP7_75t_R FILLER_242_580 ();
 FILLER_ASAP7_75t_R FILLER_242_607 ();
 DECAPx2_ASAP7_75t_R FILLER_242_623 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_629 ();
 FILLER_ASAP7_75t_R FILLER_242_644 ();
 DECAPx10_ASAP7_75t_R FILLER_242_666 ();
 FILLER_ASAP7_75t_R FILLER_242_688 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_706 ();
 DECAPx10_ASAP7_75t_R FILLER_242_719 ();
 DECAPx4_ASAP7_75t_R FILLER_242_741 ();
 FILLER_ASAP7_75t_R FILLER_242_764 ();
 DECAPx6_ASAP7_75t_R FILLER_242_832 ();
 FILLER_ASAP7_75t_R FILLER_242_846 ();
 DECAPx4_ASAP7_75t_R FILLER_242_857 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_242_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_242_898 ();
 DECAPx10_ASAP7_75t_R FILLER_243_2 ();
 DECAPx10_ASAP7_75t_R FILLER_243_24 ();
 DECAPx10_ASAP7_75t_R FILLER_243_46 ();
 DECAPx2_ASAP7_75t_R FILLER_243_68 ();
 DECAPx4_ASAP7_75t_R FILLER_243_106 ();
 FILLER_ASAP7_75t_R FILLER_243_116 ();
 DECAPx10_ASAP7_75t_R FILLER_243_121 ();
 DECAPx2_ASAP7_75t_R FILLER_243_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_149 ();
 DECAPx4_ASAP7_75t_R FILLER_243_171 ();
 DECAPx4_ASAP7_75t_R FILLER_243_210 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_220 ();
 FILLER_ASAP7_75t_R FILLER_243_238 ();
 DECAPx2_ASAP7_75t_R FILLER_243_243 ();
 FILLER_ASAP7_75t_R FILLER_243_249 ();
 DECAPx10_ASAP7_75t_R FILLER_243_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_288 ();
 DECAPx6_ASAP7_75t_R FILLER_243_292 ();
 DECAPx1_ASAP7_75t_R FILLER_243_312 ();
 DECAPx2_ASAP7_75t_R FILLER_243_322 ();
 FILLER_ASAP7_75t_R FILLER_243_328 ();
 DECAPx1_ASAP7_75t_R FILLER_243_338 ();
 DECAPx10_ASAP7_75t_R FILLER_243_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_378 ();
 FILLER_ASAP7_75t_R FILLER_243_385 ();
 DECAPx10_ASAP7_75t_R FILLER_243_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_415 ();
 DECAPx10_ASAP7_75t_R FILLER_243_436 ();
 DECAPx2_ASAP7_75t_R FILLER_243_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_467 ();
 DECAPx1_ASAP7_75t_R FILLER_243_479 ();
 DECAPx1_ASAP7_75t_R FILLER_243_491 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_495 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_499 ();
 DECAPx6_ASAP7_75t_R FILLER_243_516 ();
 FILLER_ASAP7_75t_R FILLER_243_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_545 ();
 DECAPx6_ASAP7_75t_R FILLER_243_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_575 ();
 DECAPx2_ASAP7_75t_R FILLER_243_583 ();
 DECAPx2_ASAP7_75t_R FILLER_243_627 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_633 ();
 DECAPx2_ASAP7_75t_R FILLER_243_640 ();
 FILLER_ASAP7_75t_R FILLER_243_646 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_654 ();
 DECAPx10_ASAP7_75t_R FILLER_243_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_697 ();
 FILLER_ASAP7_75t_R FILLER_243_704 ();
 DECAPx2_ASAP7_75t_R FILLER_243_716 ();
 FILLER_ASAP7_75t_R FILLER_243_722 ();
 DECAPx6_ASAP7_75t_R FILLER_243_730 ();
 DECAPx1_ASAP7_75t_R FILLER_243_744 ();
 DECAPx2_ASAP7_75t_R FILLER_243_774 ();
 FILLER_ASAP7_75t_R FILLER_243_789 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_243_802 ();
 DECAPx4_ASAP7_75t_R FILLER_243_808 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_818 ();
 DECAPx2_ASAP7_75t_R FILLER_243_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_833 ();
 DECAPx6_ASAP7_75t_R FILLER_243_847 ();
 DECAPx1_ASAP7_75t_R FILLER_243_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_898 ();
 FILLERxp5_ASAP7_75t_R FILLER_243_924 ();
 FILLER_ASAP7_75t_R FILLER_243_927 ();
 DECAPx10_ASAP7_75t_R FILLER_244_2 ();
 DECAPx10_ASAP7_75t_R FILLER_244_24 ();
 DECAPx10_ASAP7_75t_R FILLER_244_46 ();
 DECAPx4_ASAP7_75t_R FILLER_244_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_87 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_91 ();
 DECAPx10_ASAP7_75t_R FILLER_244_100 ();
 DECAPx10_ASAP7_75t_R FILLER_244_128 ();
 DECAPx10_ASAP7_75t_R FILLER_244_150 ();
 DECAPx2_ASAP7_75t_R FILLER_244_172 ();
 DECAPx4_ASAP7_75t_R FILLER_244_206 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_216 ();
 DECAPx4_ASAP7_75t_R FILLER_244_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_250 ();
 DECAPx4_ASAP7_75t_R FILLER_244_279 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_299 ();
 DECAPx1_ASAP7_75t_R FILLER_244_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_341 ();
 DECAPx2_ASAP7_75t_R FILLER_244_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_402 ();
 DECAPx1_ASAP7_75t_R FILLER_244_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_419 ();
 DECAPx6_ASAP7_75t_R FILLER_244_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_440 ();
 DECAPx4_ASAP7_75t_R FILLER_244_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_458 ();
 DECAPx10_ASAP7_75t_R FILLER_244_478 ();
 DECAPx4_ASAP7_75t_R FILLER_244_500 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_522 ();
 DECAPx4_ASAP7_75t_R FILLER_244_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_538 ();
 DECAPx1_ASAP7_75t_R FILLER_244_584 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_588 ();
 DECAPx1_ASAP7_75t_R FILLER_244_595 ();
 DECAPx6_ASAP7_75t_R FILLER_244_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_629 ();
 DECAPx4_ASAP7_75t_R FILLER_244_638 ();
 DECAPx1_ASAP7_75t_R FILLER_244_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_658 ();
 DECAPx2_ASAP7_75t_R FILLER_244_665 ();
 FILLER_ASAP7_75t_R FILLER_244_671 ();
 FILLER_ASAP7_75t_R FILLER_244_679 ();
 DECAPx10_ASAP7_75t_R FILLER_244_687 ();
 DECAPx1_ASAP7_75t_R FILLER_244_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_713 ();
 DECAPx1_ASAP7_75t_R FILLER_244_720 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_739 ();
 DECAPx4_ASAP7_75t_R FILLER_244_765 ();
 DECAPx2_ASAP7_75t_R FILLER_244_790 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_244_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_806 ();
 DECAPx2_ASAP7_75t_R FILLER_244_814 ();
 FILLER_ASAP7_75t_R FILLER_244_820 ();
 DECAPx2_ASAP7_75t_R FILLER_244_856 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_244_928 ();
 DECAPx10_ASAP7_75t_R FILLER_245_2 ();
 DECAPx10_ASAP7_75t_R FILLER_245_24 ();
 DECAPx10_ASAP7_75t_R FILLER_245_46 ();
 DECAPx10_ASAP7_75t_R FILLER_245_68 ();
 DECAPx10_ASAP7_75t_R FILLER_245_90 ();
 DECAPx6_ASAP7_75t_R FILLER_245_112 ();
 DECAPx1_ASAP7_75t_R FILLER_245_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_130 ();
 DECAPx2_ASAP7_75t_R FILLER_245_137 ();
 FILLER_ASAP7_75t_R FILLER_245_143 ();
 DECAPx10_ASAP7_75t_R FILLER_245_151 ();
 DECAPx10_ASAP7_75t_R FILLER_245_176 ();
 DECAPx4_ASAP7_75t_R FILLER_245_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_208 ();
 DECAPx6_ASAP7_75t_R FILLER_245_215 ();
 DECAPx1_ASAP7_75t_R FILLER_245_229 ();
 DECAPx6_ASAP7_75t_R FILLER_245_245 ();
 DECAPx1_ASAP7_75t_R FILLER_245_259 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_272 ();
 DECAPx1_ASAP7_75t_R FILLER_245_322 ();
 DECAPx1_ASAP7_75t_R FILLER_245_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_351 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_378 ();
 DECAPx10_ASAP7_75t_R FILLER_245_420 ();
 DECAPx1_ASAP7_75t_R FILLER_245_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_450 ();
 DECAPx4_ASAP7_75t_R FILLER_245_479 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_489 ();
 DECAPx4_ASAP7_75t_R FILLER_245_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_508 ();
 DECAPx2_ASAP7_75t_R FILLER_245_537 ();
 FILLER_ASAP7_75t_R FILLER_245_543 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_571 ();
 DECAPx6_ASAP7_75t_R FILLER_245_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_594 ();
 DECAPx2_ASAP7_75t_R FILLER_245_609 ();
 DECAPx4_ASAP7_75t_R FILLER_245_628 ();
 DECAPx10_ASAP7_75t_R FILLER_245_644 ();
 DECAPx10_ASAP7_75t_R FILLER_245_666 ();
 DECAPx10_ASAP7_75t_R FILLER_245_688 ();
 DECAPx1_ASAP7_75t_R FILLER_245_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_730 ();
 DECAPx1_ASAP7_75t_R FILLER_245_738 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_742 ();
 DECAPx10_ASAP7_75t_R FILLER_245_750 ();
 DECAPx10_ASAP7_75t_R FILLER_245_772 ();
 DECAPx1_ASAP7_75t_R FILLER_245_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_245_798 ();
 FILLER_ASAP7_75t_R FILLER_245_807 ();
 DECAPx10_ASAP7_75t_R FILLER_245_817 ();
 DECAPx2_ASAP7_75t_R FILLER_245_839 ();
 DECAPx4_ASAP7_75t_R FILLER_245_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_245_858 ();
 DECAPx10_ASAP7_75t_R FILLER_246_2 ();
 DECAPx10_ASAP7_75t_R FILLER_246_24 ();
 DECAPx10_ASAP7_75t_R FILLER_246_46 ();
 DECAPx10_ASAP7_75t_R FILLER_246_68 ();
 DECAPx4_ASAP7_75t_R FILLER_246_90 ();
 FILLER_ASAP7_75t_R FILLER_246_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_123 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_132 ();
 FILLER_ASAP7_75t_R FILLER_246_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_159 ();
 FILLER_ASAP7_75t_R FILLER_246_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_168 ();
 DECAPx10_ASAP7_75t_R FILLER_246_189 ();
 DECAPx6_ASAP7_75t_R FILLER_246_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_225 ();
 DECAPx2_ASAP7_75t_R FILLER_246_264 ();
 DECAPx4_ASAP7_75t_R FILLER_246_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_335 ();
 DECAPx4_ASAP7_75t_R FILLER_246_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_353 ();
 DECAPx1_ASAP7_75t_R FILLER_246_362 ();
 DECAPx6_ASAP7_75t_R FILLER_246_369 ();
 DECAPx1_ASAP7_75t_R FILLER_246_383 ();
 DECAPx4_ASAP7_75t_R FILLER_246_416 ();
 DECAPx1_ASAP7_75t_R FILLER_246_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_459 ();
 DECAPx10_ASAP7_75t_R FILLER_246_464 ();
 DECAPx10_ASAP7_75t_R FILLER_246_486 ();
 DECAPx2_ASAP7_75t_R FILLER_246_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_514 ();
 DECAPx10_ASAP7_75t_R FILLER_246_525 ();
 DECAPx2_ASAP7_75t_R FILLER_246_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_553 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_557 ();
 DECAPx4_ASAP7_75t_R FILLER_246_563 ();
 FILLER_ASAP7_75t_R FILLER_246_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_583 ();
 DECAPx2_ASAP7_75t_R FILLER_246_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_613 ();
 FILLER_ASAP7_75t_R FILLER_246_629 ();
 DECAPx10_ASAP7_75t_R FILLER_246_651 ();
 DECAPx4_ASAP7_75t_R FILLER_246_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_683 ();
 DECAPx6_ASAP7_75t_R FILLER_246_696 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_710 ();
 DECAPx6_ASAP7_75t_R FILLER_246_716 ();
 FILLER_ASAP7_75t_R FILLER_246_730 ();
 DECAPx2_ASAP7_75t_R FILLER_246_739 ();
 FILLER_ASAP7_75t_R FILLER_246_753 ();
 FILLER_ASAP7_75t_R FILLER_246_762 ();
 DECAPx6_ASAP7_75t_R FILLER_246_778 ();
 DECAPx2_ASAP7_75t_R FILLER_246_792 ();
 DECAPx10_ASAP7_75t_R FILLER_246_808 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_246_837 ();
 DECAPx6_ASAP7_75t_R FILLER_246_852 ();
 FILLER_ASAP7_75t_R FILLER_246_880 ();
 FILLERxp5_ASAP7_75t_R FILLER_246_933 ();
 DECAPx10_ASAP7_75t_R FILLER_247_2 ();
 DECAPx10_ASAP7_75t_R FILLER_247_24 ();
 DECAPx10_ASAP7_75t_R FILLER_247_46 ();
 DECAPx6_ASAP7_75t_R FILLER_247_68 ();
 DECAPx2_ASAP7_75t_R FILLER_247_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_94 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_124 ();
 FILLER_ASAP7_75t_R FILLER_247_171 ();
 DECAPx4_ASAP7_75t_R FILLER_247_179 ();
 FILLER_ASAP7_75t_R FILLER_247_189 ();
 DECAPx1_ASAP7_75t_R FILLER_247_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_204 ();
 DECAPx4_ASAP7_75t_R FILLER_247_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_218 ();
 FILLER_ASAP7_75t_R FILLER_247_256 ();
 DECAPx6_ASAP7_75t_R FILLER_247_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_278 ();
 DECAPx10_ASAP7_75t_R FILLER_247_288 ();
 FILLER_ASAP7_75t_R FILLER_247_310 ();
 DECAPx1_ASAP7_75t_R FILLER_247_326 ();
 DECAPx2_ASAP7_75t_R FILLER_247_341 ();
 DECAPx10_ASAP7_75t_R FILLER_247_353 ();
 DECAPx4_ASAP7_75t_R FILLER_247_375 ();
 FILLER_ASAP7_75t_R FILLER_247_385 ();
 DECAPx2_ASAP7_75t_R FILLER_247_393 ();
 DECAPx6_ASAP7_75t_R FILLER_247_402 ();
 DECAPx2_ASAP7_75t_R FILLER_247_416 ();
 DECAPx2_ASAP7_75t_R FILLER_247_441 ();
 DECAPx10_ASAP7_75t_R FILLER_247_450 ();
 DECAPx4_ASAP7_75t_R FILLER_247_472 ();
 DECAPx2_ASAP7_75t_R FILLER_247_492 ();
 DECAPx6_ASAP7_75t_R FILLER_247_505 ();
 DECAPx1_ASAP7_75t_R FILLER_247_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_523 ();
 DECAPx2_ASAP7_75t_R FILLER_247_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_536 ();
 DECAPx10_ASAP7_75t_R FILLER_247_551 ();
 DECAPx2_ASAP7_75t_R FILLER_247_579 ();
 DECAPx4_ASAP7_75t_R FILLER_247_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_608 ();
 DECAPx4_ASAP7_75t_R FILLER_247_635 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_645 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_655 ();
 DECAPx4_ASAP7_75t_R FILLER_247_678 ();
 DECAPx4_ASAP7_75t_R FILLER_247_716 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_726 ();
 DECAPx10_ASAP7_75t_R FILLER_247_781 ();
 DECAPx4_ASAP7_75t_R FILLER_247_803 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_247_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_852 ();
 DECAPx1_ASAP7_75t_R FILLER_247_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_899 ();
 FILLERxp5_ASAP7_75t_R FILLER_247_927 ();
 DECAPx10_ASAP7_75t_R FILLER_248_2 ();
 DECAPx10_ASAP7_75t_R FILLER_248_24 ();
 DECAPx10_ASAP7_75t_R FILLER_248_46 ();
 DECAPx2_ASAP7_75t_R FILLER_248_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_106 ();
 DECAPx10_ASAP7_75t_R FILLER_248_116 ();
 DECAPx4_ASAP7_75t_R FILLER_248_138 ();
 FILLER_ASAP7_75t_R FILLER_248_148 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_156 ();
 DECAPx4_ASAP7_75t_R FILLER_248_171 ();
 FILLER_ASAP7_75t_R FILLER_248_181 ();
 DECAPx2_ASAP7_75t_R FILLER_248_217 ();
 DECAPx6_ASAP7_75t_R FILLER_248_238 ();
 FILLER_ASAP7_75t_R FILLER_248_252 ();
 DECAPx6_ASAP7_75t_R FILLER_248_262 ();
 DECAPx2_ASAP7_75t_R FILLER_248_276 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_282 ();
 DECAPx10_ASAP7_75t_R FILLER_248_286 ();
 FILLER_ASAP7_75t_R FILLER_248_329 ();
 DECAPx10_ASAP7_75t_R FILLER_248_383 ();
 DECAPx4_ASAP7_75t_R FILLER_248_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_415 ();
 DECAPx1_ASAP7_75t_R FILLER_248_427 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_431 ();
 DECAPx10_ASAP7_75t_R FILLER_248_435 ();
 DECAPx1_ASAP7_75t_R FILLER_248_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_461 ();
 DECAPx2_ASAP7_75t_R FILLER_248_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_509 ();
 DECAPx1_ASAP7_75t_R FILLER_248_516 ();
 DECAPx1_ASAP7_75t_R FILLER_248_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_532 ();
 DECAPx2_ASAP7_75t_R FILLER_248_540 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_546 ();
 DECAPx1_ASAP7_75t_R FILLER_248_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_560 ();
 DECAPx4_ASAP7_75t_R FILLER_248_583 ();
 FILLER_ASAP7_75t_R FILLER_248_593 ();
 DECAPx2_ASAP7_75t_R FILLER_248_610 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_616 ();
 DECAPx2_ASAP7_75t_R FILLER_248_625 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_248_631 ();
 DECAPx2_ASAP7_75t_R FILLER_248_642 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_654 ();
 FILLER_ASAP7_75t_R FILLER_248_670 ();
 DECAPx1_ASAP7_75t_R FILLER_248_694 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_708 ();
 DECAPx6_ASAP7_75t_R FILLER_248_719 ();
 DECAPx2_ASAP7_75t_R FILLER_248_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_739 ();
 DECAPx6_ASAP7_75t_R FILLER_248_749 ();
 DECAPx1_ASAP7_75t_R FILLER_248_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_767 ();
 DECAPx4_ASAP7_75t_R FILLER_248_771 ();
 FILLER_ASAP7_75t_R FILLER_248_781 ();
 FILLER_ASAP7_75t_R FILLER_248_797 ();
 FILLER_ASAP7_75t_R FILLER_248_830 ();
 DECAPx6_ASAP7_75t_R FILLER_248_848 ();
 DECAPx1_ASAP7_75t_R FILLER_248_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_248_928 ();
 DECAPx10_ASAP7_75t_R FILLER_249_2 ();
 DECAPx10_ASAP7_75t_R FILLER_249_24 ();
 DECAPx10_ASAP7_75t_R FILLER_249_46 ();
 DECAPx6_ASAP7_75t_R FILLER_249_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_82 ();
 FILLER_ASAP7_75t_R FILLER_249_89 ();
 DECAPx6_ASAP7_75t_R FILLER_249_94 ();
 DECAPx10_ASAP7_75t_R FILLER_249_114 ();
 DECAPx6_ASAP7_75t_R FILLER_249_136 ();
 DECAPx1_ASAP7_75t_R FILLER_249_150 ();
 DECAPx2_ASAP7_75t_R FILLER_249_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_186 ();
 DECAPx1_ASAP7_75t_R FILLER_249_193 ();
 FILLER_ASAP7_75t_R FILLER_249_217 ();
 DECAPx10_ASAP7_75t_R FILLER_249_225 ();
 DECAPx6_ASAP7_75t_R FILLER_249_247 ();
 FILLER_ASAP7_75t_R FILLER_249_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_295 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_249_302 ();
 DECAPx10_ASAP7_75t_R FILLER_249_311 ();
 DECAPx4_ASAP7_75t_R FILLER_249_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_343 ();
 DECAPx2_ASAP7_75t_R FILLER_249_353 ();
 FILLER_ASAP7_75t_R FILLER_249_359 ();
 DECAPx6_ASAP7_75t_R FILLER_249_390 ();
 DECAPx1_ASAP7_75t_R FILLER_249_404 ();
 DECAPx2_ASAP7_75t_R FILLER_249_414 ();
 DECAPx6_ASAP7_75t_R FILLER_249_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_452 ();
 DECAPx2_ASAP7_75t_R FILLER_249_456 ();
 FILLER_ASAP7_75t_R FILLER_249_487 ();
 DECAPx1_ASAP7_75t_R FILLER_249_492 ();
 FILLER_ASAP7_75t_R FILLER_249_505 ();
 DECAPx1_ASAP7_75t_R FILLER_249_514 ();
 FILLER_ASAP7_75t_R FILLER_249_544 ();
 DECAPx4_ASAP7_75t_R FILLER_249_572 ();
 DECAPx10_ASAP7_75t_R FILLER_249_588 ();
 DECAPx6_ASAP7_75t_R FILLER_249_610 ();
 DECAPx1_ASAP7_75t_R FILLER_249_637 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_641 ();
 FILLER_ASAP7_75t_R FILLER_249_695 ();
 DECAPx1_ASAP7_75t_R FILLER_249_704 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_708 ();
 DECAPx10_ASAP7_75t_R FILLER_249_715 ();
 DECAPx10_ASAP7_75t_R FILLER_249_737 ();
 DECAPx1_ASAP7_75t_R FILLER_249_759 ();
 DECAPx2_ASAP7_75t_R FILLER_249_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_776 ();
 DECAPx2_ASAP7_75t_R FILLER_249_789 ();
 DECAPx2_ASAP7_75t_R FILLER_249_805 ();
 FILLER_ASAP7_75t_R FILLER_249_816 ();
 DECAPx10_ASAP7_75t_R FILLER_249_821 ();
 DECAPx6_ASAP7_75t_R FILLER_249_843 ();
 FILLER_ASAP7_75t_R FILLER_249_857 ();
 DECAPx1_ASAP7_75t_R FILLER_249_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_249_919 ();
 FILLER_ASAP7_75t_R FILLER_249_927 ();
 DECAPx10_ASAP7_75t_R FILLER_250_2 ();
 DECAPx10_ASAP7_75t_R FILLER_250_24 ();
 DECAPx10_ASAP7_75t_R FILLER_250_46 ();
 DECAPx10_ASAP7_75t_R FILLER_250_68 ();
 DECAPx2_ASAP7_75t_R FILLER_250_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_96 ();
 DECAPx10_ASAP7_75t_R FILLER_250_128 ();
 DECAPx6_ASAP7_75t_R FILLER_250_150 ();
 DECAPx1_ASAP7_75t_R FILLER_250_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_168 ();
 DECAPx4_ASAP7_75t_R FILLER_250_172 ();
 DECAPx2_ASAP7_75t_R FILLER_250_208 ();
 FILLER_ASAP7_75t_R FILLER_250_214 ();
 DECAPx10_ASAP7_75t_R FILLER_250_222 ();
 DECAPx6_ASAP7_75t_R FILLER_250_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_258 ();
 DECAPx6_ASAP7_75t_R FILLER_250_317 ();
 FILLER_ASAP7_75t_R FILLER_250_331 ();
 DECAPx4_ASAP7_75t_R FILLER_250_342 ();
 FILLER_ASAP7_75t_R FILLER_250_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_378 ();
 FILLER_ASAP7_75t_R FILLER_250_385 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_436 ();
 DECAPx2_ASAP7_75t_R FILLER_250_440 ();
 FILLER_ASAP7_75t_R FILLER_250_446 ();
 FILLER_ASAP7_75t_R FILLER_250_467 ();
 DECAPx4_ASAP7_75t_R FILLER_250_482 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_492 ();
 DECAPx2_ASAP7_75t_R FILLER_250_501 ();
 DECAPx4_ASAP7_75t_R FILLER_250_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_523 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_543 ();
 DECAPx6_ASAP7_75t_R FILLER_250_565 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_579 ();
 DECAPx2_ASAP7_75t_R FILLER_250_586 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_592 ();
 DECAPx10_ASAP7_75t_R FILLER_250_601 ();
 DECAPx10_ASAP7_75t_R FILLER_250_623 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_645 ();
 DECAPx10_ASAP7_75t_R FILLER_250_654 ();
 DECAPx2_ASAP7_75t_R FILLER_250_676 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_250_682 ();
 DECAPx6_ASAP7_75t_R FILLER_250_691 ();
 DECAPx2_ASAP7_75t_R FILLER_250_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_711 ();
 FILLER_ASAP7_75t_R FILLER_250_718 ();
 DECAPx1_ASAP7_75t_R FILLER_250_725 ();
 DECAPx10_ASAP7_75t_R FILLER_250_735 ();
 FILLER_ASAP7_75t_R FILLER_250_757 ();
 DECAPx1_ASAP7_75t_R FILLER_250_785 ();
 DECAPx10_ASAP7_75t_R FILLER_250_815 ();
 DECAPx4_ASAP7_75t_R FILLER_250_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_250_847 ();
 DECAPx2_ASAP7_75t_R FILLER_250_874 ();
 FILLER_ASAP7_75t_R FILLER_250_911 ();
 DECAPx10_ASAP7_75t_R FILLER_251_2 ();
 DECAPx10_ASAP7_75t_R FILLER_251_24 ();
 DECAPx10_ASAP7_75t_R FILLER_251_46 ();
 DECAPx10_ASAP7_75t_R FILLER_251_68 ();
 DECAPx6_ASAP7_75t_R FILLER_251_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_104 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_111 ();
 DECAPx1_ASAP7_75t_R FILLER_251_117 ();
 DECAPx10_ASAP7_75t_R FILLER_251_152 ();
 DECAPx4_ASAP7_75t_R FILLER_251_174 ();
 FILLER_ASAP7_75t_R FILLER_251_184 ();
 DECAPx6_ASAP7_75t_R FILLER_251_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_215 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_249 ();
 DECAPx2_ASAP7_75t_R FILLER_251_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_303 ();
 DECAPx2_ASAP7_75t_R FILLER_251_310 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_316 ();
 DECAPx10_ASAP7_75t_R FILLER_251_349 ();
 FILLER_ASAP7_75t_R FILLER_251_371 ();
 DECAPx2_ASAP7_75t_R FILLER_251_379 ();
 FILLER_ASAP7_75t_R FILLER_251_385 ();
 DECAPx2_ASAP7_75t_R FILLER_251_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_419 ();
 DECAPx6_ASAP7_75t_R FILLER_251_426 ();
 DECAPx1_ASAP7_75t_R FILLER_251_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_444 ();
 DECAPx10_ASAP7_75t_R FILLER_251_448 ();
 DECAPx6_ASAP7_75t_R FILLER_251_470 ();
 DECAPx10_ASAP7_75t_R FILLER_251_487 ();
 DECAPx10_ASAP7_75t_R FILLER_251_509 ();
 FILLER_ASAP7_75t_R FILLER_251_531 ();
 DECAPx6_ASAP7_75t_R FILLER_251_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_550 ();
 DECAPx10_ASAP7_75t_R FILLER_251_563 ();
 DECAPx2_ASAP7_75t_R FILLER_251_585 ();
 DECAPx1_ASAP7_75t_R FILLER_251_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_609 ();
 DECAPx10_ASAP7_75t_R FILLER_251_620 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_251_642 ();
 DECAPx10_ASAP7_75t_R FILLER_251_661 ();
 DECAPx2_ASAP7_75t_R FILLER_251_683 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_689 ();
 DECAPx4_ASAP7_75t_R FILLER_251_699 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_786 ();
 FILLER_ASAP7_75t_R FILLER_251_810 ();
 DECAPx2_ASAP7_75t_R FILLER_251_815 ();
 FILLER_ASAP7_75t_R FILLER_251_821 ();
 DECAPx2_ASAP7_75t_R FILLER_251_826 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_843 ();
 DECAPx1_ASAP7_75t_R FILLER_251_854 ();
 DECAPx1_ASAP7_75t_R FILLER_251_869 ();
 FILLER_ASAP7_75t_R FILLER_251_879 ();
 DECAPx1_ASAP7_75t_R FILLER_251_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_251_933 ();
 DECAPx10_ASAP7_75t_R FILLER_252_2 ();
 DECAPx10_ASAP7_75t_R FILLER_252_24 ();
 DECAPx10_ASAP7_75t_R FILLER_252_46 ();
 DECAPx6_ASAP7_75t_R FILLER_252_68 ();
 DECAPx10_ASAP7_75t_R FILLER_252_91 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_113 ();
 DECAPx2_ASAP7_75t_R FILLER_252_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_132 ();
 DECAPx2_ASAP7_75t_R FILLER_252_165 ();
 FILLER_ASAP7_75t_R FILLER_252_171 ();
 FILLER_ASAP7_75t_R FILLER_252_182 ();
 FILLER_ASAP7_75t_R FILLER_252_206 ();
 DECAPx1_ASAP7_75t_R FILLER_252_211 ();
 DECAPx6_ASAP7_75t_R FILLER_252_261 ();
 DECAPx2_ASAP7_75t_R FILLER_252_275 ();
 DECAPx2_ASAP7_75t_R FILLER_252_302 ();
 DECAPx4_ASAP7_75t_R FILLER_252_340 ();
 FILLER_ASAP7_75t_R FILLER_252_350 ();
 DECAPx4_ASAP7_75t_R FILLER_252_358 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_368 ();
 DECAPx4_ASAP7_75t_R FILLER_252_393 ();
 DECAPx10_ASAP7_75t_R FILLER_252_415 ();
 DECAPx6_ASAP7_75t_R FILLER_252_437 ();
 DECAPx2_ASAP7_75t_R FILLER_252_454 ();
 FILLER_ASAP7_75t_R FILLER_252_460 ();
 DECAPx1_ASAP7_75t_R FILLER_252_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_472 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_476 ();
 DECAPx1_ASAP7_75t_R FILLER_252_506 ();
 DECAPx6_ASAP7_75t_R FILLER_252_524 ();
 DECAPx1_ASAP7_75t_R FILLER_252_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_542 ();
 DECAPx6_ASAP7_75t_R FILLER_252_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_563 ();
 DECAPx2_ASAP7_75t_R FILLER_252_584 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_600 ();
 DECAPx1_ASAP7_75t_R FILLER_252_640 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_668 ();
 DECAPx6_ASAP7_75t_R FILLER_252_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_699 ();
 DECAPx1_ASAP7_75t_R FILLER_252_706 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_717 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_770 ();
 DECAPx10_ASAP7_75t_R FILLER_252_783 ();
 DECAPx2_ASAP7_75t_R FILLER_252_805 ();
 FILLER_ASAP7_75t_R FILLER_252_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_252_827 ();
 DECAPx4_ASAP7_75t_R FILLER_252_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_864 ();
 DECAPx4_ASAP7_75t_R FILLER_252_870 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_252_880 ();
 DECAPx10_ASAP7_75t_R FILLER_253_2 ();
 DECAPx10_ASAP7_75t_R FILLER_253_24 ();
 DECAPx10_ASAP7_75t_R FILLER_253_46 ();
 DECAPx2_ASAP7_75t_R FILLER_253_68 ();
 DECAPx2_ASAP7_75t_R FILLER_253_103 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_135 ();
 DECAPx1_ASAP7_75t_R FILLER_253_150 ();
 DECAPx1_ASAP7_75t_R FILLER_253_157 ();
 DECAPx1_ASAP7_75t_R FILLER_253_193 ();
 DECAPx4_ASAP7_75t_R FILLER_253_219 ();
 FILLER_ASAP7_75t_R FILLER_253_229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_238 ();
 DECAPx4_ASAP7_75t_R FILLER_253_253 ();
 DECAPx4_ASAP7_75t_R FILLER_253_278 ();
 DECAPx6_ASAP7_75t_R FILLER_253_295 ();
 DECAPx1_ASAP7_75t_R FILLER_253_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_326 ();
 DECAPx4_ASAP7_75t_R FILLER_253_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_340 ();
 DECAPx10_ASAP7_75t_R FILLER_253_367 ();
 DECAPx2_ASAP7_75t_R FILLER_253_389 ();
 FILLER_ASAP7_75t_R FILLER_253_395 ();
 DECAPx4_ASAP7_75t_R FILLER_253_419 ();
 DECAPx2_ASAP7_75t_R FILLER_253_435 ();
 DECAPx6_ASAP7_75t_R FILLER_253_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_469 ();
 FILLER_ASAP7_75t_R FILLER_253_482 ();
 DECAPx1_ASAP7_75t_R FILLER_253_508 ();
 DECAPx2_ASAP7_75t_R FILLER_253_552 ();
 DECAPx6_ASAP7_75t_R FILLER_253_566 ();
 DECAPx2_ASAP7_75t_R FILLER_253_580 ();
 DECAPx4_ASAP7_75t_R FILLER_253_592 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_602 ();
 DECAPx1_ASAP7_75t_R FILLER_253_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_621 ();
 FILLER_ASAP7_75t_R FILLER_253_629 ();
 DECAPx6_ASAP7_75t_R FILLER_253_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_671 ();
 DECAPx2_ASAP7_75t_R FILLER_253_692 ();
 DECAPx4_ASAP7_75t_R FILLER_253_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_720 ();
 DECAPx10_ASAP7_75t_R FILLER_253_753 ();
 DECAPx2_ASAP7_75t_R FILLER_253_775 ();
 FILLER_ASAP7_75t_R FILLER_253_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_806 ();
 FILLER_ASAP7_75t_R FILLER_253_840 ();
 DECAPx4_ASAP7_75t_R FILLER_253_845 ();
 FILLER_ASAP7_75t_R FILLER_253_855 ();
 DECAPx6_ASAP7_75t_R FILLER_253_863 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_253_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_253_906 ();
 FILLER_ASAP7_75t_R FILLER_253_932 ();
 DECAPx10_ASAP7_75t_R FILLER_254_2 ();
 DECAPx10_ASAP7_75t_R FILLER_254_24 ();
 DECAPx10_ASAP7_75t_R FILLER_254_46 ();
 DECAPx2_ASAP7_75t_R FILLER_254_68 ();
 DECAPx6_ASAP7_75t_R FILLER_254_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_123 ();
 DECAPx6_ASAP7_75t_R FILLER_254_127 ();
 DECAPx2_ASAP7_75t_R FILLER_254_141 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_211 ();
 DECAPx4_ASAP7_75t_R FILLER_254_218 ();
 DECAPx1_ASAP7_75t_R FILLER_254_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_258 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_294 ();
 DECAPx10_ASAP7_75t_R FILLER_254_303 ();
 DECAPx6_ASAP7_75t_R FILLER_254_325 ();
 FILLER_ASAP7_75t_R FILLER_254_345 ();
 FILLER_ASAP7_75t_R FILLER_254_353 ();
 DECAPx10_ASAP7_75t_R FILLER_254_358 ();
 DECAPx6_ASAP7_75t_R FILLER_254_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_394 ();
 DECAPx4_ASAP7_75t_R FILLER_254_409 ();
 FILLER_ASAP7_75t_R FILLER_254_419 ();
 DECAPx2_ASAP7_75t_R FILLER_254_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_451 ();
 DECAPx2_ASAP7_75t_R FILLER_254_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_464 ();
 DECAPx1_ASAP7_75t_R FILLER_254_497 ();
 DECAPx2_ASAP7_75t_R FILLER_254_527 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_533 ();
 FILLER_ASAP7_75t_R FILLER_254_570 ();
 DECAPx6_ASAP7_75t_R FILLER_254_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_612 ();
 DECAPx10_ASAP7_75t_R FILLER_254_632 ();
 DECAPx4_ASAP7_75t_R FILLER_254_654 ();
 DECAPx2_ASAP7_75t_R FILLER_254_676 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_682 ();
 DECAPx2_ASAP7_75t_R FILLER_254_695 ();
 DECAPx6_ASAP7_75t_R FILLER_254_707 ();
 DECAPx2_ASAP7_75t_R FILLER_254_721 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_732 ();
 DECAPx10_ASAP7_75t_R FILLER_254_736 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_758 ();
 DECAPx2_ASAP7_75t_R FILLER_254_770 ();
 FILLER_ASAP7_75t_R FILLER_254_776 ();
 DECAPx1_ASAP7_75t_R FILLER_254_782 ();
 DECAPx2_ASAP7_75t_R FILLER_254_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_812 ();
 DECAPx1_ASAP7_75t_R FILLER_254_819 ();
 DECAPx6_ASAP7_75t_R FILLER_254_829 ();
 DECAPx1_ASAP7_75t_R FILLER_254_843 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_847 ();
 FILLER_ASAP7_75t_R FILLER_254_855 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_254_898 ();
 FILLER_ASAP7_75t_R FILLER_254_916 ();
 FILLERxp5_ASAP7_75t_R FILLER_254_933 ();
 DECAPx10_ASAP7_75t_R FILLER_255_2 ();
 DECAPx10_ASAP7_75t_R FILLER_255_24 ();
 DECAPx10_ASAP7_75t_R FILLER_255_46 ();
 DECAPx4_ASAP7_75t_R FILLER_255_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_85 ();
 DECAPx10_ASAP7_75t_R FILLER_255_116 ();
 DECAPx6_ASAP7_75t_R FILLER_255_138 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_152 ();
 DECAPx2_ASAP7_75t_R FILLER_255_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_189 ();
 DECAPx6_ASAP7_75t_R FILLER_255_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_238 ();
 DECAPx6_ASAP7_75t_R FILLER_255_248 ();
 DECAPx2_ASAP7_75t_R FILLER_255_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_311 ();
 DECAPx4_ASAP7_75t_R FILLER_255_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_331 ();
 DECAPx6_ASAP7_75t_R FILLER_255_372 ();
 DECAPx2_ASAP7_75t_R FILLER_255_386 ();
 DECAPx2_ASAP7_75t_R FILLER_255_418 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_424 ();
 DECAPx2_ASAP7_75t_R FILLER_255_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_439 ();
 FILLER_ASAP7_75t_R FILLER_255_443 ();
 FILLER_ASAP7_75t_R FILLER_255_448 ();
 DECAPx10_ASAP7_75t_R FILLER_255_467 ();
 DECAPx10_ASAP7_75t_R FILLER_255_489 ();
 DECAPx1_ASAP7_75t_R FILLER_255_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_526 ();
 FILLER_ASAP7_75t_R FILLER_255_568 ();
 DECAPx10_ASAP7_75t_R FILLER_255_593 ();
 DECAPx10_ASAP7_75t_R FILLER_255_615 ();
 DECAPx10_ASAP7_75t_R FILLER_255_637 ();
 DECAPx2_ASAP7_75t_R FILLER_255_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_665 ();
 DECAPx6_ASAP7_75t_R FILLER_255_681 ();
 DECAPx1_ASAP7_75t_R FILLER_255_695 ();
 DECAPx1_ASAP7_75t_R FILLER_255_705 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_709 ();
 DECAPx10_ASAP7_75t_R FILLER_255_716 ();
 DECAPx6_ASAP7_75t_R FILLER_255_738 ();
 DECAPx1_ASAP7_75t_R FILLER_255_752 ();
 DECAPx10_ASAP7_75t_R FILLER_255_784 ();
 DECAPx4_ASAP7_75t_R FILLER_255_806 ();
 DECAPx10_ASAP7_75t_R FILLER_255_822 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_255_844 ();
 DECAPx4_ASAP7_75t_R FILLER_255_858 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_255_933 ();
 DECAPx10_ASAP7_75t_R FILLER_256_2 ();
 DECAPx10_ASAP7_75t_R FILLER_256_24 ();
 DECAPx10_ASAP7_75t_R FILLER_256_46 ();
 DECAPx10_ASAP7_75t_R FILLER_256_68 ();
 DECAPx2_ASAP7_75t_R FILLER_256_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_96 ();
 DECAPx6_ASAP7_75t_R FILLER_256_105 ();
 DECAPx1_ASAP7_75t_R FILLER_256_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_132 ();
 DECAPx10_ASAP7_75t_R FILLER_256_136 ();
 DECAPx10_ASAP7_75t_R FILLER_256_158 ();
 DECAPx10_ASAP7_75t_R FILLER_256_180 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_202 ();
 DECAPx1_ASAP7_75t_R FILLER_256_209 ();
 DECAPx10_ASAP7_75t_R FILLER_256_216 ();
 DECAPx4_ASAP7_75t_R FILLER_256_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_248 ();
 DECAPx1_ASAP7_75t_R FILLER_256_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_259 ();
 DECAPx6_ASAP7_75t_R FILLER_256_263 ();
 DECAPx1_ASAP7_75t_R FILLER_256_277 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_301 ();
 FILLER_ASAP7_75t_R FILLER_256_334 ();
 DECAPx1_ASAP7_75t_R FILLER_256_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_346 ();
 DECAPx2_ASAP7_75t_R FILLER_256_350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_356 ();
 DECAPx1_ASAP7_75t_R FILLER_256_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_384 ();
 DECAPx6_ASAP7_75t_R FILLER_256_393 ();
 DECAPx1_ASAP7_75t_R FILLER_256_410 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_414 ();
 DECAPx2_ASAP7_75t_R FILLER_256_425 ();
 DECAPx6_ASAP7_75t_R FILLER_256_434 ();
 DECAPx1_ASAP7_75t_R FILLER_256_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_452 ();
 DECAPx2_ASAP7_75t_R FILLER_256_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_467 ();
 DECAPx10_ASAP7_75t_R FILLER_256_477 ();
 DECAPx10_ASAP7_75t_R FILLER_256_499 ();
 DECAPx2_ASAP7_75t_R FILLER_256_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_527 ();
 DECAPx6_ASAP7_75t_R FILLER_256_534 ();
 FILLER_ASAP7_75t_R FILLER_256_548 ();
 DECAPx1_ASAP7_75t_R FILLER_256_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_557 ();
 DECAPx4_ASAP7_75t_R FILLER_256_561 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_571 ();
 DECAPx10_ASAP7_75t_R FILLER_256_608 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_630 ();
 DECAPx2_ASAP7_75t_R FILLER_256_641 ();
 FILLER_ASAP7_75t_R FILLER_256_647 ();
 DECAPx4_ASAP7_75t_R FILLER_256_657 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_667 ();
 DECAPx2_ASAP7_75t_R FILLER_256_674 ();
 FILLER_ASAP7_75t_R FILLER_256_680 ();
 DECAPx4_ASAP7_75t_R FILLER_256_689 ();
 DECAPx1_ASAP7_75t_R FILLER_256_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_711 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_722 ();
 DECAPx1_ASAP7_75t_R FILLER_256_732 ();
 DECAPx2_ASAP7_75t_R FILLER_256_742 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_748 ();
 DECAPx6_ASAP7_75t_R FILLER_256_756 ();
 DECAPx1_ASAP7_75t_R FILLER_256_770 ();
 FILLERxp5_ASAP7_75t_R FILLER_256_794 ();
 DECAPx10_ASAP7_75t_R FILLER_256_803 ();
 DECAPx4_ASAP7_75t_R FILLER_256_825 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_256_835 ();
 DECAPx10_ASAP7_75t_R FILLER_256_844 ();
 DECAPx2_ASAP7_75t_R FILLER_256_866 ();
 FILLER_ASAP7_75t_R FILLER_256_872 ();
 DECAPx10_ASAP7_75t_R FILLER_257_2 ();
 DECAPx10_ASAP7_75t_R FILLER_257_24 ();
 DECAPx10_ASAP7_75t_R FILLER_257_46 ();
 DECAPx10_ASAP7_75t_R FILLER_257_68 ();
 DECAPx6_ASAP7_75t_R FILLER_257_90 ();
 DECAPx2_ASAP7_75t_R FILLER_257_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_110 ();
 DECAPx1_ASAP7_75t_R FILLER_257_137 ();
 DECAPx10_ASAP7_75t_R FILLER_257_147 ();
 DECAPx6_ASAP7_75t_R FILLER_257_169 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_192 ();
 DECAPx4_ASAP7_75t_R FILLER_257_198 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_208 ();
 DECAPx1_ASAP7_75t_R FILLER_257_235 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_239 ();
 DECAPx6_ASAP7_75t_R FILLER_257_266 ();
 DECAPx2_ASAP7_75t_R FILLER_257_280 ();
 DECAPx2_ASAP7_75t_R FILLER_257_333 ();
 DECAPx4_ASAP7_75t_R FILLER_257_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_359 ();
 DECAPx2_ASAP7_75t_R FILLER_257_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_369 ();
 DECAPx6_ASAP7_75t_R FILLER_257_402 ();
 DECAPx2_ASAP7_75t_R FILLER_257_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_422 ();
 DECAPx2_ASAP7_75t_R FILLER_257_432 ();
 FILLER_ASAP7_75t_R FILLER_257_438 ();
 DECAPx10_ASAP7_75t_R FILLER_257_449 ();
 DECAPx6_ASAP7_75t_R FILLER_257_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_485 ();
 DECAPx2_ASAP7_75t_R FILLER_257_495 ();
 DECAPx6_ASAP7_75t_R FILLER_257_511 ();
 DECAPx2_ASAP7_75t_R FILLER_257_525 ();
 DECAPx10_ASAP7_75t_R FILLER_257_537 ();
 DECAPx10_ASAP7_75t_R FILLER_257_559 ();
 DECAPx2_ASAP7_75t_R FILLER_257_581 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_587 ();
 DECAPx2_ASAP7_75t_R FILLER_257_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_597 ();
 DECAPx2_ASAP7_75t_R FILLER_257_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_635 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_648 ();
 DECAPx10_ASAP7_75t_R FILLER_257_663 ();
 DECAPx10_ASAP7_75t_R FILLER_257_685 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_707 ();
 DECAPx1_ASAP7_75t_R FILLER_257_716 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_720 ();
 DECAPx2_ASAP7_75t_R FILLER_257_759 ();
 FILLER_ASAP7_75t_R FILLER_257_765 ();
 DECAPx1_ASAP7_75t_R FILLER_257_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_808 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_815 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_257_824 ();
 DECAPx1_ASAP7_75t_R FILLER_257_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_848 ();
 DECAPx4_ASAP7_75t_R FILLER_257_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_877 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_897 ();
 FILLER_ASAP7_75t_R FILLER_257_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_257_927 ();
 DECAPx10_ASAP7_75t_R FILLER_258_2 ();
 DECAPx10_ASAP7_75t_R FILLER_258_24 ();
 DECAPx10_ASAP7_75t_R FILLER_258_46 ();
 DECAPx4_ASAP7_75t_R FILLER_258_68 ();
 FILLER_ASAP7_75t_R FILLER_258_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_86 ();
 DECAPx4_ASAP7_75t_R FILLER_258_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_103 ();
 DECAPx2_ASAP7_75t_R FILLER_258_110 ();
 FILLER_ASAP7_75t_R FILLER_258_116 ();
 DECAPx1_ASAP7_75t_R FILLER_258_124 ();
 DECAPx2_ASAP7_75t_R FILLER_258_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_172 ();
 DECAPx4_ASAP7_75t_R FILLER_258_205 ();
 FILLER_ASAP7_75t_R FILLER_258_215 ();
 FILLER_ASAP7_75t_R FILLER_258_243 ();
 DECAPx1_ASAP7_75t_R FILLER_258_251 ();
 DECAPx4_ASAP7_75t_R FILLER_258_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_268 ();
 DECAPx6_ASAP7_75t_R FILLER_258_275 ();
 DECAPx1_ASAP7_75t_R FILLER_258_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_293 ();
 DECAPx10_ASAP7_75t_R FILLER_258_300 ();
 DECAPx6_ASAP7_75t_R FILLER_258_328 ();
 DECAPx1_ASAP7_75t_R FILLER_258_342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_372 ();
 FILLER_ASAP7_75t_R FILLER_258_381 ();
 DECAPx4_ASAP7_75t_R FILLER_258_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_412 ();
 DECAPx2_ASAP7_75t_R FILLER_258_416 ();
 DECAPx1_ASAP7_75t_R FILLER_258_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_429 ();
 DECAPx6_ASAP7_75t_R FILLER_258_433 ();
 DECAPx4_ASAP7_75t_R FILLER_258_450 ();
 FILLER_ASAP7_75t_R FILLER_258_460 ();
 DECAPx2_ASAP7_75t_R FILLER_258_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_258_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_514 ();
 DECAPx6_ASAP7_75t_R FILLER_258_523 ();
 DECAPx1_ASAP7_75t_R FILLER_258_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_541 ();
 DECAPx4_ASAP7_75t_R FILLER_258_552 ();
 DECAPx4_ASAP7_75t_R FILLER_258_594 ();
 FILLER_ASAP7_75t_R FILLER_258_604 ();
 DECAPx2_ASAP7_75t_R FILLER_258_612 ();
 DECAPx10_ASAP7_75t_R FILLER_258_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_650 ();
 DECAPx2_ASAP7_75t_R FILLER_258_673 ();
 DECAPx1_ASAP7_75t_R FILLER_258_694 ();
 DECAPx10_ASAP7_75t_R FILLER_258_704 ();
 FILLER_ASAP7_75t_R FILLER_258_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_735 ();
 FILLER_ASAP7_75t_R FILLER_258_745 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_783 ();
 FILLER_ASAP7_75t_R FILLER_258_825 ();
 DECAPx4_ASAP7_75t_R FILLER_258_879 ();
 FILLER_ASAP7_75t_R FILLER_258_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_258_903 ();
 DECAPx10_ASAP7_75t_R FILLER_259_2 ();
 DECAPx10_ASAP7_75t_R FILLER_259_24 ();
 DECAPx10_ASAP7_75t_R FILLER_259_46 ();
 DECAPx1_ASAP7_75t_R FILLER_259_68 ();
 DECAPx1_ASAP7_75t_R FILLER_259_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_102 ();
 FILLER_ASAP7_75t_R FILLER_259_145 ();
 DECAPx1_ASAP7_75t_R FILLER_259_150 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_161 ();
 FILLER_ASAP7_75t_R FILLER_259_207 ();
 DECAPx10_ASAP7_75t_R FILLER_259_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_261 ();
 DECAPx6_ASAP7_75t_R FILLER_259_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_324 ();
 DECAPx4_ASAP7_75t_R FILLER_259_337 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_347 ();
 DECAPx10_ASAP7_75t_R FILLER_259_356 ();
 DECAPx2_ASAP7_75t_R FILLER_259_378 ();
 FILLER_ASAP7_75t_R FILLER_259_384 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_441 ();
 DECAPx10_ASAP7_75t_R FILLER_259_458 ();
 DECAPx1_ASAP7_75t_R FILLER_259_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_484 ();
 DECAPx2_ASAP7_75t_R FILLER_259_496 ();
 DECAPx2_ASAP7_75t_R FILLER_259_505 ();
 DECAPx2_ASAP7_75t_R FILLER_259_537 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_543 ();
 DECAPx2_ASAP7_75t_R FILLER_259_556 ();
 FILLER_ASAP7_75t_R FILLER_259_562 ();
 DECAPx10_ASAP7_75t_R FILLER_259_570 ();
 DECAPx1_ASAP7_75t_R FILLER_259_592 ();
 FILLER_ASAP7_75t_R FILLER_259_602 ();
 DECAPx10_ASAP7_75t_R FILLER_259_612 ();
 DECAPx4_ASAP7_75t_R FILLER_259_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_644 ();
 DECAPx2_ASAP7_75t_R FILLER_259_651 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_669 ();
 DECAPx1_ASAP7_75t_R FILLER_259_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_684 ();
 FILLER_ASAP7_75t_R FILLER_259_691 ();
 DECAPx6_ASAP7_75t_R FILLER_259_705 ();
 DECAPx1_ASAP7_75t_R FILLER_259_719 ();
 DECAPx1_ASAP7_75t_R FILLER_259_749 ();
 DECAPx2_ASAP7_75t_R FILLER_259_761 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_767 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_259_783 ();
 DECAPx2_ASAP7_75t_R FILLER_259_848 ();
 FILLER_ASAP7_75t_R FILLER_259_854 ();
 DECAPx10_ASAP7_75t_R FILLER_259_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_889 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_919 ();
 FILLERxp5_ASAP7_75t_R FILLER_259_933 ();
 DECAPx10_ASAP7_75t_R FILLER_260_2 ();
 DECAPx10_ASAP7_75t_R FILLER_260_24 ();
 DECAPx6_ASAP7_75t_R FILLER_260_46 ();
 DECAPx2_ASAP7_75t_R FILLER_260_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_66 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_129 ();
 DECAPx4_ASAP7_75t_R FILLER_260_136 ();
 FILLER_ASAP7_75t_R FILLER_260_146 ();
 DECAPx6_ASAP7_75t_R FILLER_260_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_182 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_223 ();
 DECAPx6_ASAP7_75t_R FILLER_260_227 ();
 DECAPx1_ASAP7_75t_R FILLER_260_241 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_245 ();
 DECAPx1_ASAP7_75t_R FILLER_260_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_256 ();
 DECAPx1_ASAP7_75t_R FILLER_260_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_288 ();
 FILLER_ASAP7_75t_R FILLER_260_336 ();
 DECAPx10_ASAP7_75t_R FILLER_260_346 ();
 DECAPx10_ASAP7_75t_R FILLER_260_368 ();
 DECAPx6_ASAP7_75t_R FILLER_260_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_404 ();
 DECAPx10_ASAP7_75t_R FILLER_260_411 ();
 DECAPx2_ASAP7_75t_R FILLER_260_445 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_451 ();
 FILLER_ASAP7_75t_R FILLER_260_457 ();
 DECAPx4_ASAP7_75t_R FILLER_260_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_491 ();
 DECAPx2_ASAP7_75t_R FILLER_260_498 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_504 ();
 DECAPx2_ASAP7_75t_R FILLER_260_511 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_260_517 ();
 DECAPx1_ASAP7_75t_R FILLER_260_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_565 ();
 FILLER_ASAP7_75t_R FILLER_260_574 ();
 DECAPx6_ASAP7_75t_R FILLER_260_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_597 ();
 DECAPx1_ASAP7_75t_R FILLER_260_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_609 ();
 DECAPx4_ASAP7_75t_R FILLER_260_616 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_645 ();
 DECAPx4_ASAP7_75t_R FILLER_260_655 ();
 FILLER_ASAP7_75t_R FILLER_260_665 ();
 DECAPx10_ASAP7_75t_R FILLER_260_673 ();
 DECAPx4_ASAP7_75t_R FILLER_260_701 ();
 DECAPx6_ASAP7_75t_R FILLER_260_723 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_740 ();
 DECAPx10_ASAP7_75t_R FILLER_260_746 ();
 DECAPx10_ASAP7_75t_R FILLER_260_768 ();
 DECAPx2_ASAP7_75t_R FILLER_260_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_796 ();
 DECAPx2_ASAP7_75t_R FILLER_260_800 ();
 DECAPx10_ASAP7_75t_R FILLER_260_831 ();
 DECAPx10_ASAP7_75t_R FILLER_260_853 ();
 DECAPx1_ASAP7_75t_R FILLER_260_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_260_933 ();
 DECAPx10_ASAP7_75t_R FILLER_261_2 ();
 DECAPx10_ASAP7_75t_R FILLER_261_24 ();
 DECAPx10_ASAP7_75t_R FILLER_261_46 ();
 DECAPx1_ASAP7_75t_R FILLER_261_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_72 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_85 ();
 DECAPx6_ASAP7_75t_R FILLER_261_127 ();
 DECAPx1_ASAP7_75t_R FILLER_261_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_145 ();
 DECAPx10_ASAP7_75t_R FILLER_261_152 ();
 DECAPx4_ASAP7_75t_R FILLER_261_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_184 ();
 DECAPx2_ASAP7_75t_R FILLER_261_229 ();
 FILLER_ASAP7_75t_R FILLER_261_235 ();
 DECAPx4_ASAP7_75t_R FILLER_261_271 ();
 DECAPx1_ASAP7_75t_R FILLER_261_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_361 ();
 DECAPx1_ASAP7_75t_R FILLER_261_396 ();
 DECAPx6_ASAP7_75t_R FILLER_261_406 ();
 FILLER_ASAP7_75t_R FILLER_261_420 ();
 DECAPx6_ASAP7_75t_R FILLER_261_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_439 ();
 DECAPx2_ASAP7_75t_R FILLER_261_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_449 ();
 DECAPx1_ASAP7_75t_R FILLER_261_490 ();
 DECAPx2_ASAP7_75t_R FILLER_261_501 ();
 DECAPx6_ASAP7_75t_R FILLER_261_514 ();
 FILLER_ASAP7_75t_R FILLER_261_528 ();
 DECAPx10_ASAP7_75t_R FILLER_261_538 ();
 DECAPx6_ASAP7_75t_R FILLER_261_560 ();
 FILLER_ASAP7_75t_R FILLER_261_574 ();
 DECAPx1_ASAP7_75t_R FILLER_261_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_587 ();
 DECAPx6_ASAP7_75t_R FILLER_261_596 ();
 DECAPx2_ASAP7_75t_R FILLER_261_610 ();
 DECAPx2_ASAP7_75t_R FILLER_261_623 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_629 ();
 DECAPx10_ASAP7_75t_R FILLER_261_652 ();
 DECAPx2_ASAP7_75t_R FILLER_261_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_680 ();
 DECAPx6_ASAP7_75t_R FILLER_261_687 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_701 ();
 DECAPx10_ASAP7_75t_R FILLER_261_726 ();
 DECAPx1_ASAP7_75t_R FILLER_261_748 ();
 DECAPx10_ASAP7_75t_R FILLER_261_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_777 ();
 DECAPx10_ASAP7_75t_R FILLER_261_785 ();
 DECAPx10_ASAP7_75t_R FILLER_261_807 ();
 DECAPx4_ASAP7_75t_R FILLER_261_829 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_261_839 ();
 DECAPx1_ASAP7_75t_R FILLER_261_849 ();
 DECAPx1_ASAP7_75t_R FILLER_261_859 ();
 DECAPx1_ASAP7_75t_R FILLER_261_866 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_870 ();
 DECAPx1_ASAP7_75t_R FILLER_261_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_891 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_904 ();
 FILLER_ASAP7_75t_R FILLER_261_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_261_933 ();
 DECAPx10_ASAP7_75t_R FILLER_262_2 ();
 DECAPx10_ASAP7_75t_R FILLER_262_24 ();
 DECAPx10_ASAP7_75t_R FILLER_262_46 ();
 DECAPx10_ASAP7_75t_R FILLER_262_68 ();
 DECAPx10_ASAP7_75t_R FILLER_262_90 ();
 DECAPx2_ASAP7_75t_R FILLER_262_118 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_124 ();
 DECAPx2_ASAP7_75t_R FILLER_262_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_145 ();
 DECAPx4_ASAP7_75t_R FILLER_262_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_182 ();
 DECAPx4_ASAP7_75t_R FILLER_262_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_254 ();
 DECAPx2_ASAP7_75t_R FILLER_262_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_273 ();
 FILLER_ASAP7_75t_R FILLER_262_300 ();
 DECAPx1_ASAP7_75t_R FILLER_262_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_340 ();
 DECAPx1_ASAP7_75t_R FILLER_262_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_351 ();
 DECAPx1_ASAP7_75t_R FILLER_262_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_390 ();
 DECAPx6_ASAP7_75t_R FILLER_262_417 ();
 FILLER_ASAP7_75t_R FILLER_262_431 ();
 DECAPx4_ASAP7_75t_R FILLER_262_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_446 ();
 DECAPx2_ASAP7_75t_R FILLER_262_456 ();
 DECAPx2_ASAP7_75t_R FILLER_262_464 ();
 FILLER_ASAP7_75t_R FILLER_262_470 ();
 DECAPx4_ASAP7_75t_R FILLER_262_489 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_499 ();
 DECAPx1_ASAP7_75t_R FILLER_262_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_514 ();
 DECAPx10_ASAP7_75t_R FILLER_262_518 ();
 DECAPx6_ASAP7_75t_R FILLER_262_540 ();
 DECAPx1_ASAP7_75t_R FILLER_262_554 ();
 DECAPx6_ASAP7_75t_R FILLER_262_564 ();
 DECAPx2_ASAP7_75t_R FILLER_262_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_584 ();
 DECAPx2_ASAP7_75t_R FILLER_262_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_599 ();
 DECAPx1_ASAP7_75t_R FILLER_262_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_624 ();
 DECAPx10_ASAP7_75t_R FILLER_262_633 ();
 DECAPx10_ASAP7_75t_R FILLER_262_655 ();
 DECAPx6_ASAP7_75t_R FILLER_262_677 ();
 DECAPx2_ASAP7_75t_R FILLER_262_691 ();
 DECAPx2_ASAP7_75t_R FILLER_262_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_732 ();
 FILLER_ASAP7_75t_R FILLER_262_752 ();
 FILLER_ASAP7_75t_R FILLER_262_775 ();
 DECAPx10_ASAP7_75t_R FILLER_262_788 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_262_810 ();
 DECAPx6_ASAP7_75t_R FILLER_262_818 ();
 DECAPx2_ASAP7_75t_R FILLER_262_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_262_838 ();
 FILLER_ASAP7_75t_R FILLER_262_847 ();
 DECAPx10_ASAP7_75t_R FILLER_263_2 ();
 DECAPx10_ASAP7_75t_R FILLER_263_24 ();
 DECAPx10_ASAP7_75t_R FILLER_263_46 ();
 DECAPx10_ASAP7_75t_R FILLER_263_68 ();
 DECAPx6_ASAP7_75t_R FILLER_263_90 ();
 DECAPx1_ASAP7_75t_R FILLER_263_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_108 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_115 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_124 ();
 FILLER_ASAP7_75t_R FILLER_263_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_229 ();
 DECAPx4_ASAP7_75t_R FILLER_263_244 ();
 DECAPx6_ASAP7_75t_R FILLER_263_260 ();
 DECAPx1_ASAP7_75t_R FILLER_263_274 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_284 ();
 FILLER_ASAP7_75t_R FILLER_263_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_299 ();
 DECAPx1_ASAP7_75t_R FILLER_263_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_310 ();
 DECAPx1_ASAP7_75t_R FILLER_263_317 ();
 FILLER_ASAP7_75t_R FILLER_263_324 ();
 DECAPx4_ASAP7_75t_R FILLER_263_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_342 ();
 DECAPx2_ASAP7_75t_R FILLER_263_349 ();
 FILLER_ASAP7_75t_R FILLER_263_355 ();
 DECAPx1_ASAP7_75t_R FILLER_263_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_373 ();
 DECAPx6_ASAP7_75t_R FILLER_263_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_394 ();
 DECAPx1_ASAP7_75t_R FILLER_263_401 ();
 DECAPx6_ASAP7_75t_R FILLER_263_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_425 ();
 DECAPx6_ASAP7_75t_R FILLER_263_435 ();
 DECAPx1_ASAP7_75t_R FILLER_263_449 ();
 DECAPx4_ASAP7_75t_R FILLER_263_459 ();
 FILLER_ASAP7_75t_R FILLER_263_469 ();
 DECAPx2_ASAP7_75t_R FILLER_263_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_498 ();
 FILLER_ASAP7_75t_R FILLER_263_533 ();
 DECAPx4_ASAP7_75t_R FILLER_263_549 ();
 FILLER_ASAP7_75t_R FILLER_263_559 ();
 DECAPx4_ASAP7_75t_R FILLER_263_579 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_589 ();
 DECAPx6_ASAP7_75t_R FILLER_263_598 ();
 DECAPx2_ASAP7_75t_R FILLER_263_612 ();
 DECAPx4_ASAP7_75t_R FILLER_263_630 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_646 ();
 DECAPx2_ASAP7_75t_R FILLER_263_653 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_659 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_674 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_690 ();
 DECAPx4_ASAP7_75t_R FILLER_263_713 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_776 ();
 DECAPx2_ASAP7_75t_R FILLER_263_791 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_797 ();
 DECAPx6_ASAP7_75t_R FILLER_263_803 ();
 DECAPx1_ASAP7_75t_R FILLER_263_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_821 ();
 DECAPx6_ASAP7_75t_R FILLER_263_828 ();
 DECAPx1_ASAP7_75t_R FILLER_263_842 ();
 DECAPx2_ASAP7_75t_R FILLER_263_849 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_855 ();
 DECAPx2_ASAP7_75t_R FILLER_263_861 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_263_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_917 ();
 FILLERxp5_ASAP7_75t_R FILLER_263_924 ();
 FILLER_ASAP7_75t_R FILLER_263_932 ();
 DECAPx10_ASAP7_75t_R FILLER_264_2 ();
 DECAPx10_ASAP7_75t_R FILLER_264_24 ();
 DECAPx10_ASAP7_75t_R FILLER_264_46 ();
 DECAPx2_ASAP7_75t_R FILLER_264_97 ();
 FILLER_ASAP7_75t_R FILLER_264_103 ();
 DECAPx2_ASAP7_75t_R FILLER_264_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_140 ();
 DECAPx6_ASAP7_75t_R FILLER_264_152 ();
 FILLER_ASAP7_75t_R FILLER_264_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_177 ();
 DECAPx1_ASAP7_75t_R FILLER_264_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_217 ();
 DECAPx2_ASAP7_75t_R FILLER_264_224 ();
 FILLER_ASAP7_75t_R FILLER_264_230 ();
 DECAPx10_ASAP7_75t_R FILLER_264_264 ();
 FILLER_ASAP7_75t_R FILLER_264_286 ();
 DECAPx10_ASAP7_75t_R FILLER_264_291 ();
 DECAPx6_ASAP7_75t_R FILLER_264_313 ();
 DECAPx2_ASAP7_75t_R FILLER_264_327 ();
 DECAPx6_ASAP7_75t_R FILLER_264_359 ();
 DECAPx1_ASAP7_75t_R FILLER_264_373 ();
 DECAPx10_ASAP7_75t_R FILLER_264_391 ();
 DECAPx2_ASAP7_75t_R FILLER_264_413 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_419 ();
 DECAPx1_ASAP7_75t_R FILLER_264_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_432 ();
 DECAPx6_ASAP7_75t_R FILLER_264_442 ();
 DECAPx2_ASAP7_75t_R FILLER_264_456 ();
 DECAPx2_ASAP7_75t_R FILLER_264_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_470 ();
 DECAPx1_ASAP7_75t_R FILLER_264_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_487 ();
 DECAPx4_ASAP7_75t_R FILLER_264_510 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_520 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_551 ();
 DECAPx2_ASAP7_75t_R FILLER_264_563 ();
 DECAPx1_ASAP7_75t_R FILLER_264_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_580 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_587 ();
 DECAPx6_ASAP7_75t_R FILLER_264_604 ();
 DECAPx2_ASAP7_75t_R FILLER_264_630 ();
 FILLER_ASAP7_75t_R FILLER_264_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_690 ();
 DECAPx10_ASAP7_75t_R FILLER_264_705 ();
 DECAPx4_ASAP7_75t_R FILLER_264_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_737 ();
 DECAPx6_ASAP7_75t_R FILLER_264_771 ();
 DECAPx2_ASAP7_75t_R FILLER_264_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_264_791 ();
 DECAPx2_ASAP7_75t_R FILLER_264_799 ();
 FILLER_ASAP7_75t_R FILLER_264_805 ();
 DECAPx2_ASAP7_75t_R FILLER_264_813 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_264_819 ();
 DECAPx10_ASAP7_75t_R FILLER_264_858 ();
 DECAPx4_ASAP7_75t_R FILLER_264_880 ();
 FILLER_ASAP7_75t_R FILLER_264_890 ();
 FILLER_ASAP7_75t_R FILLER_264_932 ();
 DECAPx10_ASAP7_75t_R FILLER_265_2 ();
 DECAPx10_ASAP7_75t_R FILLER_265_24 ();
 DECAPx10_ASAP7_75t_R FILLER_265_46 ();
 DECAPx4_ASAP7_75t_R FILLER_265_68 ();
 FILLER_ASAP7_75t_R FILLER_265_84 ();
 DECAPx6_ASAP7_75t_R FILLER_265_95 ();
 DECAPx1_ASAP7_75t_R FILLER_265_109 ();
 DECAPx10_ASAP7_75t_R FILLER_265_127 ();
 DECAPx10_ASAP7_75t_R FILLER_265_149 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_171 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_180 ();
 DECAPx10_ASAP7_75t_R FILLER_265_198 ();
 DECAPx4_ASAP7_75t_R FILLER_265_220 ();
 FILLER_ASAP7_75t_R FILLER_265_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_238 ();
 DECAPx6_ASAP7_75t_R FILLER_265_277 ();
 DECAPx1_ASAP7_75t_R FILLER_265_291 ();
 FILLER_ASAP7_75t_R FILLER_265_301 ();
 DECAPx10_ASAP7_75t_R FILLER_265_309 ();
 DECAPx2_ASAP7_75t_R FILLER_265_331 ();
 FILLER_ASAP7_75t_R FILLER_265_337 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_345 ();
 DECAPx4_ASAP7_75t_R FILLER_265_351 ();
 FILLER_ASAP7_75t_R FILLER_265_361 ();
 DECAPx6_ASAP7_75t_R FILLER_265_369 ();
 DECAPx1_ASAP7_75t_R FILLER_265_383 ();
 DECAPx6_ASAP7_75t_R FILLER_265_394 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_408 ();
 DECAPx1_ASAP7_75t_R FILLER_265_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_435 ();
 DECAPx2_ASAP7_75t_R FILLER_265_443 ();
 DECAPx10_ASAP7_75t_R FILLER_265_459 ();
 DECAPx2_ASAP7_75t_R FILLER_265_481 ();
 FILLER_ASAP7_75t_R FILLER_265_487 ();
 DECAPx10_ASAP7_75t_R FILLER_265_499 ();
 FILLER_ASAP7_75t_R FILLER_265_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_533 ();
 DECAPx4_ASAP7_75t_R FILLER_265_562 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_572 ();
 DECAPx1_ASAP7_75t_R FILLER_265_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_605 ();
 DECAPx10_ASAP7_75t_R FILLER_265_613 ();
 DECAPx2_ASAP7_75t_R FILLER_265_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_649 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_656 ();
 FILLER_ASAP7_75t_R FILLER_265_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_265_698 ();
 DECAPx10_ASAP7_75t_R FILLER_265_713 ();
 DECAPx2_ASAP7_75t_R FILLER_265_735 ();
 FILLER_ASAP7_75t_R FILLER_265_741 ();
 DECAPx6_ASAP7_75t_R FILLER_265_746 ();
 DECAPx10_ASAP7_75t_R FILLER_265_763 ();
 DECAPx1_ASAP7_75t_R FILLER_265_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_834 ();
 DECAPx10_ASAP7_75t_R FILLER_265_843 ();
 DECAPx10_ASAP7_75t_R FILLER_265_865 ();
 DECAPx2_ASAP7_75t_R FILLER_265_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_265_893 ();
 FILLER_ASAP7_75t_R FILLER_265_923 ();
 FILLER_ASAP7_75t_R FILLER_265_927 ();
 DECAPx10_ASAP7_75t_R FILLER_266_2 ();
 DECAPx10_ASAP7_75t_R FILLER_266_24 ();
 DECAPx10_ASAP7_75t_R FILLER_266_46 ();
 DECAPx4_ASAP7_75t_R FILLER_266_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_78 ();
 DECAPx10_ASAP7_75t_R FILLER_266_85 ();
 DECAPx10_ASAP7_75t_R FILLER_266_107 ();
 DECAPx10_ASAP7_75t_R FILLER_266_129 ();
 DECAPx4_ASAP7_75t_R FILLER_266_151 ();
 DECAPx2_ASAP7_75t_R FILLER_266_169 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_181 ();
 DECAPx6_ASAP7_75t_R FILLER_266_191 ();
 DECAPx2_ASAP7_75t_R FILLER_266_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_217 ();
 DECAPx10_ASAP7_75t_R FILLER_266_221 ();
 FILLER_ASAP7_75t_R FILLER_266_249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_289 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_322 ();
 DECAPx6_ASAP7_75t_R FILLER_266_331 ();
 DECAPx2_ASAP7_75t_R FILLER_266_345 ();
 DECAPx6_ASAP7_75t_R FILLER_266_386 ();
 DECAPx4_ASAP7_75t_R FILLER_266_426 ();
 FILLER_ASAP7_75t_R FILLER_266_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_467 ();
 DECAPx10_ASAP7_75t_R FILLER_266_472 ();
 FILLER_ASAP7_75t_R FILLER_266_501 ();
 DECAPx6_ASAP7_75t_R FILLER_266_529 ();
 DECAPx2_ASAP7_75t_R FILLER_266_543 ();
 DECAPx1_ASAP7_75t_R FILLER_266_562 ();
 DECAPx6_ASAP7_75t_R FILLER_266_580 ();
 FILLER_ASAP7_75t_R FILLER_266_594 ();
 DECAPx1_ASAP7_75t_R FILLER_266_602 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_606 ();
 DECAPx10_ASAP7_75t_R FILLER_266_621 ();
 DECAPx4_ASAP7_75t_R FILLER_266_643 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_653 ();
 DECAPx10_ASAP7_75t_R FILLER_266_668 ();
 DECAPx6_ASAP7_75t_R FILLER_266_690 ();
 DECAPx1_ASAP7_75t_R FILLER_266_704 ();
 DECAPx10_ASAP7_75t_R FILLER_266_714 ();
 DECAPx6_ASAP7_75t_R FILLER_266_736 ();
 DECAPx6_ASAP7_75t_R FILLER_266_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_767 ();
 FILLER_ASAP7_75t_R FILLER_266_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_266_805 ();
 DECAPx6_ASAP7_75t_R FILLER_266_815 ();
 DECAPx2_ASAP7_75t_R FILLER_266_829 ();
 DECAPx2_ASAP7_75t_R FILLER_266_843 ();
 FILLER_ASAP7_75t_R FILLER_266_849 ();
 DECAPx6_ASAP7_75t_R FILLER_266_860 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_874 ();
 FILLER_ASAP7_75t_R FILLER_266_893 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_266_905 ();
 DECAPx10_ASAP7_75t_R FILLER_267_2 ();
 DECAPx10_ASAP7_75t_R FILLER_267_24 ();
 DECAPx6_ASAP7_75t_R FILLER_267_46 ();
 DECAPx2_ASAP7_75t_R FILLER_267_60 ();
 DECAPx2_ASAP7_75t_R FILLER_267_95 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_267_101 ();
 DECAPx4_ASAP7_75t_R FILLER_267_110 ();
 DECAPx4_ASAP7_75t_R FILLER_267_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_267_144 ();
 DECAPx10_ASAP7_75t_R FILLER_267_173 ();
 DECAPx2_ASAP7_75t_R FILLER_267_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_267_201 ();
 DECAPx10_ASAP7_75t_R FILLER_267_233 ();
 DECAPx2_ASAP7_75t_R FILLER_267_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_268 ();
 FILLER_ASAP7_75t_R FILLER_267_321 ();
 DECAPx1_ASAP7_75t_R FILLER_267_337 ();
 DECAPx1_ASAP7_75t_R FILLER_267_367 ();
 DECAPx4_ASAP7_75t_R FILLER_267_374 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_384 ();
 DECAPx4_ASAP7_75t_R FILLER_267_425 ();
 FILLER_ASAP7_75t_R FILLER_267_435 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_456 ();
 DECAPx10_ASAP7_75t_R FILLER_267_471 ();
 DECAPx6_ASAP7_75t_R FILLER_267_493 ();
 DECAPx10_ASAP7_75t_R FILLER_267_533 ();
 DECAPx10_ASAP7_75t_R FILLER_267_555 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_267_577 ();
 DECAPx10_ASAP7_75t_R FILLER_267_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_267_612 ();
 DECAPx10_ASAP7_75t_R FILLER_267_627 ();
 DECAPx10_ASAP7_75t_R FILLER_267_649 ();
 DECAPx10_ASAP7_75t_R FILLER_267_671 ();
 DECAPx4_ASAP7_75t_R FILLER_267_693 ();
 FILLER_ASAP7_75t_R FILLER_267_703 ();
 DECAPx2_ASAP7_75t_R FILLER_267_711 ();
 FILLER_ASAP7_75t_R FILLER_267_717 ();
 DECAPx6_ASAP7_75t_R FILLER_267_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_744 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_763 ();
 FILLER_ASAP7_75t_R FILLER_267_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_267_794 ();
 DECAPx10_ASAP7_75t_R FILLER_267_801 ();
 DECAPx6_ASAP7_75t_R FILLER_267_839 ();
 DECAPx1_ASAP7_75t_R FILLER_267_868 ();
 FILLER_ASAP7_75t_R FILLER_267_898 ();
 FILLER_ASAP7_75t_R FILLER_267_927 ();
 DECAPx10_ASAP7_75t_R FILLER_268_2 ();
 DECAPx10_ASAP7_75t_R FILLER_268_24 ();
 DECAPx10_ASAP7_75t_R FILLER_268_46 ();
 DECAPx2_ASAP7_75t_R FILLER_268_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_74 ();
 DECAPx1_ASAP7_75t_R FILLER_268_84 ();
 DECAPx6_ASAP7_75t_R FILLER_268_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_144 ();
 DECAPx6_ASAP7_75t_R FILLER_268_156 ();
 DECAPx1_ASAP7_75t_R FILLER_268_170 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_182 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_268_195 ();
 DECAPx1_ASAP7_75t_R FILLER_268_201 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_205 ();
 DECAPx10_ASAP7_75t_R FILLER_268_212 ();
 FILLER_ASAP7_75t_R FILLER_268_234 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_248 ();
 DECAPx6_ASAP7_75t_R FILLER_268_252 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_268_266 ();
 DECAPx1_ASAP7_75t_R FILLER_268_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_276 ();
 FILLER_ASAP7_75t_R FILLER_268_283 ();
 DECAPx6_ASAP7_75t_R FILLER_268_288 ();
 FILLER_ASAP7_75t_R FILLER_268_302 ();
 FILLER_ASAP7_75t_R FILLER_268_319 ();
 DECAPx2_ASAP7_75t_R FILLER_268_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_345 ();
 DECAPx6_ASAP7_75t_R FILLER_268_361 ();
 DECAPx1_ASAP7_75t_R FILLER_268_375 ();
 FILLER_ASAP7_75t_R FILLER_268_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_409 ();
 DECAPx2_ASAP7_75t_R FILLER_268_416 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_422 ();
 DECAPx10_ASAP7_75t_R FILLER_268_426 ();
 DECAPx4_ASAP7_75t_R FILLER_268_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_458 ();
 FILLER_ASAP7_75t_R FILLER_268_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_469 ();
 DECAPx6_ASAP7_75t_R FILLER_268_494 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_508 ();
 DECAPx1_ASAP7_75t_R FILLER_268_515 ();
 DECAPx2_ASAP7_75t_R FILLER_268_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_538 ();
 FILLER_ASAP7_75t_R FILLER_268_545 ();
 DECAPx2_ASAP7_75t_R FILLER_268_557 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_268_563 ();
 DECAPx10_ASAP7_75t_R FILLER_268_592 ();
 DECAPx2_ASAP7_75t_R FILLER_268_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_268_620 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_629 ();
 DECAPx2_ASAP7_75t_R FILLER_268_643 ();
 DECAPx6_ASAP7_75t_R FILLER_268_659 ();
 DECAPx2_ASAP7_75t_R FILLER_268_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_679 ();
 DECAPx6_ASAP7_75t_R FILLER_268_686 ();
 FILLER_ASAP7_75t_R FILLER_268_700 ();
 DECAPx1_ASAP7_75t_R FILLER_268_714 ();
 DECAPx10_ASAP7_75t_R FILLER_268_750 ();
 DECAPx10_ASAP7_75t_R FILLER_268_772 ();
 DECAPx4_ASAP7_75t_R FILLER_268_794 ();
 FILLER_ASAP7_75t_R FILLER_268_804 ();
 DECAPx2_ASAP7_75t_R FILLER_268_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_817 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_844 ();
 DECAPx1_ASAP7_75t_R FILLER_268_896 ();
 FILLERxp5_ASAP7_75t_R FILLER_268_900 ();
 DECAPx10_ASAP7_75t_R FILLER_269_2 ();
 DECAPx10_ASAP7_75t_R FILLER_269_24 ();
 DECAPx10_ASAP7_75t_R FILLER_269_46 ();
 DECAPx6_ASAP7_75t_R FILLER_269_68 ();
 DECAPx1_ASAP7_75t_R FILLER_269_82 ();
 FILLER_ASAP7_75t_R FILLER_269_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_126 ();
 DECAPx2_ASAP7_75t_R FILLER_269_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_141 ();
 DECAPx10_ASAP7_75t_R FILLER_269_154 ();
 FILLER_ASAP7_75t_R FILLER_269_176 ();
 DECAPx1_ASAP7_75t_R FILLER_269_210 ();
 DECAPx1_ASAP7_75t_R FILLER_269_260 ();
 DECAPx10_ASAP7_75t_R FILLER_269_270 ();
 DECAPx6_ASAP7_75t_R FILLER_269_292 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_306 ();
 DECAPx2_ASAP7_75t_R FILLER_269_312 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_347 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_394 ();
 DECAPx2_ASAP7_75t_R FILLER_269_413 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_419 ();
 DECAPx10_ASAP7_75t_R FILLER_269_436 ();
 DECAPx6_ASAP7_75t_R FILLER_269_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_472 ();
 DECAPx10_ASAP7_75t_R FILLER_269_503 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_535 ();
 DECAPx10_ASAP7_75t_R FILLER_269_570 ();
 DECAPx2_ASAP7_75t_R FILLER_269_592 ();
 FILLER_ASAP7_75t_R FILLER_269_598 ();
 DECAPx4_ASAP7_75t_R FILLER_269_606 ();
 FILLER_ASAP7_75t_R FILLER_269_622 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_630 ();
 DECAPx1_ASAP7_75t_R FILLER_269_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_645 ();
 DECAPx1_ASAP7_75t_R FILLER_269_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_657 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_664 ();
 FILLER_ASAP7_75t_R FILLER_269_673 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_690 ();
 DECAPx2_ASAP7_75t_R FILLER_269_713 ();
 FILLER_ASAP7_75t_R FILLER_269_719 ();
 FILLER_ASAP7_75t_R FILLER_269_733 ();
 DECAPx4_ASAP7_75t_R FILLER_269_743 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_792 ();
 FILLER_ASAP7_75t_R FILLER_269_801 ();
 DECAPx2_ASAP7_75t_R FILLER_269_838 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_269_857 ();
 DECAPx10_ASAP7_75t_R FILLER_269_866 ();
 DECAPx1_ASAP7_75t_R FILLER_269_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_269_892 ();
 FILLER_ASAP7_75t_R FILLER_269_908 ();
 FILLER_ASAP7_75t_R FILLER_269_927 ();
 DECAPx10_ASAP7_75t_R FILLER_270_2 ();
 DECAPx10_ASAP7_75t_R FILLER_270_24 ();
 DECAPx10_ASAP7_75t_R FILLER_270_46 ();
 DECAPx10_ASAP7_75t_R FILLER_270_68 ();
 DECAPx2_ASAP7_75t_R FILLER_270_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_96 ();
 DECAPx6_ASAP7_75t_R FILLER_270_141 ();
 FILLER_ASAP7_75t_R FILLER_270_155 ();
 DECAPx1_ASAP7_75t_R FILLER_270_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_187 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_231 ();
 DECAPx6_ASAP7_75t_R FILLER_270_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_311 ();
 DECAPx6_ASAP7_75t_R FILLER_270_318 ();
 DECAPx1_ASAP7_75t_R FILLER_270_332 ();
 FILLER_ASAP7_75t_R FILLER_270_339 ();
 DECAPx1_ASAP7_75t_R FILLER_270_362 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_366 ();
 DECAPx2_ASAP7_75t_R FILLER_270_414 ();
 DECAPx6_ASAP7_75t_R FILLER_270_446 ();
 FILLER_ASAP7_75t_R FILLER_270_460 ();
 DECAPx6_ASAP7_75t_R FILLER_270_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_488 ();
 DECAPx1_ASAP7_75t_R FILLER_270_500 ();
 DECAPx6_ASAP7_75t_R FILLER_270_519 ();
 DECAPx2_ASAP7_75t_R FILLER_270_533 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_539 ();
 DECAPx1_ASAP7_75t_R FILLER_270_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_552 ();
 DECAPx4_ASAP7_75t_R FILLER_270_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_566 ();
 FILLER_ASAP7_75t_R FILLER_270_573 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_270_581 ();
 FILLER_ASAP7_75t_R FILLER_270_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_270_679 ();
 DECAPx4_ASAP7_75t_R FILLER_270_708 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_270_718 ();
 DECAPx10_ASAP7_75t_R FILLER_270_728 ();
 DECAPx4_ASAP7_75t_R FILLER_270_758 ();
 FILLER_ASAP7_75t_R FILLER_270_768 ();
 DECAPx1_ASAP7_75t_R FILLER_270_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_799 ();
 DECAPx10_ASAP7_75t_R FILLER_270_826 ();
 DECAPx10_ASAP7_75t_R FILLER_270_848 ();
 FILLERxp5_ASAP7_75t_R FILLER_270_870 ();
 DECAPx4_ASAP7_75t_R FILLER_270_877 ();
 FILLER_ASAP7_75t_R FILLER_270_927 ();
 DECAPx10_ASAP7_75t_R FILLER_271_2 ();
 DECAPx10_ASAP7_75t_R FILLER_271_24 ();
 DECAPx10_ASAP7_75t_R FILLER_271_46 ();
 DECAPx4_ASAP7_75t_R FILLER_271_68 ();
 DECAPx10_ASAP7_75t_R FILLER_271_90 ();
 FILLER_ASAP7_75t_R FILLER_271_112 ();
 DECAPx1_ASAP7_75t_R FILLER_271_120 ();
 DECAPx6_ASAP7_75t_R FILLER_271_127 ();
 DECAPx1_ASAP7_75t_R FILLER_271_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_145 ();
 DECAPx6_ASAP7_75t_R FILLER_271_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_192 ();
 DECAPx4_ASAP7_75t_R FILLER_271_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_206 ();
 FILLER_ASAP7_75t_R FILLER_271_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_251 ();
 DECAPx2_ASAP7_75t_R FILLER_271_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_271_311 ();
 DECAPx6_ASAP7_75t_R FILLER_271_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_336 ();
 FILLER_ASAP7_75t_R FILLER_271_366 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_382 ();
 DECAPx1_ASAP7_75t_R FILLER_271_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_390 ();
 DECAPx6_ASAP7_75t_R FILLER_271_397 ();
 DECAPx1_ASAP7_75t_R FILLER_271_411 ();
 DECAPx4_ASAP7_75t_R FILLER_271_420 ();
 FILLER_ASAP7_75t_R FILLER_271_430 ();
 DECAPx4_ASAP7_75t_R FILLER_271_441 ();
 DECAPx1_ASAP7_75t_R FILLER_271_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_481 ();
 DECAPx4_ASAP7_75t_R FILLER_271_492 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_505 ();
 DECAPx10_ASAP7_75t_R FILLER_271_509 ();
 DECAPx10_ASAP7_75t_R FILLER_271_531 ();
 DECAPx6_ASAP7_75t_R FILLER_271_553 ();
 DECAPx2_ASAP7_75t_R FILLER_271_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_573 ();
 DECAPx1_ASAP7_75t_R FILLER_271_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_584 ();
 FILLER_ASAP7_75t_R FILLER_271_608 ();
 DECAPx10_ASAP7_75t_R FILLER_271_619 ();
 DECAPx10_ASAP7_75t_R FILLER_271_641 ();
 DECAPx6_ASAP7_75t_R FILLER_271_663 ();
 DECAPx10_ASAP7_75t_R FILLER_271_695 ();
 DECAPx4_ASAP7_75t_R FILLER_271_717 ();
 FILLER_ASAP7_75t_R FILLER_271_727 ();
 FILLER_ASAP7_75t_R FILLER_271_761 ();
 DECAPx2_ASAP7_75t_R FILLER_271_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_271_779 ();
 DECAPx10_ASAP7_75t_R FILLER_271_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_813 ();
 DECAPx10_ASAP7_75t_R FILLER_271_817 ();
 DECAPx10_ASAP7_75t_R FILLER_271_839 ();
 DECAPx6_ASAP7_75t_R FILLER_271_861 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_271_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_271_890 ();
 FILLER_ASAP7_75t_R FILLER_271_907 ();
 FILLER_ASAP7_75t_R FILLER_271_923 ();
 FILLER_ASAP7_75t_R FILLER_271_927 ();
 DECAPx10_ASAP7_75t_R FILLER_272_7 ();
 DECAPx10_ASAP7_75t_R FILLER_272_29 ();
 DECAPx6_ASAP7_75t_R FILLER_272_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_65 ();
 DECAPx10_ASAP7_75t_R FILLER_272_97 ();
 DECAPx6_ASAP7_75t_R FILLER_272_119 ();
 DECAPx1_ASAP7_75t_R FILLER_272_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_137 ();
 DECAPx2_ASAP7_75t_R FILLER_272_144 ();
 FILLER_ASAP7_75t_R FILLER_272_150 ();
 FILLER_ASAP7_75t_R FILLER_272_158 ();
 DECAPx10_ASAP7_75t_R FILLER_272_172 ();
 DECAPx10_ASAP7_75t_R FILLER_272_194 ();
 DECAPx10_ASAP7_75t_R FILLER_272_216 ();
 DECAPx6_ASAP7_75t_R FILLER_272_238 ();
 DECAPx2_ASAP7_75t_R FILLER_272_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_284 ();
 FILLER_ASAP7_75t_R FILLER_272_288 ();
 FILLER_ASAP7_75t_R FILLER_272_302 ();
 DECAPx10_ASAP7_75t_R FILLER_272_310 ();
 DECAPx4_ASAP7_75t_R FILLER_272_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_355 ();
 DECAPx10_ASAP7_75t_R FILLER_272_372 ();
 DECAPx2_ASAP7_75t_R FILLER_272_394 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_400 ();
 DECAPx1_ASAP7_75t_R FILLER_272_409 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_427 ();
 FILLER_ASAP7_75t_R FILLER_272_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_461 ();
 DECAPx10_ASAP7_75t_R FILLER_272_483 ();
 DECAPx6_ASAP7_75t_R FILLER_272_505 ();
 DECAPx1_ASAP7_75t_R FILLER_272_519 ();
 DECAPx4_ASAP7_75t_R FILLER_272_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_547 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_559 ();
 DECAPx2_ASAP7_75t_R FILLER_272_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_574 ();
 DECAPx6_ASAP7_75t_R FILLER_272_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_605 ();
 DECAPx10_ASAP7_75t_R FILLER_272_612 ();
 DECAPx10_ASAP7_75t_R FILLER_272_634 ();
 DECAPx10_ASAP7_75t_R FILLER_272_656 ();
 DECAPx10_ASAP7_75t_R FILLER_272_678 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_700 ();
 DECAPx1_ASAP7_75t_R FILLER_272_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_719 ();
 FILLER_ASAP7_75t_R FILLER_272_764 ();
 DECAPx6_ASAP7_75t_R FILLER_272_778 ();
 FILLER_ASAP7_75t_R FILLER_272_792 ();
 DECAPx10_ASAP7_75t_R FILLER_272_800 ();
 DECAPx4_ASAP7_75t_R FILLER_272_822 ();
 DECAPx1_ASAP7_75t_R FILLER_272_838 ();
 FILLERxp5_ASAP7_75t_R FILLER_272_855 ();
 DECAPx4_ASAP7_75t_R FILLER_272_868 ();
 FILLER_ASAP7_75t_R FILLER_272_878 ();
 DECAPx6_ASAP7_75t_R FILLER_272_883 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_272_897 ();
 DECAPx10_ASAP7_75t_R FILLER_273_7 ();
 DECAPx10_ASAP7_75t_R FILLER_273_29 ();
 DECAPx10_ASAP7_75t_R FILLER_273_51 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_73 ();
 DECAPx2_ASAP7_75t_R FILLER_273_102 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_108 ();
 FILLER_ASAP7_75t_R FILLER_273_117 ();
 DECAPx2_ASAP7_75t_R FILLER_273_122 ();
 FILLER_ASAP7_75t_R FILLER_273_128 ();
 DECAPx10_ASAP7_75t_R FILLER_273_159 ();
 DECAPx10_ASAP7_75t_R FILLER_273_181 ();
 DECAPx10_ASAP7_75t_R FILLER_273_203 ();
 DECAPx10_ASAP7_75t_R FILLER_273_225 ();
 DECAPx10_ASAP7_75t_R FILLER_273_247 ();
 DECAPx10_ASAP7_75t_R FILLER_273_269 ();
 DECAPx1_ASAP7_75t_R FILLER_273_291 ();
 DECAPx6_ASAP7_75t_R FILLER_273_298 ();
 DECAPx2_ASAP7_75t_R FILLER_273_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_318 ();
 DECAPx2_ASAP7_75t_R FILLER_273_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_351 ();
 DECAPx10_ASAP7_75t_R FILLER_273_361 ();
 DECAPx4_ASAP7_75t_R FILLER_273_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_407 ();
 DECAPx10_ASAP7_75t_R FILLER_273_422 ();
 DECAPx2_ASAP7_75t_R FILLER_273_444 ();
 DECAPx4_ASAP7_75t_R FILLER_273_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_463 ();
 DECAPx10_ASAP7_75t_R FILLER_273_467 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_489 ();
 DECAPx4_ASAP7_75t_R FILLER_273_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_509 ();
 DECAPx10_ASAP7_75t_R FILLER_273_536 ();
 DECAPx1_ASAP7_75t_R FILLER_273_558 ();
 DECAPx6_ASAP7_75t_R FILLER_273_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_596 ();
 DECAPx10_ASAP7_75t_R FILLER_273_603 ();
 DECAPx6_ASAP7_75t_R FILLER_273_625 ();
 DECAPx2_ASAP7_75t_R FILLER_273_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_645 ();
 FILLER_ASAP7_75t_R FILLER_273_661 ();
 DECAPx10_ASAP7_75t_R FILLER_273_669 ();
 DECAPx4_ASAP7_75t_R FILLER_273_691 ();
 FILLER_ASAP7_75t_R FILLER_273_701 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_765 ();
 DECAPx2_ASAP7_75t_R FILLER_273_778 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_273_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_273_829 ();
 FILLER_ASAP7_75t_R FILLER_273_840 ();
 FILLER_ASAP7_75t_R FILLER_273_854 ();
 DECAPx6_ASAP7_75t_R FILLER_273_891 ();
 DECAPx1_ASAP7_75t_R FILLER_273_905 ();
 FILLER_ASAP7_75t_R FILLER_273_927 ();
 DECAPx10_ASAP7_75t_R FILLER_274_2 ();
 DECAPx10_ASAP7_75t_R FILLER_274_24 ();
 DECAPx10_ASAP7_75t_R FILLER_274_46 ();
 DECAPx4_ASAP7_75t_R FILLER_274_68 ();
 FILLER_ASAP7_75t_R FILLER_274_78 ();
 DECAPx1_ASAP7_75t_R FILLER_274_95 ();
 DECAPx1_ASAP7_75t_R FILLER_274_131 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_141 ();
 DECAPx10_ASAP7_75t_R FILLER_274_147 ();
 FILLER_ASAP7_75t_R FILLER_274_169 ();
 DECAPx2_ASAP7_75t_R FILLER_274_186 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_192 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_201 ();
 DECAPx2_ASAP7_75t_R FILLER_274_219 ();
 DECAPx1_ASAP7_75t_R FILLER_274_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_243 ();
 FILLER_ASAP7_75t_R FILLER_274_250 ();
 DECAPx10_ASAP7_75t_R FILLER_274_258 ();
 FILLER_ASAP7_75t_R FILLER_274_280 ();
 DECAPx2_ASAP7_75t_R FILLER_274_288 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_294 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_313 ();
 DECAPx10_ASAP7_75t_R FILLER_274_354 ();
 DECAPx6_ASAP7_75t_R FILLER_274_376 ();
 DECAPx2_ASAP7_75t_R FILLER_274_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_396 ();
 FILLER_ASAP7_75t_R FILLER_274_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_408 ();
 DECAPx10_ASAP7_75t_R FILLER_274_415 ();
 DECAPx2_ASAP7_75t_R FILLER_274_437 ();
 DECAPx2_ASAP7_75t_R FILLER_274_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_464 ();
 DECAPx10_ASAP7_75t_R FILLER_274_470 ();
 DECAPx2_ASAP7_75t_R FILLER_274_492 ();
 DECAPx4_ASAP7_75t_R FILLER_274_521 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_531 ();
 FILLER_ASAP7_75t_R FILLER_274_542 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_547 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_554 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_575 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_592 ();
 DECAPx1_ASAP7_75t_R FILLER_274_603 ();
 DECAPx1_ASAP7_75t_R FILLER_274_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_659 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_675 ();
 DECAPx6_ASAP7_75t_R FILLER_274_686 ();
 DECAPx1_ASAP7_75t_R FILLER_274_700 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_722 ();
 DECAPx1_ASAP7_75t_R FILLER_274_746 ();
 FILLER_ASAP7_75t_R FILLER_274_761 ();
 DECAPx6_ASAP7_75t_R FILLER_274_773 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_274_787 ();
 DECAPx1_ASAP7_75t_R FILLER_274_797 ();
 FILLER_ASAP7_75t_R FILLER_274_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_274_817 ();
 DECAPx1_ASAP7_75t_R FILLER_274_853 ();
 DECAPx4_ASAP7_75t_R FILLER_274_869 ();
 DECAPx2_ASAP7_75t_R FILLER_274_887 ();
 FILLER_ASAP7_75t_R FILLER_274_893 ();
 DECAPx4_ASAP7_75t_R FILLER_274_901 ();
 DECAPx10_ASAP7_75t_R FILLER_275_2 ();
 DECAPx10_ASAP7_75t_R FILLER_275_24 ();
 DECAPx10_ASAP7_75t_R FILLER_275_46 ();
 DECAPx10_ASAP7_75t_R FILLER_275_68 ();
 DECAPx6_ASAP7_75t_R FILLER_275_90 ();
 DECAPx2_ASAP7_75t_R FILLER_275_104 ();
 DECAPx1_ASAP7_75t_R FILLER_275_119 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_129 ();
 DECAPx4_ASAP7_75t_R FILLER_275_136 ();
 FILLER_ASAP7_75t_R FILLER_275_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_164 ();
 FILLER_ASAP7_75t_R FILLER_275_196 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_235 ();
 FILLER_ASAP7_75t_R FILLER_275_258 ();
 DECAPx1_ASAP7_75t_R FILLER_275_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_305 ();
 FILLER_ASAP7_75t_R FILLER_275_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_328 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_343 ();
 DECAPx10_ASAP7_75t_R FILLER_275_352 ();
 DECAPx1_ASAP7_75t_R FILLER_275_374 ();
 DECAPx4_ASAP7_75t_R FILLER_275_416 ();
 DECAPx4_ASAP7_75t_R FILLER_275_429 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_439 ();
 DECAPx4_ASAP7_75t_R FILLER_275_445 ();
 DECAPx6_ASAP7_75t_R FILLER_275_507 ();
 DECAPx1_ASAP7_75t_R FILLER_275_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_525 ();
 DECAPx6_ASAP7_75t_R FILLER_275_568 ();
 DECAPx1_ASAP7_75t_R FILLER_275_582 ();
 DECAPx1_ASAP7_75t_R FILLER_275_592 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_596 ();
 DECAPx4_ASAP7_75t_R FILLER_275_603 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_275_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_631 ();
 DECAPx1_ASAP7_75t_R FILLER_275_645 ();
 DECAPx1_ASAP7_75t_R FILLER_275_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_673 ();
 DECAPx6_ASAP7_75t_R FILLER_275_715 ();
 DECAPx2_ASAP7_75t_R FILLER_275_729 ();
 DECAPx10_ASAP7_75t_R FILLER_275_738 ();
 FILLER_ASAP7_75t_R FILLER_275_760 ();
 DECAPx4_ASAP7_75t_R FILLER_275_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_782 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_797 ();
 FILLER_ASAP7_75t_R FILLER_275_831 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_842 ();
 DECAPx10_ASAP7_75t_R FILLER_275_846 ();
 DECAPx4_ASAP7_75t_R FILLER_275_868 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_878 ();
 FILLERxp5_ASAP7_75t_R FILLER_275_905 ();
 FILLER_ASAP7_75t_R FILLER_275_913 ();
 FILLER_ASAP7_75t_R FILLER_275_927 ();
 DECAPx10_ASAP7_75t_R FILLER_276_2 ();
 DECAPx10_ASAP7_75t_R FILLER_276_24 ();
 DECAPx10_ASAP7_75t_R FILLER_276_46 ();
 DECAPx10_ASAP7_75t_R FILLER_276_68 ();
 DECAPx10_ASAP7_75t_R FILLER_276_90 ();
 DECAPx1_ASAP7_75t_R FILLER_276_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_116 ();
 DECAPx4_ASAP7_75t_R FILLER_276_143 ();
 DECAPx1_ASAP7_75t_R FILLER_276_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_220 ();
 DECAPx2_ASAP7_75t_R FILLER_276_253 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_276 ();
 DECAPx1_ASAP7_75t_R FILLER_276_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_287 ();
 DECAPx2_ASAP7_75t_R FILLER_276_291 ();
 FILLER_ASAP7_75t_R FILLER_276_297 ();
 DECAPx4_ASAP7_75t_R FILLER_276_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_367 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_376 ();
 FILLER_ASAP7_75t_R FILLER_276_391 ();
 DECAPx10_ASAP7_75t_R FILLER_276_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_430 ();
 DECAPx6_ASAP7_75t_R FILLER_276_446 ();
 FILLER_ASAP7_75t_R FILLER_276_460 ();
 DECAPx1_ASAP7_75t_R FILLER_276_464 ();
 DECAPx4_ASAP7_75t_R FILLER_276_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_509 ();
 DECAPx4_ASAP7_75t_R FILLER_276_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_523 ();
 DECAPx10_ASAP7_75t_R FILLER_276_540 ();
 DECAPx2_ASAP7_75t_R FILLER_276_562 ();
 FILLER_ASAP7_75t_R FILLER_276_568 ();
 DECAPx6_ASAP7_75t_R FILLER_276_590 ();
 DECAPx1_ASAP7_75t_R FILLER_276_604 ();
 DECAPx1_ASAP7_75t_R FILLER_276_614 ();
 DECAPx2_ASAP7_75t_R FILLER_276_624 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_639 ();
 DECAPx1_ASAP7_75t_R FILLER_276_658 ();
 FILLER_ASAP7_75t_R FILLER_276_690 ();
 DECAPx10_ASAP7_75t_R FILLER_276_708 ();
 DECAPx10_ASAP7_75t_R FILLER_276_730 ();
 DECAPx6_ASAP7_75t_R FILLER_276_752 ();
 DECAPx2_ASAP7_75t_R FILLER_276_766 ();
 DECAPx10_ASAP7_75t_R FILLER_276_786 ();
 DECAPx10_ASAP7_75t_R FILLER_276_808 ();
 DECAPx6_ASAP7_75t_R FILLER_276_830 ();
 DECAPx1_ASAP7_75t_R FILLER_276_844 ();
 FILLERxp5_ASAP7_75t_R FILLER_276_848 ();
 DECAPx6_ASAP7_75t_R FILLER_276_854 ();
 DECAPx2_ASAP7_75t_R FILLER_276_868 ();
 DECAPx2_ASAP7_75t_R FILLER_276_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_891 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_276_897 ();
 DECAPx10_ASAP7_75t_R FILLER_277_2 ();
 DECAPx10_ASAP7_75t_R FILLER_277_24 ();
 DECAPx10_ASAP7_75t_R FILLER_277_46 ();
 DECAPx4_ASAP7_75t_R FILLER_277_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_78 ();
 FILLER_ASAP7_75t_R FILLER_277_88 ();
 DECAPx10_ASAP7_75t_R FILLER_277_110 ();
 FILLER_ASAP7_75t_R FILLER_277_135 ();
 DECAPx2_ASAP7_75t_R FILLER_277_153 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_159 ();
 DECAPx4_ASAP7_75t_R FILLER_277_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_181 ();
 DECAPx1_ASAP7_75t_R FILLER_277_196 ();
 DECAPx1_ASAP7_75t_R FILLER_277_239 ();
 DECAPx1_ASAP7_75t_R FILLER_277_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_261 ();
 DECAPx10_ASAP7_75t_R FILLER_277_268 ();
 DECAPx6_ASAP7_75t_R FILLER_277_290 ();
 DECAPx1_ASAP7_75t_R FILLER_277_304 ();
 DECAPx10_ASAP7_75t_R FILLER_277_314 ();
 DECAPx4_ASAP7_75t_R FILLER_277_336 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_346 ();
 DECAPx10_ASAP7_75t_R FILLER_277_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_418 ();
 DECAPx2_ASAP7_75t_R FILLER_277_442 ();
 FILLER_ASAP7_75t_R FILLER_277_448 ();
 DECAPx2_ASAP7_75t_R FILLER_277_460 ();
 FILLER_ASAP7_75t_R FILLER_277_466 ();
 DECAPx1_ASAP7_75t_R FILLER_277_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_475 ();
 DECAPx2_ASAP7_75t_R FILLER_277_488 ();
 DECAPx2_ASAP7_75t_R FILLER_277_525 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_531 ();
 DECAPx10_ASAP7_75t_R FILLER_277_540 ();
 DECAPx1_ASAP7_75t_R FILLER_277_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_566 ();
 DECAPx10_ASAP7_75t_R FILLER_277_621 ();
 DECAPx6_ASAP7_75t_R FILLER_277_643 ();
 DECAPx6_ASAP7_75t_R FILLER_277_663 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_677 ();
 DECAPx2_ASAP7_75t_R FILLER_277_684 ();
 DECAPx2_ASAP7_75t_R FILLER_277_710 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_716 ();
 DECAPx6_ASAP7_75t_R FILLER_277_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_740 ();
 DECAPx6_ASAP7_75t_R FILLER_277_751 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_765 ();
 DECAPx10_ASAP7_75t_R FILLER_277_797 ();
 DECAPx2_ASAP7_75t_R FILLER_277_819 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_825 ();
 DECAPx4_ASAP7_75t_R FILLER_277_834 ();
 FILLER_ASAP7_75t_R FILLER_277_844 ();
 DECAPx2_ASAP7_75t_R FILLER_277_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_868 ();
 DECAPx2_ASAP7_75t_R FILLER_277_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_887 ();
 DECAPx4_ASAP7_75t_R FILLER_277_895 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_277_905 ();
 DECAPx4_ASAP7_75t_R FILLER_277_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_277_924 ();
 DECAPx1_ASAP7_75t_R FILLER_277_930 ();
 DECAPx10_ASAP7_75t_R FILLER_278_2 ();
 DECAPx10_ASAP7_75t_R FILLER_278_24 ();
 DECAPx10_ASAP7_75t_R FILLER_278_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_95 ();
 DECAPx10_ASAP7_75t_R FILLER_278_110 ();
 DECAPx2_ASAP7_75t_R FILLER_278_132 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_138 ();
 DECAPx2_ASAP7_75t_R FILLER_278_145 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_151 ();
 DECAPx10_ASAP7_75t_R FILLER_278_158 ();
 DECAPx10_ASAP7_75t_R FILLER_278_180 ();
 DECAPx2_ASAP7_75t_R FILLER_278_208 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_226 ();
 DECAPx10_ASAP7_75t_R FILLER_278_230 ();
 DECAPx6_ASAP7_75t_R FILLER_278_252 ();
 DECAPx1_ASAP7_75t_R FILLER_278_266 ();
 DECAPx6_ASAP7_75t_R FILLER_278_302 ();
 FILLER_ASAP7_75t_R FILLER_278_316 ();
 DECAPx10_ASAP7_75t_R FILLER_278_324 ();
 DECAPx1_ASAP7_75t_R FILLER_278_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_350 ();
 FILLER_ASAP7_75t_R FILLER_278_371 ();
 FILLER_ASAP7_75t_R FILLER_278_379 ();
 DECAPx4_ASAP7_75t_R FILLER_278_392 ();
 DECAPx2_ASAP7_75t_R FILLER_278_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_420 ();
 DECAPx10_ASAP7_75t_R FILLER_278_427 ();
 DECAPx1_ASAP7_75t_R FILLER_278_449 ();
 DECAPx10_ASAP7_75t_R FILLER_278_467 ();
 DECAPx6_ASAP7_75t_R FILLER_278_489 ();
 FILLER_ASAP7_75t_R FILLER_278_503 ();
 DECAPx2_ASAP7_75t_R FILLER_278_508 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_514 ();
 DECAPx4_ASAP7_75t_R FILLER_278_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_537 ();
 DECAPx6_ASAP7_75t_R FILLER_278_549 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_563 ();
 DECAPx10_ASAP7_75t_R FILLER_278_597 ();
 FILLER_ASAP7_75t_R FILLER_278_619 ();
 DECAPx10_ASAP7_75t_R FILLER_278_629 ();
 DECAPx10_ASAP7_75t_R FILLER_278_651 ();
 DECAPx10_ASAP7_75t_R FILLER_278_673 ();
 DECAPx10_ASAP7_75t_R FILLER_278_695 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_746 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_278_750 ();
 DECAPx6_ASAP7_75t_R FILLER_278_759 ();
 FILLER_ASAP7_75t_R FILLER_278_773 ();
 DECAPx4_ASAP7_75t_R FILLER_278_792 ();
 FILLER_ASAP7_75t_R FILLER_278_802 ();
 DECAPx6_ASAP7_75t_R FILLER_278_812 ();
 FILLER_ASAP7_75t_R FILLER_278_836 ();
 DECAPx4_ASAP7_75t_R FILLER_278_877 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_278_887 ();
 FILLERxp5_ASAP7_75t_R FILLER_278_904 ();
 DECAPx10_ASAP7_75t_R FILLER_278_908 ();
 DECAPx1_ASAP7_75t_R FILLER_278_930 ();
 DECAPx10_ASAP7_75t_R FILLER_279_2 ();
 DECAPx10_ASAP7_75t_R FILLER_279_24 ();
 DECAPx10_ASAP7_75t_R FILLER_279_46 ();
 DECAPx2_ASAP7_75t_R FILLER_279_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_74 ();
 FILLER_ASAP7_75t_R FILLER_279_81 ();
 DECAPx1_ASAP7_75t_R FILLER_279_89 ();
 DECAPx4_ASAP7_75t_R FILLER_279_99 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_116 ();
 DECAPx10_ASAP7_75t_R FILLER_279_131 ();
 DECAPx6_ASAP7_75t_R FILLER_279_153 ();
 DECAPx1_ASAP7_75t_R FILLER_279_167 ();
 FILLER_ASAP7_75t_R FILLER_279_177 ();
 DECAPx10_ASAP7_75t_R FILLER_279_188 ();
 DECAPx10_ASAP7_75t_R FILLER_279_210 ();
 DECAPx2_ASAP7_75t_R FILLER_279_232 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_238 ();
 DECAPx6_ASAP7_75t_R FILLER_279_244 ();
 DECAPx1_ASAP7_75t_R FILLER_279_258 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_269 ();
 DECAPx2_ASAP7_75t_R FILLER_279_308 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_321 ();
 DECAPx6_ASAP7_75t_R FILLER_279_347 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_361 ();
 DECAPx10_ASAP7_75t_R FILLER_279_370 ();
 DECAPx1_ASAP7_75t_R FILLER_279_392 ();
 DECAPx6_ASAP7_75t_R FILLER_279_422 ();
 DECAPx1_ASAP7_75t_R FILLER_279_436 ();
 DECAPx1_ASAP7_75t_R FILLER_279_449 ();
 DECAPx10_ASAP7_75t_R FILLER_279_467 ();
 DECAPx4_ASAP7_75t_R FILLER_279_489 ();
 DECAPx10_ASAP7_75t_R FILLER_279_502 ();
 DECAPx4_ASAP7_75t_R FILLER_279_524 ();
 FILLER_ASAP7_75t_R FILLER_279_534 ();
 FILLER_ASAP7_75t_R FILLER_279_558 ();
 DECAPx10_ASAP7_75t_R FILLER_279_566 ();
 DECAPx10_ASAP7_75t_R FILLER_279_588 ();
 DECAPx10_ASAP7_75t_R FILLER_279_610 ();
 DECAPx2_ASAP7_75t_R FILLER_279_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_644 ();
 DECAPx10_ASAP7_75t_R FILLER_279_650 ();
 DECAPx6_ASAP7_75t_R FILLER_279_672 ();
 DECAPx2_ASAP7_75t_R FILLER_279_686 ();
 DECAPx4_ASAP7_75t_R FILLER_279_698 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_708 ();
 FILLER_ASAP7_75t_R FILLER_279_758 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_768 ();
 DECAPx6_ASAP7_75t_R FILLER_279_772 ();
 DECAPx1_ASAP7_75t_R FILLER_279_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_279_790 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_279_823 ();
 DECAPx2_ASAP7_75t_R FILLER_279_882 ();
 FILLER_ASAP7_75t_R FILLER_279_898 ();
 DECAPx1_ASAP7_75t_R FILLER_279_921 ();
 FILLER_ASAP7_75t_R FILLER_279_927 ();
 DECAPx10_ASAP7_75t_R FILLER_280_2 ();
 DECAPx10_ASAP7_75t_R FILLER_280_24 ();
 DECAPx10_ASAP7_75t_R FILLER_280_46 ();
 DECAPx2_ASAP7_75t_R FILLER_280_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_280_135 ();
 DECAPx4_ASAP7_75t_R FILLER_280_144 ();
 FILLER_ASAP7_75t_R FILLER_280_154 ();
 FILLER_ASAP7_75t_R FILLER_280_165 ();
 DECAPx4_ASAP7_75t_R FILLER_280_193 ();
 DECAPx6_ASAP7_75t_R FILLER_280_209 ();
 DECAPx1_ASAP7_75t_R FILLER_280_230 ();
 DECAPx4_ASAP7_75t_R FILLER_280_240 ();
 FILLER_ASAP7_75t_R FILLER_280_250 ();
 DECAPx2_ASAP7_75t_R FILLER_280_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_284 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_280_288 ();
 DECAPx4_ASAP7_75t_R FILLER_280_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_313 ();
 FILLER_ASAP7_75t_R FILLER_280_322 ();
 DECAPx10_ASAP7_75t_R FILLER_280_356 ();
 DECAPx2_ASAP7_75t_R FILLER_280_378 ();
 FILLER_ASAP7_75t_R FILLER_280_384 ();
 DECAPx2_ASAP7_75t_R FILLER_280_403 ();
 FILLER_ASAP7_75t_R FILLER_280_409 ();
 DECAPx4_ASAP7_75t_R FILLER_280_414 ();
 DECAPx6_ASAP7_75t_R FILLER_280_441 ();
 DECAPx2_ASAP7_75t_R FILLER_280_455 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_461 ();
 DECAPx4_ASAP7_75t_R FILLER_280_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_474 ();
 DECAPx2_ASAP7_75t_R FILLER_280_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_484 ();
 DECAPx2_ASAP7_75t_R FILLER_280_497 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_280_503 ();
 FILLER_ASAP7_75t_R FILLER_280_520 ();
 DECAPx2_ASAP7_75t_R FILLER_280_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_537 ();
 DECAPx6_ASAP7_75t_R FILLER_280_564 ();
 FILLER_ASAP7_75t_R FILLER_280_578 ();
 DECAPx2_ASAP7_75t_R FILLER_280_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_589 ();
 FILLER_ASAP7_75t_R FILLER_280_596 ();
 DECAPx4_ASAP7_75t_R FILLER_280_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_617 ();
 DECAPx6_ASAP7_75t_R FILLER_280_624 ();
 DECAPx2_ASAP7_75t_R FILLER_280_638 ();
 FILLER_ASAP7_75t_R FILLER_280_677 ();
 DECAPx6_ASAP7_75t_R FILLER_280_685 ();
 FILLER_ASAP7_75t_R FILLER_280_699 ();
 DECAPx1_ASAP7_75t_R FILLER_280_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_739 ();
 FILLER_ASAP7_75t_R FILLER_280_743 ();
 DECAPx6_ASAP7_75t_R FILLER_280_780 ();
 DECAPx2_ASAP7_75t_R FILLER_280_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_820 ();
 DECAPx2_ASAP7_75t_R FILLER_280_834 ();
 FILLERxp5_ASAP7_75t_R FILLER_280_840 ();
 DECAPx2_ASAP7_75t_R FILLER_280_844 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_280_850 ();
 DECAPx2_ASAP7_75t_R FILLER_280_856 ();
 FILLER_ASAP7_75t_R FILLER_280_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_280_926 ();
 DECAPx10_ASAP7_75t_R FILLER_281_2 ();
 DECAPx10_ASAP7_75t_R FILLER_281_24 ();
 DECAPx10_ASAP7_75t_R FILLER_281_46 ();
 DECAPx2_ASAP7_75t_R FILLER_281_68 ();
 FILLER_ASAP7_75t_R FILLER_281_74 ();
 DECAPx10_ASAP7_75t_R FILLER_281_85 ();
 DECAPx2_ASAP7_75t_R FILLER_281_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_113 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_281_123 ();
 FILLER_ASAP7_75t_R FILLER_281_137 ();
 DECAPx1_ASAP7_75t_R FILLER_281_177 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_281_187 ();
 DECAPx1_ASAP7_75t_R FILLER_281_209 ();
 DECAPx2_ASAP7_75t_R FILLER_281_245 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_281_264 ();
 DECAPx10_ASAP7_75t_R FILLER_281_270 ();
 DECAPx4_ASAP7_75t_R FILLER_281_292 ();
 FILLER_ASAP7_75t_R FILLER_281_302 ();
 DECAPx2_ASAP7_75t_R FILLER_281_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_318 ();
 FILLER_ASAP7_75t_R FILLER_281_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_355 ();
 DECAPx6_ASAP7_75t_R FILLER_281_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_389 ();
 DECAPx10_ASAP7_75t_R FILLER_281_398 ();
 DECAPx4_ASAP7_75t_R FILLER_281_420 ();
 FILLER_ASAP7_75t_R FILLER_281_430 ();
 DECAPx2_ASAP7_75t_R FILLER_281_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_444 ();
 FILLER_ASAP7_75t_R FILLER_281_451 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_281_462 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_488 ();
 DECAPx1_ASAP7_75t_R FILLER_281_503 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_507 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_522 ();
 FILLER_ASAP7_75t_R FILLER_281_537 ();
 DECAPx2_ASAP7_75t_R FILLER_281_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_570 ();
 DECAPx2_ASAP7_75t_R FILLER_281_593 ();
 DECAPx1_ASAP7_75t_R FILLER_281_658 ();
 FILLER_ASAP7_75t_R FILLER_281_673 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_691 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_281_700 ();
 DECAPx4_ASAP7_75t_R FILLER_281_710 ();
 DECAPx2_ASAP7_75t_R FILLER_281_726 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_732 ();
 DECAPx4_ASAP7_75t_R FILLER_281_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_281_749 ();
 DECAPx1_ASAP7_75t_R FILLER_281_758 ();
 DECAPx2_ASAP7_75t_R FILLER_281_776 ();
 FILLER_ASAP7_75t_R FILLER_281_782 ();
 DECAPx10_ASAP7_75t_R FILLER_281_792 ();
 DECAPx10_ASAP7_75t_R FILLER_281_814 ();
 DECAPx10_ASAP7_75t_R FILLER_281_836 ();
 DECAPx6_ASAP7_75t_R FILLER_281_858 ();
 DECAPx1_ASAP7_75t_R FILLER_281_872 ();
 FILLER_ASAP7_75t_R FILLER_281_879 ();
 DECAPx2_ASAP7_75t_R FILLER_281_884 ();
 FILLER_ASAP7_75t_R FILLER_281_890 ();
 FILLER_ASAP7_75t_R FILLER_281_898 ();
 DECAPx2_ASAP7_75t_R FILLER_281_903 ();
 FILLER_ASAP7_75t_R FILLER_281_927 ();
 DECAPx10_ASAP7_75t_R FILLER_282_2 ();
 DECAPx10_ASAP7_75t_R FILLER_282_24 ();
 DECAPx10_ASAP7_75t_R FILLER_282_46 ();
 DECAPx10_ASAP7_75t_R FILLER_282_68 ();
 DECAPx10_ASAP7_75t_R FILLER_282_90 ();
 DECAPx6_ASAP7_75t_R FILLER_282_112 ();
 DECAPx2_ASAP7_75t_R FILLER_282_126 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_132 ();
 DECAPx2_ASAP7_75t_R FILLER_282_139 ();
 DECAPx1_ASAP7_75t_R FILLER_282_151 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_282_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_233 ();
 DECAPx1_ASAP7_75t_R FILLER_282_237 ();
 DECAPx10_ASAP7_75t_R FILLER_282_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_282_298 ();
 DECAPx2_ASAP7_75t_R FILLER_282_307 ();
 FILLER_ASAP7_75t_R FILLER_282_313 ();
 DECAPx6_ASAP7_75t_R FILLER_282_323 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_337 ();
 DECAPx1_ASAP7_75t_R FILLER_282_341 ();
 DECAPx1_ASAP7_75t_R FILLER_282_371 ();
 DECAPx6_ASAP7_75t_R FILLER_282_383 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_397 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_405 ();
 DECAPx4_ASAP7_75t_R FILLER_282_418 ();
 DECAPx4_ASAP7_75t_R FILLER_282_451 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_461 ();
 DECAPx2_ASAP7_75t_R FILLER_282_467 ();
 FILLER_ASAP7_75t_R FILLER_282_473 ();
 DECAPx10_ASAP7_75t_R FILLER_282_484 ();
 FILLER_ASAP7_75t_R FILLER_282_506 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_514 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_282_518 ();
 DECAPx6_ASAP7_75t_R FILLER_282_530 ();
 DECAPx1_ASAP7_75t_R FILLER_282_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_548 ();
 FILLER_ASAP7_75t_R FILLER_282_556 ();
 DECAPx1_ASAP7_75t_R FILLER_282_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_572 ();
 DECAPx1_ASAP7_75t_R FILLER_282_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_603 ();
 DECAPx1_ASAP7_75t_R FILLER_282_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_282_628 ();
 DECAPx2_ASAP7_75t_R FILLER_282_656 ();
 FILLER_ASAP7_75t_R FILLER_282_697 ();
 DECAPx6_ASAP7_75t_R FILLER_282_714 ();
 DECAPx2_ASAP7_75t_R FILLER_282_728 ();
 DECAPx10_ASAP7_75t_R FILLER_282_740 ();
 DECAPx6_ASAP7_75t_R FILLER_282_762 ();
 FILLER_ASAP7_75t_R FILLER_282_776 ();
 DECAPx1_ASAP7_75t_R FILLER_282_781 ();
 DECAPx6_ASAP7_75t_R FILLER_282_802 ();
 DECAPx10_ASAP7_75t_R FILLER_282_826 ();
 DECAPx10_ASAP7_75t_R FILLER_282_848 ();
 DECAPx10_ASAP7_75t_R FILLER_282_870 ();
 DECAPx10_ASAP7_75t_R FILLER_282_892 ();
 DECAPx2_ASAP7_75t_R FILLER_282_914 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_282_920 ();
 FILLER_ASAP7_75t_R FILLER_282_932 ();
 DECAPx10_ASAP7_75t_R FILLER_283_2 ();
 DECAPx10_ASAP7_75t_R FILLER_283_24 ();
 DECAPx10_ASAP7_75t_R FILLER_283_46 ();
 DECAPx4_ASAP7_75t_R FILLER_283_68 ();
 FILLER_ASAP7_75t_R FILLER_283_78 ();
 DECAPx10_ASAP7_75t_R FILLER_283_114 ();
 DECAPx4_ASAP7_75t_R FILLER_283_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_146 ();
 DECAPx1_ASAP7_75t_R FILLER_283_161 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_171 ();
 DECAPx1_ASAP7_75t_R FILLER_283_178 ();
 DECAPx2_ASAP7_75t_R FILLER_283_185 ();
 FILLER_ASAP7_75t_R FILLER_283_191 ();
 FILLER_ASAP7_75t_R FILLER_283_205 ();
 DECAPx4_ASAP7_75t_R FILLER_283_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_249 ();
 DECAPx1_ASAP7_75t_R FILLER_283_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_269 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_296 ();
 FILLER_ASAP7_75t_R FILLER_283_311 ();
 DECAPx10_ASAP7_75t_R FILLER_283_319 ();
 DECAPx4_ASAP7_75t_R FILLER_283_341 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_283_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_283_363 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_380 ();
 DECAPx6_ASAP7_75t_R FILLER_283_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_409 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_283_424 ();
 DECAPx10_ASAP7_75t_R FILLER_283_442 ();
 DECAPx10_ASAP7_75t_R FILLER_283_464 ();
 DECAPx1_ASAP7_75t_R FILLER_283_486 ();
 DECAPx6_ASAP7_75t_R FILLER_283_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_527 ();
 DECAPx6_ASAP7_75t_R FILLER_283_534 ();
 FILLER_ASAP7_75t_R FILLER_283_548 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_283_561 ();
 DECAPx10_ASAP7_75t_R FILLER_283_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_618 ();
 DECAPx6_ASAP7_75t_R FILLER_283_632 ();
 FILLER_ASAP7_75t_R FILLER_283_646 ();
 DECAPx10_ASAP7_75t_R FILLER_283_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_680 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_283_691 ();
 DECAPx1_ASAP7_75t_R FILLER_283_700 ();
 DECAPx10_ASAP7_75t_R FILLER_283_710 ();
 DECAPx1_ASAP7_75t_R FILLER_283_732 ();
 DECAPx6_ASAP7_75t_R FILLER_283_742 ();
 DECAPx2_ASAP7_75t_R FILLER_283_756 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_762 ();
 FILLER_ASAP7_75t_R FILLER_283_778 ();
 FILLER_ASAP7_75t_R FILLER_283_786 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_791 ();
 FILLER_ASAP7_75t_R FILLER_283_800 ();
 DECAPx2_ASAP7_75t_R FILLER_283_805 ();
 FILLER_ASAP7_75t_R FILLER_283_811 ();
 DECAPx6_ASAP7_75t_R FILLER_283_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_283_835 ();
 DECAPx2_ASAP7_75t_R FILLER_283_850 ();
 DECAPx4_ASAP7_75t_R FILLER_283_864 ();
 DECAPx10_ASAP7_75t_R FILLER_283_877 ();
 DECAPx10_ASAP7_75t_R FILLER_283_899 ();
 DECAPx1_ASAP7_75t_R FILLER_283_921 ();
 FILLER_ASAP7_75t_R FILLER_283_927 ();
 DECAPx10_ASAP7_75t_R FILLER_284_2 ();
 DECAPx10_ASAP7_75t_R FILLER_284_24 ();
 DECAPx10_ASAP7_75t_R FILLER_284_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_95 ();
 DECAPx4_ASAP7_75t_R FILLER_284_102 ();
 DECAPx2_ASAP7_75t_R FILLER_284_118 ();
 DECAPx4_ASAP7_75t_R FILLER_284_132 ();
 FILLER_ASAP7_75t_R FILLER_284_142 ();
 DECAPx10_ASAP7_75t_R FILLER_284_152 ();
 DECAPx4_ASAP7_75t_R FILLER_284_174 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_190 ();
 DECAPx4_ASAP7_75t_R FILLER_284_197 ();
 FILLER_ASAP7_75t_R FILLER_284_207 ();
 DECAPx10_ASAP7_75t_R FILLER_284_215 ();
 DECAPx10_ASAP7_75t_R FILLER_284_237 ();
 DECAPx6_ASAP7_75t_R FILLER_284_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_273 ();
 FILLER_ASAP7_75t_R FILLER_284_312 ();
 DECAPx2_ASAP7_75t_R FILLER_284_320 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_284_326 ();
 DECAPx10_ASAP7_75t_R FILLER_284_335 ();
 DECAPx10_ASAP7_75t_R FILLER_284_357 ();
 DECAPx1_ASAP7_75t_R FILLER_284_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_383 ();
 DECAPx1_ASAP7_75t_R FILLER_284_396 ();
 DECAPx10_ASAP7_75t_R FILLER_284_428 ();
 DECAPx2_ASAP7_75t_R FILLER_284_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_456 ();
 FILLER_ASAP7_75t_R FILLER_284_460 ();
 DECAPx1_ASAP7_75t_R FILLER_284_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_468 ();
 DECAPx4_ASAP7_75t_R FILLER_284_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_284_496 ();
 DECAPx10_ASAP7_75t_R FILLER_284_508 ();
 DECAPx10_ASAP7_75t_R FILLER_284_530 ();
 DECAPx4_ASAP7_75t_R FILLER_284_552 ();
 FILLER_ASAP7_75t_R FILLER_284_562 ();
 DECAPx1_ASAP7_75t_R FILLER_284_574 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_578 ();
 DECAPx1_ASAP7_75t_R FILLER_284_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_586 ();
 DECAPx10_ASAP7_75t_R FILLER_284_590 ();
 DECAPx10_ASAP7_75t_R FILLER_284_612 ();
 DECAPx6_ASAP7_75t_R FILLER_284_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_648 ();
 DECAPx10_ASAP7_75t_R FILLER_284_659 ();
 DECAPx2_ASAP7_75t_R FILLER_284_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_697 ();
 DECAPx6_ASAP7_75t_R FILLER_284_718 ();
 DECAPx1_ASAP7_75t_R FILLER_284_732 ();
 DECAPx10_ASAP7_75t_R FILLER_284_743 ();
 DECAPx4_ASAP7_75t_R FILLER_284_765 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_284_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_284_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_787 ();
 FILLER_ASAP7_75t_R FILLER_284_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_836 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_854 ();
 DECAPx2_ASAP7_75t_R FILLER_284_864 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_870 ();
 DECAPx1_ASAP7_75t_R FILLER_284_888 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_892 ();
 DECAPx1_ASAP7_75t_R FILLER_284_903 ();
 FILLERxp5_ASAP7_75t_R FILLER_284_907 ();
 DECAPx10_ASAP7_75t_R FILLER_285_2 ();
 DECAPx10_ASAP7_75t_R FILLER_285_24 ();
 DECAPx10_ASAP7_75t_R FILLER_285_46 ();
 DECAPx6_ASAP7_75t_R FILLER_285_68 ();
 FILLER_ASAP7_75t_R FILLER_285_82 ();
 DECAPx1_ASAP7_75t_R FILLER_285_87 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_91 ();
 DECAPx2_ASAP7_75t_R FILLER_285_95 ();
 DECAPx2_ASAP7_75t_R FILLER_285_133 ();
 FILLER_ASAP7_75t_R FILLER_285_139 ();
 DECAPx2_ASAP7_75t_R FILLER_285_147 ();
 DECAPx6_ASAP7_75t_R FILLER_285_159 ();
 DECAPx1_ASAP7_75t_R FILLER_285_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_177 ();
 DECAPx10_ASAP7_75t_R FILLER_285_204 ();
 DECAPx4_ASAP7_75t_R FILLER_285_226 ();
 DECAPx6_ASAP7_75t_R FILLER_285_242 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_285_256 ();
 DECAPx4_ASAP7_75t_R FILLER_285_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_275 ();
 DECAPx2_ASAP7_75t_R FILLER_285_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_285_321 ();
 DECAPx2_ASAP7_75t_R FILLER_285_350 ();
 FILLER_ASAP7_75t_R FILLER_285_356 ();
 DECAPx4_ASAP7_75t_R FILLER_285_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_378 ();
 DECAPx10_ASAP7_75t_R FILLER_285_405 ();
 DECAPx10_ASAP7_75t_R FILLER_285_427 ();
 DECAPx1_ASAP7_75t_R FILLER_285_479 ();
 DECAPx10_ASAP7_75t_R FILLER_285_486 ();
 DECAPx6_ASAP7_75t_R FILLER_285_508 ();
 DECAPx1_ASAP7_75t_R FILLER_285_522 ();
 DECAPx2_ASAP7_75t_R FILLER_285_540 ();
 FILLER_ASAP7_75t_R FILLER_285_546 ();
 DECAPx10_ASAP7_75t_R FILLER_285_554 ();
 DECAPx10_ASAP7_75t_R FILLER_285_576 ();
 DECAPx4_ASAP7_75t_R FILLER_285_598 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_285_608 ();
 DECAPx1_ASAP7_75t_R FILLER_285_615 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_619 ();
 DECAPx6_ASAP7_75t_R FILLER_285_626 ();
 DECAPx2_ASAP7_75t_R FILLER_285_660 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_285_666 ();
 DECAPx6_ASAP7_75t_R FILLER_285_675 ();
 DECAPx1_ASAP7_75t_R FILLER_285_689 ();
 DECAPx2_ASAP7_75t_R FILLER_285_710 ();
 FILLER_ASAP7_75t_R FILLER_285_716 ();
 FILLER_ASAP7_75t_R FILLER_285_732 ();
 DECAPx2_ASAP7_75t_R FILLER_285_770 ();
 FILLER_ASAP7_75t_R FILLER_285_776 ();
 DECAPx10_ASAP7_75t_R FILLER_285_790 ();
 DECAPx2_ASAP7_75t_R FILLER_285_812 ();
 FILLER_ASAP7_75t_R FILLER_285_818 ();
 DECAPx1_ASAP7_75t_R FILLER_285_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_285_924 ();
 DECAPx1_ASAP7_75t_R FILLER_285_930 ();
 DECAPx10_ASAP7_75t_R FILLER_286_2 ();
 DECAPx10_ASAP7_75t_R FILLER_286_24 ();
 DECAPx10_ASAP7_75t_R FILLER_286_46 ();
 DECAPx2_ASAP7_75t_R FILLER_286_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_74 ();
 DECAPx6_ASAP7_75t_R FILLER_286_89 ();
 DECAPx1_ASAP7_75t_R FILLER_286_103 ();
 FILLER_ASAP7_75t_R FILLER_286_113 ();
 DECAPx1_ASAP7_75t_R FILLER_286_118 ();
 FILLER_ASAP7_75t_R FILLER_286_125 ();
 FILLER_ASAP7_75t_R FILLER_286_130 ();
 DECAPx6_ASAP7_75t_R FILLER_286_146 ();
 DECAPx2_ASAP7_75t_R FILLER_286_160 ();
 DECAPx6_ASAP7_75t_R FILLER_286_172 ();
 DECAPx2_ASAP7_75t_R FILLER_286_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_192 ();
 DECAPx2_ASAP7_75t_R FILLER_286_196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_202 ();
 DECAPx1_ASAP7_75t_R FILLER_286_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_246 ();
 DECAPx2_ASAP7_75t_R FILLER_286_275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_281 ();
 DECAPx2_ASAP7_75t_R FILLER_286_287 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_293 ();
 DECAPx6_ASAP7_75t_R FILLER_286_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_311 ();
 DECAPx1_ASAP7_75t_R FILLER_286_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_338 ();
 DECAPx1_ASAP7_75t_R FILLER_286_359 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_363 ();
 DECAPx6_ASAP7_75t_R FILLER_286_379 ();
 DECAPx10_ASAP7_75t_R FILLER_286_396 ();
 DECAPx10_ASAP7_75t_R FILLER_286_418 ();
 DECAPx2_ASAP7_75t_R FILLER_286_440 ();
 FILLER_ASAP7_75t_R FILLER_286_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_464 ();
 DECAPx2_ASAP7_75t_R FILLER_286_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_485 ();
 DECAPx6_ASAP7_75t_R FILLER_286_505 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_519 ();
 DECAPx10_ASAP7_75t_R FILLER_286_571 ();
 DECAPx1_ASAP7_75t_R FILLER_286_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_605 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_620 ();
 DECAPx6_ASAP7_75t_R FILLER_286_636 ();
 DECAPx2_ASAP7_75t_R FILLER_286_650 ();
 FILLER_ASAP7_75t_R FILLER_286_663 ();
 DECAPx2_ASAP7_75t_R FILLER_286_678 ();
 FILLER_ASAP7_75t_R FILLER_286_684 ();
 DECAPx6_ASAP7_75t_R FILLER_286_696 ();
 FILLER_ASAP7_75t_R FILLER_286_710 ();
 DECAPx1_ASAP7_75t_R FILLER_286_737 ();
 DECAPx6_ASAP7_75t_R FILLER_286_780 ();
 DECAPx2_ASAP7_75t_R FILLER_286_794 ();
 DECAPx6_ASAP7_75t_R FILLER_286_806 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_824 ();
 DECAPx2_ASAP7_75t_R FILLER_286_832 ();
 FILLER_ASAP7_75t_R FILLER_286_838 ();
 DECAPx1_ASAP7_75t_R FILLER_286_843 ();
 DECAPx4_ASAP7_75t_R FILLER_286_853 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_286_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_286_875 ();
 FILLER_ASAP7_75t_R FILLER_286_884 ();
 DECAPx2_ASAP7_75t_R FILLER_286_905 ();
 DECAPx6_ASAP7_75t_R FILLER_286_920 ();
 DECAPx10_ASAP7_75t_R FILLER_287_2 ();
 DECAPx10_ASAP7_75t_R FILLER_287_24 ();
 DECAPx10_ASAP7_75t_R FILLER_287_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_68 ();
 DECAPx4_ASAP7_75t_R FILLER_287_97 ();
 DECAPx10_ASAP7_75t_R FILLER_287_119 ();
 DECAPx1_ASAP7_75t_R FILLER_287_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_151 ();
 FILLER_ASAP7_75t_R FILLER_287_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_183 ();
 FILLER_ASAP7_75t_R FILLER_287_192 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_211 ();
 DECAPx4_ASAP7_75t_R FILLER_287_240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_250 ();
 DECAPx1_ASAP7_75t_R FILLER_287_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_263 ();
 DECAPx10_ASAP7_75t_R FILLER_287_267 ();
 DECAPx6_ASAP7_75t_R FILLER_287_289 ();
 DECAPx1_ASAP7_75t_R FILLER_287_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_307 ();
 FILLER_ASAP7_75t_R FILLER_287_314 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_319 ();
 DECAPx6_ASAP7_75t_R FILLER_287_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_337 ();
 DECAPx4_ASAP7_75t_R FILLER_287_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_353 ();
 DECAPx2_ASAP7_75t_R FILLER_287_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_386 ();
 DECAPx6_ASAP7_75t_R FILLER_287_395 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_409 ();
 FILLER_ASAP7_75t_R FILLER_287_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_482 ();
 FILLER_ASAP7_75t_R FILLER_287_509 ();
 DECAPx2_ASAP7_75t_R FILLER_287_526 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_532 ();
 FILLER_ASAP7_75t_R FILLER_287_538 ();
 DECAPx2_ASAP7_75t_R FILLER_287_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_549 ();
 DECAPx6_ASAP7_75t_R FILLER_287_555 ();
 DECAPx1_ASAP7_75t_R FILLER_287_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_583 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_596 ();
 DECAPx1_ASAP7_75t_R FILLER_287_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_610 ();
 DECAPx2_ASAP7_75t_R FILLER_287_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_623 ();
 DECAPx10_ASAP7_75t_R FILLER_287_634 ();
 DECAPx6_ASAP7_75t_R FILLER_287_656 ();
 DECAPx2_ASAP7_75t_R FILLER_287_670 ();
 DECAPx10_ASAP7_75t_R FILLER_287_682 ();
 DECAPx4_ASAP7_75t_R FILLER_287_704 ();
 DECAPx6_ASAP7_75t_R FILLER_287_743 ();
 DECAPx1_ASAP7_75t_R FILLER_287_757 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_761 ();
 DECAPx10_ASAP7_75t_R FILLER_287_772 ();
 DECAPx1_ASAP7_75t_R FILLER_287_794 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_825 ();
 DECAPx10_ASAP7_75t_R FILLER_287_852 ();
 DECAPx10_ASAP7_75t_R FILLER_287_874 ();
 DECAPx4_ASAP7_75t_R FILLER_287_896 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_287_906 ();
 DECAPx1_ASAP7_75t_R FILLER_287_921 ();
 DECAPx2_ASAP7_75t_R FILLER_287_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_287_933 ();
 DECAPx10_ASAP7_75t_R FILLER_288_2 ();
 DECAPx10_ASAP7_75t_R FILLER_288_24 ();
 DECAPx10_ASAP7_75t_R FILLER_288_46 ();
 DECAPx6_ASAP7_75t_R FILLER_288_68 ();
 DECAPx1_ASAP7_75t_R FILLER_288_82 ();
 DECAPx4_ASAP7_75t_R FILLER_288_89 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_99 ();
 DECAPx2_ASAP7_75t_R FILLER_288_128 ();
 FILLER_ASAP7_75t_R FILLER_288_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_168 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_174 ();
 DECAPx2_ASAP7_75t_R FILLER_288_201 ();
 DECAPx2_ASAP7_75t_R FILLER_288_213 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_228 ();
 DECAPx6_ASAP7_75t_R FILLER_288_232 ();
 FILLER_ASAP7_75t_R FILLER_288_246 ();
 DECAPx2_ASAP7_75t_R FILLER_288_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_260 ();
 DECAPx6_ASAP7_75t_R FILLER_288_267 ();
 DECAPx1_ASAP7_75t_R FILLER_288_281 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_291 ();
 FILLER_ASAP7_75t_R FILLER_288_300 ();
 DECAPx10_ASAP7_75t_R FILLER_288_328 ();
 DECAPx4_ASAP7_75t_R FILLER_288_350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_360 ();
 DECAPx2_ASAP7_75t_R FILLER_288_372 ();
 FILLER_ASAP7_75t_R FILLER_288_407 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_417 ();
 FILLER_ASAP7_75t_R FILLER_288_460 ();
 DECAPx1_ASAP7_75t_R FILLER_288_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_468 ();
 DECAPx1_ASAP7_75t_R FILLER_288_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_487 ();
 DECAPx1_ASAP7_75t_R FILLER_288_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_532 ();
 DECAPx4_ASAP7_75t_R FILLER_288_536 ();
 FILLER_ASAP7_75t_R FILLER_288_546 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_568 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_288_591 ();
 DECAPx1_ASAP7_75t_R FILLER_288_601 ();
 DECAPx2_ASAP7_75t_R FILLER_288_613 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_619 ();
 DECAPx2_ASAP7_75t_R FILLER_288_630 ();
 FILLER_ASAP7_75t_R FILLER_288_646 ();
 DECAPx10_ASAP7_75t_R FILLER_288_651 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_673 ();
 FILLER_ASAP7_75t_R FILLER_288_690 ();
 DECAPx10_ASAP7_75t_R FILLER_288_698 ();
 DECAPx4_ASAP7_75t_R FILLER_288_720 ();
 DECAPx2_ASAP7_75t_R FILLER_288_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_288_745 ();
 DECAPx10_ASAP7_75t_R FILLER_288_755 ();
 DECAPx2_ASAP7_75t_R FILLER_288_777 ();
 DECAPx1_ASAP7_75t_R FILLER_288_791 ();
 DECAPx10_ASAP7_75t_R FILLER_288_821 ();
 DECAPx10_ASAP7_75t_R FILLER_288_843 ();
 DECAPx1_ASAP7_75t_R FILLER_288_865 ();
 DECAPx10_ASAP7_75t_R FILLER_288_872 ();
 DECAPx10_ASAP7_75t_R FILLER_288_894 ();
 DECAPx6_ASAP7_75t_R FILLER_288_916 ();
 DECAPx1_ASAP7_75t_R FILLER_288_930 ();
 DECAPx10_ASAP7_75t_R FILLER_289_2 ();
 DECAPx10_ASAP7_75t_R FILLER_289_24 ();
 DECAPx10_ASAP7_75t_R FILLER_289_46 ();
 DECAPx1_ASAP7_75t_R FILLER_289_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_72 ();
 DECAPx6_ASAP7_75t_R FILLER_289_99 ();
 DECAPx1_ASAP7_75t_R FILLER_289_113 ();
 DECAPx6_ASAP7_75t_R FILLER_289_120 ();
 DECAPx1_ASAP7_75t_R FILLER_289_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_138 ();
 DECAPx2_ASAP7_75t_R FILLER_289_145 ();
 DECAPx10_ASAP7_75t_R FILLER_289_154 ();
 DECAPx1_ASAP7_75t_R FILLER_289_176 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_289_186 ();
 DECAPx10_ASAP7_75t_R FILLER_289_192 ();
 DECAPx2_ASAP7_75t_R FILLER_289_214 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_289_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_285 ();
 DECAPx4_ASAP7_75t_R FILLER_289_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_304 ();
 DECAPx6_ASAP7_75t_R FILLER_289_311 ();
 DECAPx2_ASAP7_75t_R FILLER_289_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_337 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_352 ();
 DECAPx1_ASAP7_75t_R FILLER_289_379 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_383 ();
 FILLER_ASAP7_75t_R FILLER_289_390 ();
 DECAPx1_ASAP7_75t_R FILLER_289_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_405 ();
 DECAPx1_ASAP7_75t_R FILLER_289_413 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_417 ();
 DECAPx1_ASAP7_75t_R FILLER_289_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_461 ();
 FILLER_ASAP7_75t_R FILLER_289_476 ();
 DECAPx4_ASAP7_75t_R FILLER_289_484 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_289_494 ();
 DECAPx2_ASAP7_75t_R FILLER_289_500 ();
 FILLER_ASAP7_75t_R FILLER_289_506 ();
 FILLER_ASAP7_75t_R FILLER_289_514 ();
 DECAPx10_ASAP7_75t_R FILLER_289_519 ();
 DECAPx6_ASAP7_75t_R FILLER_289_541 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_289_555 ();
 DECAPx6_ASAP7_75t_R FILLER_289_573 ();
 FILLER_ASAP7_75t_R FILLER_289_587 ();
 DECAPx10_ASAP7_75t_R FILLER_289_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_618 ();
 FILLER_ASAP7_75t_R FILLER_289_629 ();
 FILLER_ASAP7_75t_R FILLER_289_668 ();
 DECAPx4_ASAP7_75t_R FILLER_289_688 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_698 ();
 DECAPx10_ASAP7_75t_R FILLER_289_717 ();
 DECAPx6_ASAP7_75t_R FILLER_289_739 ();
 DECAPx1_ASAP7_75t_R FILLER_289_753 ();
 DECAPx10_ASAP7_75t_R FILLER_289_819 ();
 DECAPx6_ASAP7_75t_R FILLER_289_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_289_855 ();
 DECAPx2_ASAP7_75t_R FILLER_289_873 ();
 FILLER_ASAP7_75t_R FILLER_289_879 ();
 DECAPx6_ASAP7_75t_R FILLER_289_884 ();
 FILLER_ASAP7_75t_R FILLER_289_898 ();
 DECAPx6_ASAP7_75t_R FILLER_289_909 ();
 FILLER_ASAP7_75t_R FILLER_289_923 ();
 DECAPx2_ASAP7_75t_R FILLER_289_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_289_933 ();
 DECAPx10_ASAP7_75t_R FILLER_290_2 ();
 DECAPx10_ASAP7_75t_R FILLER_290_24 ();
 DECAPx10_ASAP7_75t_R FILLER_290_46 ();
 DECAPx4_ASAP7_75t_R FILLER_290_68 ();
 FILLER_ASAP7_75t_R FILLER_290_78 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_86 ();
 FILLER_ASAP7_75t_R FILLER_290_93 ();
 DECAPx1_ASAP7_75t_R FILLER_290_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_128 ();
 DECAPx10_ASAP7_75t_R FILLER_290_138 ();
 DECAPx1_ASAP7_75t_R FILLER_290_160 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_164 ();
 DECAPx6_ASAP7_75t_R FILLER_290_177 ();
 DECAPx1_ASAP7_75t_R FILLER_290_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_195 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_290_202 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_211 ();
 DECAPx2_ASAP7_75t_R FILLER_290_238 ();
 DECAPx1_ASAP7_75t_R FILLER_290_269 ();
 DECAPx1_ASAP7_75t_R FILLER_290_305 ();
 DECAPx1_ASAP7_75t_R FILLER_290_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_321 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_357 ();
 DECAPx1_ASAP7_75t_R FILLER_290_364 ();
 DECAPx10_ASAP7_75t_R FILLER_290_371 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_290_393 ();
 FILLER_ASAP7_75t_R FILLER_290_404 ();
 DECAPx10_ASAP7_75t_R FILLER_290_432 ();
 DECAPx2_ASAP7_75t_R FILLER_290_454 ();
 FILLER_ASAP7_75t_R FILLER_290_460 ();
 DECAPx2_ASAP7_75t_R FILLER_290_464 ();
 FILLER_ASAP7_75t_R FILLER_290_470 ();
 DECAPx10_ASAP7_75t_R FILLER_290_478 ();
 DECAPx6_ASAP7_75t_R FILLER_290_500 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_290_514 ();
 DECAPx2_ASAP7_75t_R FILLER_290_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_532 ();
 DECAPx6_ASAP7_75t_R FILLER_290_542 ();
 DECAPx1_ASAP7_75t_R FILLER_290_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_560 ();
 DECAPx10_ASAP7_75t_R FILLER_290_564 ();
 DECAPx1_ASAP7_75t_R FILLER_290_586 ();
 DECAPx10_ASAP7_75t_R FILLER_290_609 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_631 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_638 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_662 ();
 DECAPx2_ASAP7_75t_R FILLER_290_687 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_693 ();
 DECAPx10_ASAP7_75t_R FILLER_290_713 ();
 DECAPx1_ASAP7_75t_R FILLER_290_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_739 ();
 DECAPx10_ASAP7_75t_R FILLER_290_746 ();
 DECAPx1_ASAP7_75t_R FILLER_290_768 ();
 DECAPx2_ASAP7_75t_R FILLER_290_775 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_781 ();
 DECAPx10_ASAP7_75t_R FILLER_290_793 ();
 DECAPx10_ASAP7_75t_R FILLER_290_815 ();
 DECAPx2_ASAP7_75t_R FILLER_290_837 ();
 FILLERxp5_ASAP7_75t_R FILLER_290_843 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_290_856 ();
 FILLER_ASAP7_75t_R FILLER_290_893 ();
 FILLER_ASAP7_75t_R FILLER_290_904 ();
 FILLER_ASAP7_75t_R FILLER_290_932 ();
 DECAPx10_ASAP7_75t_R FILLER_291_2 ();
 DECAPx10_ASAP7_75t_R FILLER_291_24 ();
 DECAPx10_ASAP7_75t_R FILLER_291_46 ();
 DECAPx6_ASAP7_75t_R FILLER_291_68 ();
 DECAPx1_ASAP7_75t_R FILLER_291_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_86 ();
 DECAPx6_ASAP7_75t_R FILLER_291_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_104 ();
 DECAPx2_ASAP7_75t_R FILLER_291_113 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_119 ();
 DECAPx2_ASAP7_75t_R FILLER_291_146 ();
 DECAPx2_ASAP7_75t_R FILLER_291_178 ();
 FILLER_ASAP7_75t_R FILLER_291_184 ();
 FILLER_ASAP7_75t_R FILLER_291_224 ();
 DECAPx2_ASAP7_75t_R FILLER_291_229 ();
 DECAPx4_ASAP7_75t_R FILLER_291_241 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_251 ();
 DECAPx2_ASAP7_75t_R FILLER_291_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_263 ();
 DECAPx1_ASAP7_75t_R FILLER_291_272 ();
 FILLER_ASAP7_75t_R FILLER_291_282 ();
 FILLER_ASAP7_75t_R FILLER_291_290 ();
 DECAPx1_ASAP7_75t_R FILLER_291_298 ();
 DECAPx6_ASAP7_75t_R FILLER_291_355 ();
 DECAPx2_ASAP7_75t_R FILLER_291_369 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_375 ();
 DECAPx4_ASAP7_75t_R FILLER_291_391 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_401 ();
 DECAPx1_ASAP7_75t_R FILLER_291_412 ();
 DECAPx2_ASAP7_75t_R FILLER_291_425 ();
 DECAPx6_ASAP7_75t_R FILLER_291_438 ();
 DECAPx1_ASAP7_75t_R FILLER_291_452 ();
 DECAPx10_ASAP7_75t_R FILLER_291_459 ();
 DECAPx6_ASAP7_75t_R FILLER_291_481 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_495 ();
 DECAPx4_ASAP7_75t_R FILLER_291_504 ();
 DECAPx2_ASAP7_75t_R FILLER_291_528 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_534 ();
 DECAPx6_ASAP7_75t_R FILLER_291_540 ();
 DECAPx2_ASAP7_75t_R FILLER_291_554 ();
 DECAPx10_ASAP7_75t_R FILLER_291_563 ();
 DECAPx1_ASAP7_75t_R FILLER_291_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_589 ();
 DECAPx10_ASAP7_75t_R FILLER_291_602 ();
 DECAPx10_ASAP7_75t_R FILLER_291_624 ();
 FILLER_ASAP7_75t_R FILLER_291_646 ();
 FILLER_ASAP7_75t_R FILLER_291_654 ();
 DECAPx2_ASAP7_75t_R FILLER_291_674 ();
 FILLER_ASAP7_75t_R FILLER_291_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_688 ();
 DECAPx10_ASAP7_75t_R FILLER_291_699 ();
 DECAPx2_ASAP7_75t_R FILLER_291_721 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_727 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_749 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_760 ();
 DECAPx10_ASAP7_75t_R FILLER_291_773 ();
 DECAPx6_ASAP7_75t_R FILLER_291_795 ();
 DECAPx1_ASAP7_75t_R FILLER_291_809 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_813 ();
 FILLER_ASAP7_75t_R FILLER_291_826 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_291_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_291_924 ();
 DECAPx1_ASAP7_75t_R FILLER_291_930 ();
 DECAPx10_ASAP7_75t_R FILLER_292_2 ();
 DECAPx10_ASAP7_75t_R FILLER_292_24 ();
 DECAPx10_ASAP7_75t_R FILLER_292_46 ();
 DECAPx4_ASAP7_75t_R FILLER_292_68 ();
 DECAPx1_ASAP7_75t_R FILLER_292_90 ();
 DECAPx4_ASAP7_75t_R FILLER_292_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_110 ();
 DECAPx1_ASAP7_75t_R FILLER_292_120 ();
 DECAPx1_ASAP7_75t_R FILLER_292_130 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_134 ();
 DECAPx2_ASAP7_75t_R FILLER_292_141 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_292_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_205 ();
 DECAPx6_ASAP7_75t_R FILLER_292_209 ();
 DECAPx2_ASAP7_75t_R FILLER_292_223 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_229 ();
 DECAPx10_ASAP7_75t_R FILLER_292_256 ();
 DECAPx10_ASAP7_75t_R FILLER_292_278 ();
 DECAPx10_ASAP7_75t_R FILLER_292_300 ();
 DECAPx10_ASAP7_75t_R FILLER_292_322 ();
 DECAPx4_ASAP7_75t_R FILLER_292_344 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_292_354 ();
 DECAPx1_ASAP7_75t_R FILLER_292_363 ();
 DECAPx6_ASAP7_75t_R FILLER_292_394 ();
 DECAPx10_ASAP7_75t_R FILLER_292_414 ();
 DECAPx4_ASAP7_75t_R FILLER_292_436 ();
 FILLER_ASAP7_75t_R FILLER_292_446 ();
 DECAPx6_ASAP7_75t_R FILLER_292_473 ();
 DECAPx2_ASAP7_75t_R FILLER_292_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_493 ();
 DECAPx6_ASAP7_75t_R FILLER_292_517 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_531 ();
 DECAPx2_ASAP7_75t_R FILLER_292_563 ();
 DECAPx1_ASAP7_75t_R FILLER_292_575 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_579 ();
 DECAPx1_ASAP7_75t_R FILLER_292_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_612 ();
 DECAPx4_ASAP7_75t_R FILLER_292_620 ();
 FILLER_ASAP7_75t_R FILLER_292_630 ();
 DECAPx6_ASAP7_75t_R FILLER_292_639 ();
 DECAPx1_ASAP7_75t_R FILLER_292_653 ();
 DECAPx6_ASAP7_75t_R FILLER_292_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_292_677 ();
 DECAPx6_ASAP7_75t_R FILLER_292_703 ();
 DECAPx1_ASAP7_75t_R FILLER_292_717 ();
 DECAPx1_ASAP7_75t_R FILLER_292_764 ();
 DECAPx4_ASAP7_75t_R FILLER_292_787 ();
 FILLER_ASAP7_75t_R FILLER_292_797 ();
 FILLER_ASAP7_75t_R FILLER_292_802 ();
 FILLER_ASAP7_75t_R FILLER_292_837 ();
 DECAPx2_ASAP7_75t_R FILLER_292_865 ();
 DECAPx4_ASAP7_75t_R FILLER_292_897 ();
 FILLERxp5_ASAP7_75t_R FILLER_292_907 ();
 DECAPx10_ASAP7_75t_R FILLER_293_2 ();
 DECAPx10_ASAP7_75t_R FILLER_293_24 ();
 DECAPx10_ASAP7_75t_R FILLER_293_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_68 ();
 DECAPx6_ASAP7_75t_R FILLER_293_113 ();
 DECAPx1_ASAP7_75t_R FILLER_293_127 ();
 FILLER_ASAP7_75t_R FILLER_293_160 ();
 DECAPx6_ASAP7_75t_R FILLER_293_165 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_179 ();
 DECAPx2_ASAP7_75t_R FILLER_293_188 ();
 DECAPx6_ASAP7_75t_R FILLER_293_197 ();
 DECAPx2_ASAP7_75t_R FILLER_293_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_217 ();
 DECAPx6_ASAP7_75t_R FILLER_293_224 ();
 DECAPx1_ASAP7_75t_R FILLER_293_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_251 ();
 DECAPx10_ASAP7_75t_R FILLER_293_255 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_277 ();
 DECAPx2_ASAP7_75t_R FILLER_293_284 ();
 DECAPx2_ASAP7_75t_R FILLER_293_293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_299 ();
 DECAPx10_ASAP7_75t_R FILLER_293_312 ();
 DECAPx6_ASAP7_75t_R FILLER_293_334 ();
 DECAPx1_ASAP7_75t_R FILLER_293_348 ();
 DECAPx10_ASAP7_75t_R FILLER_293_381 ();
 DECAPx10_ASAP7_75t_R FILLER_293_403 ();
 DECAPx6_ASAP7_75t_R FILLER_293_425 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_494 ();
 DECAPx4_ASAP7_75t_R FILLER_293_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_519 ();
 DECAPx1_ASAP7_75t_R FILLER_293_529 ();
 DECAPx2_ASAP7_75t_R FILLER_293_553 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_559 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_565 ();
 DECAPx6_ASAP7_75t_R FILLER_293_584 ();
 DECAPx2_ASAP7_75t_R FILLER_293_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_604 ();
 DECAPx2_ASAP7_75t_R FILLER_293_611 ();
 DECAPx10_ASAP7_75t_R FILLER_293_645 ();
 DECAPx6_ASAP7_75t_R FILLER_293_667 ();
 DECAPx1_ASAP7_75t_R FILLER_293_681 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_685 ();
 DECAPx10_ASAP7_75t_R FILLER_293_692 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_714 ();
 FILLER_ASAP7_75t_R FILLER_293_751 ();
 DECAPx10_ASAP7_75t_R FILLER_293_762 ();
 DECAPx2_ASAP7_75t_R FILLER_293_788 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_794 ();
 DECAPx4_ASAP7_75t_R FILLER_293_804 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_814 ();
 DECAPx4_ASAP7_75t_R FILLER_293_841 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_851 ();
 DECAPx10_ASAP7_75t_R FILLER_293_857 ();
 DECAPx2_ASAP7_75t_R FILLER_293_879 ();
 FILLERxp5_ASAP7_75t_R FILLER_293_885 ();
 DECAPx10_ASAP7_75t_R FILLER_293_889 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_911 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_293_922 ();
 DECAPx1_ASAP7_75t_R FILLER_293_930 ();
 DECAPx10_ASAP7_75t_R FILLER_294_2 ();
 DECAPx10_ASAP7_75t_R FILLER_294_24 ();
 DECAPx10_ASAP7_75t_R FILLER_294_46 ();
 DECAPx6_ASAP7_75t_R FILLER_294_68 ();
 DECAPx1_ASAP7_75t_R FILLER_294_82 ();
 DECAPx2_ASAP7_75t_R FILLER_294_89 ();
 DECAPx10_ASAP7_75t_R FILLER_294_101 ();
 DECAPx6_ASAP7_75t_R FILLER_294_123 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_144 ();
 DECAPx10_ASAP7_75t_R FILLER_294_148 ();
 DECAPx1_ASAP7_75t_R FILLER_294_170 ();
 DECAPx6_ASAP7_75t_R FILLER_294_193 ();
 FILLER_ASAP7_75t_R FILLER_294_207 ();
 DECAPx10_ASAP7_75t_R FILLER_294_235 ();
 DECAPx4_ASAP7_75t_R FILLER_294_257 ();
 FILLER_ASAP7_75t_R FILLER_294_293 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_294_301 ();
 DECAPx4_ASAP7_75t_R FILLER_294_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_329 ();
 DECAPx10_ASAP7_75t_R FILLER_294_336 ();
 DECAPx1_ASAP7_75t_R FILLER_294_358 ();
 DECAPx6_ASAP7_75t_R FILLER_294_371 ();
 DECAPx1_ASAP7_75t_R FILLER_294_385 ();
 DECAPx1_ASAP7_75t_R FILLER_294_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_416 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_294_423 ();
 DECAPx1_ASAP7_75t_R FILLER_294_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_444 ();
 DECAPx2_ASAP7_75t_R FILLER_294_454 ();
 FILLER_ASAP7_75t_R FILLER_294_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_294_470 ();
 DECAPx10_ASAP7_75t_R FILLER_294_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_294_515 ();
 DECAPx6_ASAP7_75t_R FILLER_294_530 ();
 DECAPx1_ASAP7_75t_R FILLER_294_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_548 ();
 DECAPx10_ASAP7_75t_R FILLER_294_575 ();
 DECAPx1_ASAP7_75t_R FILLER_294_597 ();
 DECAPx1_ASAP7_75t_R FILLER_294_615 ();
 DECAPx2_ASAP7_75t_R FILLER_294_626 ();
 DECAPx10_ASAP7_75t_R FILLER_294_639 ();
 DECAPx10_ASAP7_75t_R FILLER_294_661 ();
 DECAPx10_ASAP7_75t_R FILLER_294_683 ();
 DECAPx4_ASAP7_75t_R FILLER_294_705 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_294_715 ();
 DECAPx6_ASAP7_75t_R FILLER_294_740 ();
 DECAPx1_ASAP7_75t_R FILLER_294_754 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_758 ();
 DECAPx4_ASAP7_75t_R FILLER_294_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_772 ();
 DECAPx1_ASAP7_75t_R FILLER_294_776 ();
 FILLER_ASAP7_75t_R FILLER_294_786 ();
 DECAPx4_ASAP7_75t_R FILLER_294_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_294_828 ();
 DECAPx10_ASAP7_75t_R FILLER_294_832 ();
 DECAPx10_ASAP7_75t_R FILLER_294_854 ();
 DECAPx6_ASAP7_75t_R FILLER_294_876 ();
 FILLER_ASAP7_75t_R FILLER_294_890 ();
 DECAPx10_ASAP7_75t_R FILLER_294_900 ();
 DECAPx4_ASAP7_75t_R FILLER_294_922 ();
 FILLER_ASAP7_75t_R FILLER_294_932 ();
 DECAPx10_ASAP7_75t_R FILLER_295_2 ();
 DECAPx10_ASAP7_75t_R FILLER_295_24 ();
 DECAPx10_ASAP7_75t_R FILLER_295_46 ();
 DECAPx2_ASAP7_75t_R FILLER_295_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_74 ();
 DECAPx10_ASAP7_75t_R FILLER_295_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_103 ();
 DECAPx10_ASAP7_75t_R FILLER_295_130 ();
 DECAPx4_ASAP7_75t_R FILLER_295_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_162 ();
 DECAPx1_ASAP7_75t_R FILLER_295_194 ();
 DECAPx4_ASAP7_75t_R FILLER_295_204 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_295_220 ();
 DECAPx6_ASAP7_75t_R FILLER_295_226 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_240 ();
 DECAPx1_ASAP7_75t_R FILLER_295_247 ();
 FILLER_ASAP7_75t_R FILLER_295_271 ();
 FILLER_ASAP7_75t_R FILLER_295_279 ();
 DECAPx2_ASAP7_75t_R FILLER_295_284 ();
 DECAPx1_ASAP7_75t_R FILLER_295_316 ();
 DECAPx10_ASAP7_75t_R FILLER_295_355 ();
 DECAPx1_ASAP7_75t_R FILLER_295_377 ();
 FILLER_ASAP7_75t_R FILLER_295_413 ();
 DECAPx10_ASAP7_75t_R FILLER_295_453 ();
 DECAPx2_ASAP7_75t_R FILLER_295_475 ();
 DECAPx10_ASAP7_75t_R FILLER_295_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_515 ();
 DECAPx10_ASAP7_75t_R FILLER_295_530 ();
 DECAPx10_ASAP7_75t_R FILLER_295_552 ();
 DECAPx2_ASAP7_75t_R FILLER_295_574 ();
 DECAPx2_ASAP7_75t_R FILLER_295_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_592 ();
 DECAPx1_ASAP7_75t_R FILLER_295_599 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_610 ();
 DECAPx10_ASAP7_75t_R FILLER_295_614 ();
 DECAPx4_ASAP7_75t_R FILLER_295_636 ();
 DECAPx10_ASAP7_75t_R FILLER_295_652 ();
 DECAPx10_ASAP7_75t_R FILLER_295_674 ();
 DECAPx10_ASAP7_75t_R FILLER_295_696 ();
 DECAPx10_ASAP7_75t_R FILLER_295_718 ();
 DECAPx6_ASAP7_75t_R FILLER_295_740 ();
 DECAPx2_ASAP7_75t_R FILLER_295_754 ();
 DECAPx2_ASAP7_75t_R FILLER_295_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_295_783 ();
 DECAPx1_ASAP7_75t_R FILLER_295_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_793 ();
 DECAPx4_ASAP7_75t_R FILLER_295_820 ();
 DECAPx2_ASAP7_75t_R FILLER_295_839 ();
 FILLER_ASAP7_75t_R FILLER_295_845 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_295_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_868 ();
 DECAPx4_ASAP7_75t_R FILLER_295_879 ();
 DECAPx6_ASAP7_75t_R FILLER_295_906 ();
 DECAPx1_ASAP7_75t_R FILLER_295_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_924 ();
 FILLERxp5_ASAP7_75t_R FILLER_295_933 ();
 DECAPx10_ASAP7_75t_R FILLER_296_2 ();
 DECAPx10_ASAP7_75t_R FILLER_296_24 ();
 DECAPx6_ASAP7_75t_R FILLER_296_46 ();
 DECAPx2_ASAP7_75t_R FILLER_296_60 ();
 DECAPx6_ASAP7_75t_R FILLER_296_92 ();
 DECAPx1_ASAP7_75t_R FILLER_296_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_110 ();
 FILLER_ASAP7_75t_R FILLER_296_123 ();
 DECAPx6_ASAP7_75t_R FILLER_296_131 ();
 DECAPx2_ASAP7_75t_R FILLER_296_145 ();
 DECAPx1_ASAP7_75t_R FILLER_296_183 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_187 ();
 FILLER_ASAP7_75t_R FILLER_296_213 ();
 DECAPx6_ASAP7_75t_R FILLER_296_221 ();
 FILLER_ASAP7_75t_R FILLER_296_235 ();
 DECAPx6_ASAP7_75t_R FILLER_296_271 ();
 DECAPx2_ASAP7_75t_R FILLER_296_285 ();
 DECAPx6_ASAP7_75t_R FILLER_296_297 ();
 DECAPx2_ASAP7_75t_R FILLER_296_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_317 ();
 DECAPx2_ASAP7_75t_R FILLER_296_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_330 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_296_339 ();
 DECAPx2_ASAP7_75t_R FILLER_296_353 ();
 DECAPx6_ASAP7_75t_R FILLER_296_365 ();
 DECAPx2_ASAP7_75t_R FILLER_296_379 ();
 DECAPx1_ASAP7_75t_R FILLER_296_391 ();
 DECAPx6_ASAP7_75t_R FILLER_296_398 ();
 DECAPx1_ASAP7_75t_R FILLER_296_412 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_416 ();
 DECAPx2_ASAP7_75t_R FILLER_296_423 ();
 FILLER_ASAP7_75t_R FILLER_296_429 ();
 DECAPx6_ASAP7_75t_R FILLER_296_443 ();
 DECAPx1_ASAP7_75t_R FILLER_296_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_461 ();
 DECAPx4_ASAP7_75t_R FILLER_296_464 ();
 FILLER_ASAP7_75t_R FILLER_296_474 ();
 DECAPx10_ASAP7_75t_R FILLER_296_479 ();
 DECAPx10_ASAP7_75t_R FILLER_296_501 ();
 DECAPx2_ASAP7_75t_R FILLER_296_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_529 ();
 DECAPx4_ASAP7_75t_R FILLER_296_539 ();
 FILLER_ASAP7_75t_R FILLER_296_549 ();
 DECAPx4_ASAP7_75t_R FILLER_296_554 ();
 DECAPx4_ASAP7_75t_R FILLER_296_567 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_577 ();
 FILLER_ASAP7_75t_R FILLER_296_590 ();
 DECAPx10_ASAP7_75t_R FILLER_296_606 ();
 DECAPx6_ASAP7_75t_R FILLER_296_628 ();
 DECAPx1_ASAP7_75t_R FILLER_296_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_672 ();
 DECAPx10_ASAP7_75t_R FILLER_296_685 ();
 DECAPx4_ASAP7_75t_R FILLER_296_707 ();
 FILLER_ASAP7_75t_R FILLER_296_717 ();
 DECAPx6_ASAP7_75t_R FILLER_296_727 ();
 FILLER_ASAP7_75t_R FILLER_296_741 ();
 DECAPx2_ASAP7_75t_R FILLER_296_753 ();
 DECAPx10_ASAP7_75t_R FILLER_296_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_807 ();
 DECAPx4_ASAP7_75t_R FILLER_296_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_821 ();
 DECAPx1_ASAP7_75t_R FILLER_296_854 ();
 FILLER_ASAP7_75t_R FILLER_296_884 ();
 DECAPx1_ASAP7_75t_R FILLER_296_912 ();
 FILLERxp5_ASAP7_75t_R FILLER_296_916 ();
 FILLER_ASAP7_75t_R FILLER_296_932 ();
 DECAPx10_ASAP7_75t_R FILLER_297_2 ();
 DECAPx10_ASAP7_75t_R FILLER_297_24 ();
 DECAPx10_ASAP7_75t_R FILLER_297_46 ();
 DECAPx4_ASAP7_75t_R FILLER_297_68 ();
 FILLER_ASAP7_75t_R FILLER_297_78 ();
 DECAPx4_ASAP7_75t_R FILLER_297_92 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_108 ();
 FILLER_ASAP7_75t_R FILLER_297_131 ();
 DECAPx1_ASAP7_75t_R FILLER_297_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_151 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_202 ();
 DECAPx2_ASAP7_75t_R FILLER_297_237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_243 ();
 DECAPx4_ASAP7_75t_R FILLER_297_261 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_271 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_282 ();
 DECAPx10_ASAP7_75t_R FILLER_297_291 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_313 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_329 ();
 DECAPx1_ASAP7_75t_R FILLER_297_338 ();
 DECAPx10_ASAP7_75t_R FILLER_297_377 ();
 DECAPx4_ASAP7_75t_R FILLER_297_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_409 ();
 DECAPx6_ASAP7_75t_R FILLER_297_424 ();
 FILLER_ASAP7_75t_R FILLER_297_438 ();
 DECAPx2_ASAP7_75t_R FILLER_297_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_456 ();
 DECAPx10_ASAP7_75t_R FILLER_297_460 ();
 DECAPx6_ASAP7_75t_R FILLER_297_482 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_496 ();
 DECAPx1_ASAP7_75t_R FILLER_297_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_529 ();
 DECAPx4_ASAP7_75t_R FILLER_297_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_554 ();
 DECAPx6_ASAP7_75t_R FILLER_297_558 ();
 FILLER_ASAP7_75t_R FILLER_297_572 ();
 DECAPx10_ASAP7_75t_R FILLER_297_588 ();
 DECAPx2_ASAP7_75t_R FILLER_297_610 ();
 DECAPx10_ASAP7_75t_R FILLER_297_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_644 ();
 DECAPx2_ASAP7_75t_R FILLER_297_648 ();
 FILLER_ASAP7_75t_R FILLER_297_654 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_659 ();
 DECAPx10_ASAP7_75t_R FILLER_297_693 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_715 ();
 DECAPx1_ASAP7_75t_R FILLER_297_726 ();
 DECAPx10_ASAP7_75t_R FILLER_297_778 ();
 DECAPx10_ASAP7_75t_R FILLER_297_800 ();
 DECAPx2_ASAP7_75t_R FILLER_297_822 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_828 ();
 DECAPx2_ASAP7_75t_R FILLER_297_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_297_840 ();
 DECAPx2_ASAP7_75t_R FILLER_297_846 ();
 FILLER_ASAP7_75t_R FILLER_297_852 ();
 DECAPx4_ASAP7_75t_R FILLER_297_872 ();
 FILLER_ASAP7_75t_R FILLER_297_882 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_890 ();
 DECAPx2_ASAP7_75t_R FILLER_297_894 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_900 ();
 FILLER_ASAP7_75t_R FILLER_297_904 ();
 DECAPx1_ASAP7_75t_R FILLER_297_921 ();
 FILLERxp5_ASAP7_75t_R FILLER_297_933 ();
 DECAPx10_ASAP7_75t_R FILLER_298_2 ();
 DECAPx10_ASAP7_75t_R FILLER_298_24 ();
 DECAPx10_ASAP7_75t_R FILLER_298_46 ();
 DECAPx10_ASAP7_75t_R FILLER_298_68 ();
 DECAPx1_ASAP7_75t_R FILLER_298_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_94 ();
 DECAPx2_ASAP7_75t_R FILLER_298_101 ();
 FILLER_ASAP7_75t_R FILLER_298_107 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_231 ();
 DECAPx6_ASAP7_75t_R FILLER_298_245 ();
 DECAPx2_ASAP7_75t_R FILLER_298_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_265 ();
 DECAPx2_ASAP7_75t_R FILLER_298_302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_298_308 ();
 DECAPx10_ASAP7_75t_R FILLER_298_331 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_298_360 ();
 DECAPx2_ASAP7_75t_R FILLER_298_366 ();
 DECAPx4_ASAP7_75t_R FILLER_298_394 ();
 FILLER_ASAP7_75t_R FILLER_298_404 ();
 DECAPx2_ASAP7_75t_R FILLER_298_432 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_298_438 ();
 DECAPx2_ASAP7_75t_R FILLER_298_464 ();
 DECAPx2_ASAP7_75t_R FILLER_298_479 ();
 DECAPx1_ASAP7_75t_R FILLER_298_488 ();
 FILLER_ASAP7_75t_R FILLER_298_521 ();
 FILLER_ASAP7_75t_R FILLER_298_526 ();
 DECAPx1_ASAP7_75t_R FILLER_298_542 ();
 DECAPx4_ASAP7_75t_R FILLER_298_555 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_565 ();
 DECAPx2_ASAP7_75t_R FILLER_298_583 ();
 FILLER_ASAP7_75t_R FILLER_298_589 ();
 DECAPx4_ASAP7_75t_R FILLER_298_601 ();
 FILLER_ASAP7_75t_R FILLER_298_611 ();
 DECAPx10_ASAP7_75t_R FILLER_298_630 ();
 DECAPx6_ASAP7_75t_R FILLER_298_652 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_666 ();
 FILLER_ASAP7_75t_R FILLER_298_676 ();
 DECAPx2_ASAP7_75t_R FILLER_298_681 ();
 DECAPx10_ASAP7_75t_R FILLER_298_690 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_298_712 ();
 DECAPx10_ASAP7_75t_R FILLER_298_761 ();
 DECAPx10_ASAP7_75t_R FILLER_298_783 ();
 DECAPx1_ASAP7_75t_R FILLER_298_805 ();
 FILLERxp5_ASAP7_75t_R FILLER_298_809 ();
 DECAPx10_ASAP7_75t_R FILLER_298_820 ();
 DECAPx10_ASAP7_75t_R FILLER_298_842 ();
 DECAPx4_ASAP7_75t_R FILLER_298_864 ();
 DECAPx10_ASAP7_75t_R FILLER_298_882 ();
 DECAPx1_ASAP7_75t_R FILLER_298_904 ();
 DECAPx10_ASAP7_75t_R FILLER_299_2 ();
 DECAPx10_ASAP7_75t_R FILLER_299_24 ();
 DECAPx10_ASAP7_75t_R FILLER_299_46 ();
 DECAPx2_ASAP7_75t_R FILLER_299_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_74 ();
 FILLER_ASAP7_75t_R FILLER_299_81 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_299_108 ();
 DECAPx2_ASAP7_75t_R FILLER_299_122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_299_128 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_149 ();
 DECAPx2_ASAP7_75t_R FILLER_299_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_299_162 ();
 DECAPx2_ASAP7_75t_R FILLER_299_171 ();
 FILLER_ASAP7_75t_R FILLER_299_177 ();
 DECAPx2_ASAP7_75t_R FILLER_299_254 ();
 FILLER_ASAP7_75t_R FILLER_299_260 ();
 FILLER_ASAP7_75t_R FILLER_299_268 ();
 DECAPx1_ASAP7_75t_R FILLER_299_276 ();
 DECAPx1_ASAP7_75t_R FILLER_299_286 ();
 DECAPx4_ASAP7_75t_R FILLER_299_293 ();
 DECAPx6_ASAP7_75t_R FILLER_299_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_299_329 ();
 FILLER_ASAP7_75t_R FILLER_299_338 ();
 DECAPx6_ASAP7_75t_R FILLER_299_343 ();
 DECAPx2_ASAP7_75t_R FILLER_299_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_363 ();
 FILLER_ASAP7_75t_R FILLER_299_376 ();
 DECAPx6_ASAP7_75t_R FILLER_299_407 ();
 DECAPx2_ASAP7_75t_R FILLER_299_424 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_430 ();
 DECAPx2_ASAP7_75t_R FILLER_299_437 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_299_443 ();
 FILLER_ASAP7_75t_R FILLER_299_458 ();
 FILLER_ASAP7_75t_R FILLER_299_494 ();
 DECAPx6_ASAP7_75t_R FILLER_299_516 ();
 DECAPx2_ASAP7_75t_R FILLER_299_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_536 ();
 DECAPx2_ASAP7_75t_R FILLER_299_543 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_577 ();
 DECAPx2_ASAP7_75t_R FILLER_299_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_629 ();
 DECAPx2_ASAP7_75t_R FILLER_299_650 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_656 ();
 DECAPx10_ASAP7_75t_R FILLER_299_671 ();
 DECAPx10_ASAP7_75t_R FILLER_299_693 ();
 DECAPx6_ASAP7_75t_R FILLER_299_715 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_729 ();
 DECAPx4_ASAP7_75t_R FILLER_299_733 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_743 ();
 FILLER_ASAP7_75t_R FILLER_299_747 ();
 DECAPx10_ASAP7_75t_R FILLER_299_752 ();
 DECAPx2_ASAP7_75t_R FILLER_299_774 ();
 FILLER_ASAP7_75t_R FILLER_299_796 ();
 DECAPx4_ASAP7_75t_R FILLER_299_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_834 ();
 DECAPx6_ASAP7_75t_R FILLER_299_841 ();
 DECAPx2_ASAP7_75t_R FILLER_299_855 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_861 ();
 FILLER_ASAP7_75t_R FILLER_299_865 ();
 DECAPx1_ASAP7_75t_R FILLER_299_870 ();
 DECAPx10_ASAP7_75t_R FILLER_299_884 ();
 DECAPx6_ASAP7_75t_R FILLER_299_906 ();
 DECAPx1_ASAP7_75t_R FILLER_299_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_299_924 ();
 DECAPx1_ASAP7_75t_R FILLER_299_930 ();
 DECAPx10_ASAP7_75t_R FILLER_300_2 ();
 DECAPx10_ASAP7_75t_R FILLER_300_24 ();
 DECAPx10_ASAP7_75t_R FILLER_300_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_68 ();
 DECAPx10_ASAP7_75t_R FILLER_300_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_139 ();
 DECAPx10_ASAP7_75t_R FILLER_300_143 ();
 DECAPx10_ASAP7_75t_R FILLER_300_165 ();
 DECAPx1_ASAP7_75t_R FILLER_300_187 ();
 DECAPx2_ASAP7_75t_R FILLER_300_194 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_233 ();
 DECAPx1_ASAP7_75t_R FILLER_300_246 ();
 DECAPx6_ASAP7_75t_R FILLER_300_281 ();
 DECAPx1_ASAP7_75t_R FILLER_300_295 ();
 DECAPx2_ASAP7_75t_R FILLER_300_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_357 ();
 DECAPx10_ASAP7_75t_R FILLER_300_364 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_386 ();
 DECAPx2_ASAP7_75t_R FILLER_300_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_402 ();
 DECAPx1_ASAP7_75t_R FILLER_300_409 ();
 DECAPx2_ASAP7_75t_R FILLER_300_422 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_300_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_300_438 ();
 DECAPx1_ASAP7_75t_R FILLER_300_448 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_461 ();
 DECAPx1_ASAP7_75t_R FILLER_300_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_468 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_300_475 ();
 DECAPx1_ASAP7_75t_R FILLER_300_499 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_503 ();
 DECAPx6_ASAP7_75t_R FILLER_300_509 ();
 FILLER_ASAP7_75t_R FILLER_300_523 ();
 DECAPx1_ASAP7_75t_R FILLER_300_528 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_532 ();
 DECAPx1_ASAP7_75t_R FILLER_300_547 ();
 DECAPx2_ASAP7_75t_R FILLER_300_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_563 ();
 DECAPx10_ASAP7_75t_R FILLER_300_570 ();
 FILLER_ASAP7_75t_R FILLER_300_592 ();
 DECAPx10_ASAP7_75t_R FILLER_300_674 ();
 DECAPx6_ASAP7_75t_R FILLER_300_696 ();
 DECAPx1_ASAP7_75t_R FILLER_300_710 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_714 ();
 DECAPx10_ASAP7_75t_R FILLER_300_718 ();
 DECAPx10_ASAP7_75t_R FILLER_300_740 ();
 DECAPx2_ASAP7_75t_R FILLER_300_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_774 ();
 FILLER_ASAP7_75t_R FILLER_300_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_868 ();
 DECAPx2_ASAP7_75t_R FILLER_300_902 ();
 DECAPx6_ASAP7_75t_R FILLER_300_915 ();
 DECAPx1_ASAP7_75t_R FILLER_300_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_300_933 ();
 DECAPx10_ASAP7_75t_R FILLER_301_2 ();
 DECAPx10_ASAP7_75t_R FILLER_301_24 ();
 DECAPx10_ASAP7_75t_R FILLER_301_46 ();
 DECAPx2_ASAP7_75t_R FILLER_301_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_74 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_86 ();
 DECAPx10_ASAP7_75t_R FILLER_301_114 ();
 DECAPx10_ASAP7_75t_R FILLER_301_136 ();
 DECAPx10_ASAP7_75t_R FILLER_301_158 ();
 DECAPx10_ASAP7_75t_R FILLER_301_180 ();
 DECAPx4_ASAP7_75t_R FILLER_301_202 ();
 DECAPx10_ASAP7_75t_R FILLER_301_221 ();
 DECAPx4_ASAP7_75t_R FILLER_301_243 ();
 DECAPx1_ASAP7_75t_R FILLER_301_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_263 ();
 DECAPx6_ASAP7_75t_R FILLER_301_267 ();
 DECAPx1_ASAP7_75t_R FILLER_301_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_285 ();
 FILLER_ASAP7_75t_R FILLER_301_312 ();
 DECAPx4_ASAP7_75t_R FILLER_301_317 ();
 DECAPx6_ASAP7_75t_R FILLER_301_333 ();
 FILLER_ASAP7_75t_R FILLER_301_347 ();
 DECAPx10_ASAP7_75t_R FILLER_301_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_423 ();
 DECAPx6_ASAP7_75t_R FILLER_301_462 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_476 ();
 FILLER_ASAP7_75t_R FILLER_301_489 ();
 DECAPx10_ASAP7_75t_R FILLER_301_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_518 ();
 DECAPx4_ASAP7_75t_R FILLER_301_522 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_532 ();
 DECAPx10_ASAP7_75t_R FILLER_301_547 ();
 DECAPx4_ASAP7_75t_R FILLER_301_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_579 ();
 DECAPx6_ASAP7_75t_R FILLER_301_591 ();
 DECAPx6_ASAP7_75t_R FILLER_301_612 ();
 DECAPx1_ASAP7_75t_R FILLER_301_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_630 ();
 DECAPx2_ASAP7_75t_R FILLER_301_646 ();
 DECAPx10_ASAP7_75t_R FILLER_301_675 ();
 DECAPx4_ASAP7_75t_R FILLER_301_697 ();
 FILLER_ASAP7_75t_R FILLER_301_707 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_721 ();
 DECAPx10_ASAP7_75t_R FILLER_301_736 ();
 DECAPx2_ASAP7_75t_R FILLER_301_758 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_793 ();
 FILLER_ASAP7_75t_R FILLER_301_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_301_807 ();
 DECAPx4_ASAP7_75t_R FILLER_301_813 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_823 ();
 DECAPx1_ASAP7_75t_R FILLER_301_830 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_881 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_895 ();
 FILLERxp5_ASAP7_75t_R FILLER_301_914 ();
 DECAPx1_ASAP7_75t_R FILLER_301_930 ();
 DECAPx10_ASAP7_75t_R FILLER_302_2 ();
 DECAPx10_ASAP7_75t_R FILLER_302_24 ();
 DECAPx10_ASAP7_75t_R FILLER_302_46 ();
 DECAPx6_ASAP7_75t_R FILLER_302_68 ();
 DECAPx2_ASAP7_75t_R FILLER_302_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_112 ();
 DECAPx2_ASAP7_75t_R FILLER_302_121 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_127 ();
 DECAPx6_ASAP7_75t_R FILLER_302_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_150 ();
 DECAPx1_ASAP7_75t_R FILLER_302_177 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_181 ();
 FILLER_ASAP7_75t_R FILLER_302_196 ();
 DECAPx10_ASAP7_75t_R FILLER_302_204 ();
 DECAPx6_ASAP7_75t_R FILLER_302_226 ();
 FILLER_ASAP7_75t_R FILLER_302_240 ();
 DECAPx10_ASAP7_75t_R FILLER_302_254 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_276 ();
 DECAPx1_ASAP7_75t_R FILLER_302_285 ();
 DECAPx10_ASAP7_75t_R FILLER_302_295 ();
 DECAPx10_ASAP7_75t_R FILLER_302_317 ();
 DECAPx1_ASAP7_75t_R FILLER_302_349 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_353 ();
 DECAPx1_ASAP7_75t_R FILLER_302_360 ();
 DECAPx10_ASAP7_75t_R FILLER_302_367 ();
 DECAPx1_ASAP7_75t_R FILLER_302_389 ();
 DECAPx4_ASAP7_75t_R FILLER_302_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_409 ();
 DECAPx4_ASAP7_75t_R FILLER_302_415 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_425 ();
 DECAPx2_ASAP7_75t_R FILLER_302_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_441 ();
 DECAPx6_ASAP7_75t_R FILLER_302_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_461 ();
 DECAPx10_ASAP7_75t_R FILLER_302_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_496 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_508 ();
 DECAPx10_ASAP7_75t_R FILLER_302_531 ();
 DECAPx4_ASAP7_75t_R FILLER_302_553 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_563 ();
 DECAPx10_ASAP7_75t_R FILLER_302_593 ();
 DECAPx10_ASAP7_75t_R FILLER_302_615 ();
 DECAPx4_ASAP7_75t_R FILLER_302_637 ();
 FILLER_ASAP7_75t_R FILLER_302_647 ();
 DECAPx10_ASAP7_75t_R FILLER_302_652 ();
 DECAPx1_ASAP7_75t_R FILLER_302_674 ();
 DECAPx6_ASAP7_75t_R FILLER_302_695 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_732 ();
 FILLER_ASAP7_75t_R FILLER_302_759 ();
 DECAPx2_ASAP7_75t_R FILLER_302_793 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_302_799 ();
 DECAPx10_ASAP7_75t_R FILLER_302_817 ();
 DECAPx1_ASAP7_75t_R FILLER_302_839 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_843 ();
 DECAPx1_ASAP7_75t_R FILLER_302_851 ();
 FILLERxp5_ASAP7_75t_R FILLER_302_855 ();
 DECAPx10_ASAP7_75t_R FILLER_302_868 ();
 FILLER_ASAP7_75t_R FILLER_302_890 ();
 DECAPx4_ASAP7_75t_R FILLER_302_898 ();
 DECAPx10_ASAP7_75t_R FILLER_303_2 ();
 DECAPx10_ASAP7_75t_R FILLER_303_24 ();
 DECAPx10_ASAP7_75t_R FILLER_303_46 ();
 DECAPx6_ASAP7_75t_R FILLER_303_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_82 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_111 ();
 DECAPx1_ASAP7_75t_R FILLER_303_132 ();
 DECAPx1_ASAP7_75t_R FILLER_303_209 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_219 ();
 DECAPx6_ASAP7_75t_R FILLER_303_223 ();
 FILLER_ASAP7_75t_R FILLER_303_237 ();
 DECAPx2_ASAP7_75t_R FILLER_303_265 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_271 ();
 DECAPx4_ASAP7_75t_R FILLER_303_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_316 ();
 DECAPx1_ASAP7_75t_R FILLER_303_320 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_324 ();
 DECAPx10_ASAP7_75t_R FILLER_303_409 ();
 DECAPx2_ASAP7_75t_R FILLER_303_431 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_437 ();
 DECAPx6_ASAP7_75t_R FILLER_303_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_457 ();
 DECAPx2_ASAP7_75t_R FILLER_303_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_470 ();
 DECAPx2_ASAP7_75t_R FILLER_303_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_489 ();
 DECAPx1_ASAP7_75t_R FILLER_303_513 ();
 DECAPx2_ASAP7_75t_R FILLER_303_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_543 ();
 DECAPx4_ASAP7_75t_R FILLER_303_560 ();
 FILLER_ASAP7_75t_R FILLER_303_570 ();
 DECAPx10_ASAP7_75t_R FILLER_303_578 ();
 DECAPx4_ASAP7_75t_R FILLER_303_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_610 ();
 DECAPx10_ASAP7_75t_R FILLER_303_625 ();
 DECAPx10_ASAP7_75t_R FILLER_303_647 ();
 DECAPx2_ASAP7_75t_R FILLER_303_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_675 ();
 DECAPx6_ASAP7_75t_R FILLER_303_699 ();
 DECAPx1_ASAP7_75t_R FILLER_303_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_717 ();
 DECAPx10_ASAP7_75t_R FILLER_303_785 ();
 DECAPx2_ASAP7_75t_R FILLER_303_807 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_303_813 ();
 DECAPx10_ASAP7_75t_R FILLER_303_826 ();
 DECAPx6_ASAP7_75t_R FILLER_303_848 ();
 DECAPx2_ASAP7_75t_R FILLER_303_862 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_868 ();
 DECAPx10_ASAP7_75t_R FILLER_303_889 ();
 DECAPx2_ASAP7_75t_R FILLER_303_917 ();
 FILLER_ASAP7_75t_R FILLER_303_923 ();
 DECAPx2_ASAP7_75t_R FILLER_303_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_303_933 ();
 DECAPx10_ASAP7_75t_R FILLER_304_2 ();
 DECAPx10_ASAP7_75t_R FILLER_304_24 ();
 DECAPx10_ASAP7_75t_R FILLER_304_46 ();
 DECAPx4_ASAP7_75t_R FILLER_304_68 ();
 FILLER_ASAP7_75t_R FILLER_304_78 ();
 DECAPx6_ASAP7_75t_R FILLER_304_86 ();
 DECAPx4_ASAP7_75t_R FILLER_304_103 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_119 ();
 DECAPx4_ASAP7_75t_R FILLER_304_126 ();
 FILLER_ASAP7_75t_R FILLER_304_136 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_176 ();
 FILLER_ASAP7_75t_R FILLER_304_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_196 ();
 DECAPx1_ASAP7_75t_R FILLER_304_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_204 ();
 DECAPx10_ASAP7_75t_R FILLER_304_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_253 ();
 DECAPx2_ASAP7_75t_R FILLER_304_257 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_274 ();
 DECAPx1_ASAP7_75t_R FILLER_304_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_287 ();
 DECAPx10_ASAP7_75t_R FILLER_304_317 ();
 DECAPx1_ASAP7_75t_R FILLER_304_348 ();
 DECAPx2_ASAP7_75t_R FILLER_304_355 ();
 FILLER_ASAP7_75t_R FILLER_304_361 ();
 DECAPx4_ASAP7_75t_R FILLER_304_378 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_394 ();
 DECAPx2_ASAP7_75t_R FILLER_304_400 ();
 DECAPx6_ASAP7_75t_R FILLER_304_409 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_423 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_461 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_474 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_487 ();
 DECAPx6_ASAP7_75t_R FILLER_304_504 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_518 ();
 DECAPx10_ASAP7_75t_R FILLER_304_525 ();
 DECAPx1_ASAP7_75t_R FILLER_304_547 ();
 DECAPx1_ASAP7_75t_R FILLER_304_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_558 ();
 DECAPx2_ASAP7_75t_R FILLER_304_562 ();
 DECAPx2_ASAP7_75t_R FILLER_304_571 ();
 FILLER_ASAP7_75t_R FILLER_304_577 ();
 DECAPx1_ASAP7_75t_R FILLER_304_582 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_586 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_593 ();
 DECAPx1_ASAP7_75t_R FILLER_304_611 ();
 DECAPx1_ASAP7_75t_R FILLER_304_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_626 ();
 DECAPx2_ASAP7_75t_R FILLER_304_630 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_636 ();
 DECAPx6_ASAP7_75t_R FILLER_304_642 ();
 DECAPx1_ASAP7_75t_R FILLER_304_656 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_660 ();
 DECAPx4_ASAP7_75t_R FILLER_304_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_674 ();
 DECAPx10_ASAP7_75t_R FILLER_304_690 ();
 DECAPx6_ASAP7_75t_R FILLER_304_712 ();
 DECAPx2_ASAP7_75t_R FILLER_304_726 ();
 DECAPx4_ASAP7_75t_R FILLER_304_735 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_745 ();
 DECAPx10_ASAP7_75t_R FILLER_304_763 ();
 DECAPx10_ASAP7_75t_R FILLER_304_785 ();
 DECAPx2_ASAP7_75t_R FILLER_304_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_813 ();
 DECAPx2_ASAP7_75t_R FILLER_304_840 ();
 FILLERxp5_ASAP7_75t_R FILLER_304_846 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_850 ();
 DECAPx10_ASAP7_75t_R FILLER_304_859 ();
 DECAPx2_ASAP7_75t_R FILLER_304_881 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_887 ();
 DECAPx6_ASAP7_75t_R FILLER_304_893 ();
 DECAPx1_ASAP7_75t_R FILLER_304_907 ();
 DECAPx6_ASAP7_75t_R FILLER_304_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_304_931 ();
 DECAPx10_ASAP7_75t_R FILLER_305_2 ();
 DECAPx10_ASAP7_75t_R FILLER_305_24 ();
 DECAPx10_ASAP7_75t_R FILLER_305_46 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_68 ();
 DECAPx6_ASAP7_75t_R FILLER_305_97 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_111 ();
 DECAPx1_ASAP7_75t_R FILLER_305_123 ();
 FILLER_ASAP7_75t_R FILLER_305_144 ();
 DECAPx1_ASAP7_75t_R FILLER_305_152 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_162 ();
 DECAPx10_ASAP7_75t_R FILLER_305_168 ();
 DECAPx6_ASAP7_75t_R FILLER_305_190 ();
 DECAPx1_ASAP7_75t_R FILLER_305_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_208 ();
 DECAPx1_ASAP7_75t_R FILLER_305_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_234 ();
 DECAPx2_ASAP7_75t_R FILLER_305_242 ();
 FILLER_ASAP7_75t_R FILLER_305_254 ();
 DECAPx1_ASAP7_75t_R FILLER_305_259 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_263 ();
 DECAPx6_ASAP7_75t_R FILLER_305_270 ();
 DECAPx2_ASAP7_75t_R FILLER_305_284 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_323 ();
 DECAPx6_ASAP7_75t_R FILLER_305_330 ();
 DECAPx1_ASAP7_75t_R FILLER_305_344 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_348 ();
 DECAPx10_ASAP7_75t_R FILLER_305_355 ();
 DECAPx10_ASAP7_75t_R FILLER_305_377 ();
 DECAPx2_ASAP7_75t_R FILLER_305_399 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_405 ();
 FILLER_ASAP7_75t_R FILLER_305_414 ();
 FILLER_ASAP7_75t_R FILLER_305_428 ();
 DECAPx1_ASAP7_75t_R FILLER_305_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_440 ();
 DECAPx10_ASAP7_75t_R FILLER_305_493 ();
 DECAPx10_ASAP7_75t_R FILLER_305_515 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_579 ();
 DECAPx1_ASAP7_75t_R FILLER_305_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_628 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_643 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_648 ();
 DECAPx10_ASAP7_75t_R FILLER_305_668 ();
 DECAPx10_ASAP7_75t_R FILLER_305_690 ();
 DECAPx10_ASAP7_75t_R FILLER_305_712 ();
 DECAPx10_ASAP7_75t_R FILLER_305_734 ();
 DECAPx10_ASAP7_75t_R FILLER_305_756 ();
 DECAPx2_ASAP7_75t_R FILLER_305_778 ();
 FILLER_ASAP7_75t_R FILLER_305_784 ();
 FILLER_ASAP7_75t_R FILLER_305_792 ();
 DECAPx2_ASAP7_75t_R FILLER_305_800 ();
 FILLER_ASAP7_75t_R FILLER_305_806 ();
 DECAPx1_ASAP7_75t_R FILLER_305_842 ();
 FILLER_ASAP7_75t_R FILLER_305_861 ();
 DECAPx6_ASAP7_75t_R FILLER_305_871 ();
 DECAPx2_ASAP7_75t_R FILLER_305_885 ();
 DECAPx1_ASAP7_75t_R FILLER_305_897 ();
 FILLER_ASAP7_75t_R FILLER_305_904 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_305_922 ();
 DECAPx2_ASAP7_75t_R FILLER_305_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_305_933 ();
 DECAPx10_ASAP7_75t_R FILLER_306_2 ();
 DECAPx10_ASAP7_75t_R FILLER_306_24 ();
 DECAPx10_ASAP7_75t_R FILLER_306_46 ();
 DECAPx6_ASAP7_75t_R FILLER_306_68 ();
 FILLER_ASAP7_75t_R FILLER_306_91 ();
 DECAPx2_ASAP7_75t_R FILLER_306_96 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_102 ();
 DECAPx1_ASAP7_75t_R FILLER_306_139 ();
 DECAPx10_ASAP7_75t_R FILLER_306_149 ();
 DECAPx6_ASAP7_75t_R FILLER_306_171 ();
 FILLER_ASAP7_75t_R FILLER_306_185 ();
 DECAPx10_ASAP7_75t_R FILLER_306_196 ();
 DECAPx1_ASAP7_75t_R FILLER_306_218 ();
 FILLER_ASAP7_75t_R FILLER_306_228 ();
 DECAPx1_ASAP7_75t_R FILLER_306_236 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_240 ();
 DECAPx1_ASAP7_75t_R FILLER_306_267 ();
 DECAPx10_ASAP7_75t_R FILLER_306_277 ();
 FILLER_ASAP7_75t_R FILLER_306_299 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_310 ();
 DECAPx10_ASAP7_75t_R FILLER_306_337 ();
 DECAPx4_ASAP7_75t_R FILLER_306_365 ();
 FILLER_ASAP7_75t_R FILLER_306_375 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_393 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_402 ();
 DECAPx1_ASAP7_75t_R FILLER_306_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_425 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_461 ();
 DECAPx1_ASAP7_75t_R FILLER_306_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_468 ();
 DECAPx4_ASAP7_75t_R FILLER_306_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_485 ();
 DECAPx10_ASAP7_75t_R FILLER_306_496 ();
 DECAPx6_ASAP7_75t_R FILLER_306_518 ();
 DECAPx2_ASAP7_75t_R FILLER_306_532 ();
 DECAPx2_ASAP7_75t_R FILLER_306_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_558 ();
 DECAPx4_ASAP7_75t_R FILLER_306_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_580 ();
 DECAPx1_ASAP7_75t_R FILLER_306_600 ();
 DECAPx4_ASAP7_75t_R FILLER_306_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_617 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_621 ();
 DECAPx10_ASAP7_75t_R FILLER_306_681 ();
 DECAPx10_ASAP7_75t_R FILLER_306_703 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_725 ();
 DECAPx10_ASAP7_75t_R FILLER_306_734 ();
 DECAPx10_ASAP7_75t_R FILLER_306_756 ();
 DECAPx1_ASAP7_75t_R FILLER_306_778 ();
 FILLER_ASAP7_75t_R FILLER_306_791 ();
 DECAPx2_ASAP7_75t_R FILLER_306_808 ();
 FILLER_ASAP7_75t_R FILLER_306_814 ();
 FILLER_ASAP7_75t_R FILLER_306_824 ();
 DECAPx2_ASAP7_75t_R FILLER_306_852 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_858 ();
 DECAPx2_ASAP7_75t_R FILLER_306_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_306_920 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_306_931 ();
 DECAPx10_ASAP7_75t_R FILLER_307_2 ();
 DECAPx10_ASAP7_75t_R FILLER_307_24 ();
 DECAPx10_ASAP7_75t_R FILLER_307_46 ();
 DECAPx6_ASAP7_75t_R FILLER_307_68 ();
 DECAPx2_ASAP7_75t_R FILLER_307_88 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_94 ();
 DECAPx1_ASAP7_75t_R FILLER_307_105 ();
 DECAPx10_ASAP7_75t_R FILLER_307_115 ();
 DECAPx10_ASAP7_75t_R FILLER_307_137 ();
 DECAPx4_ASAP7_75t_R FILLER_307_159 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_169 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_178 ();
 DECAPx10_ASAP7_75t_R FILLER_307_214 ();
 DECAPx2_ASAP7_75t_R FILLER_307_236 ();
 FILLER_ASAP7_75t_R FILLER_307_242 ();
 DECAPx1_ASAP7_75t_R FILLER_307_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_278 ();
 DECAPx6_ASAP7_75t_R FILLER_307_292 ();
 DECAPx1_ASAP7_75t_R FILLER_307_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_325 ();
 DECAPx2_ASAP7_75t_R FILLER_307_329 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_335 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_361 ();
 DECAPx1_ASAP7_75t_R FILLER_307_370 ();
 DECAPx1_ASAP7_75t_R FILLER_307_380 ();
 DECAPx2_ASAP7_75t_R FILLER_307_422 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_428 ();
 DECAPx10_ASAP7_75t_R FILLER_307_463 ();
 DECAPx4_ASAP7_75t_R FILLER_307_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_495 ();
 DECAPx2_ASAP7_75t_R FILLER_307_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_507 ();
 DECAPx1_ASAP7_75t_R FILLER_307_516 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_520 ();
 DECAPx6_ASAP7_75t_R FILLER_307_545 ();
 DECAPx1_ASAP7_75t_R FILLER_307_559 ();
 DECAPx1_ASAP7_75t_R FILLER_307_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_587 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_611 ();
 DECAPx10_ASAP7_75t_R FILLER_307_615 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_637 ();
 DECAPx1_ASAP7_75t_R FILLER_307_647 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_654 ();
 DECAPx10_ASAP7_75t_R FILLER_307_687 ();
 DECAPx2_ASAP7_75t_R FILLER_307_709 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_715 ();
 DECAPx1_ASAP7_75t_R FILLER_307_722 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_726 ();
 DECAPx1_ASAP7_75t_R FILLER_307_737 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_741 ();
 DECAPx10_ASAP7_75t_R FILLER_307_758 ();
 FILLER_ASAP7_75t_R FILLER_307_780 ();
 DECAPx2_ASAP7_75t_R FILLER_307_785 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_791 ();
 DECAPx6_ASAP7_75t_R FILLER_307_802 ();
 DECAPx2_ASAP7_75t_R FILLER_307_816 ();
 DECAPx1_ASAP7_75t_R FILLER_307_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_829 ();
 FILLER_ASAP7_75t_R FILLER_307_838 ();
 DECAPx6_ASAP7_75t_R FILLER_307_843 ();
 DECAPx2_ASAP7_75t_R FILLER_307_857 ();
 DECAPx1_ASAP7_75t_R FILLER_307_869 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_873 ();
 DECAPx2_ASAP7_75t_R FILLER_307_892 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_898 ();
 DECAPx6_ASAP7_75t_R FILLER_307_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_307_922 ();
 FILLERxp5_ASAP7_75t_R FILLER_307_933 ();
 DECAPx10_ASAP7_75t_R FILLER_308_2 ();
 DECAPx10_ASAP7_75t_R FILLER_308_24 ();
 DECAPx10_ASAP7_75t_R FILLER_308_46 ();
 FILLER_ASAP7_75t_R FILLER_308_68 ();
 DECAPx6_ASAP7_75t_R FILLER_308_110 ();
 DECAPx2_ASAP7_75t_R FILLER_308_124 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_130 ();
 DECAPx10_ASAP7_75t_R FILLER_308_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_308_156 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_188 ();
 DECAPx10_ASAP7_75t_R FILLER_308_226 ();
 DECAPx2_ASAP7_75t_R FILLER_308_248 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_254 ();
 FILLER_ASAP7_75t_R FILLER_308_261 ();
 DECAPx1_ASAP7_75t_R FILLER_308_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_274 ();
 DECAPx4_ASAP7_75t_R FILLER_308_301 ();
 DECAPx6_ASAP7_75t_R FILLER_308_318 ();
 DECAPx1_ASAP7_75t_R FILLER_308_332 ();
 FILLER_ASAP7_75t_R FILLER_308_350 ();
 DECAPx6_ASAP7_75t_R FILLER_308_387 ();
 DECAPx1_ASAP7_75t_R FILLER_308_407 ();
 DECAPx6_ASAP7_75t_R FILLER_308_414 ();
 DECAPx1_ASAP7_75t_R FILLER_308_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_432 ();
 DECAPx2_ASAP7_75t_R FILLER_308_464 ();
 DECAPx1_ASAP7_75t_R FILLER_308_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_480 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_499 ();
 FILLER_ASAP7_75t_R FILLER_308_523 ();
 DECAPx10_ASAP7_75t_R FILLER_308_539 ();
 DECAPx6_ASAP7_75t_R FILLER_308_561 ();
 DECAPx2_ASAP7_75t_R FILLER_308_589 ();
 DECAPx4_ASAP7_75t_R FILLER_308_612 ();
 FILLER_ASAP7_75t_R FILLER_308_622 ();
 DECAPx10_ASAP7_75t_R FILLER_308_627 ();
 FILLER_ASAP7_75t_R FILLER_308_649 ();
 DECAPx2_ASAP7_75t_R FILLER_308_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_660 ();
 DECAPx1_ASAP7_75t_R FILLER_308_664 ();
 DECAPx4_ASAP7_75t_R FILLER_308_671 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_681 ();
 DECAPx6_ASAP7_75t_R FILLER_308_694 ();
 DECAPx1_ASAP7_75t_R FILLER_308_708 ();
 FILLERxp5_ASAP7_75t_R FILLER_308_712 ();
 DECAPx1_ASAP7_75t_R FILLER_308_785 ();
 DECAPx10_ASAP7_75t_R FILLER_308_821 ();
 DECAPx10_ASAP7_75t_R FILLER_308_843 ();
 DECAPx10_ASAP7_75t_R FILLER_308_865 ();
 DECAPx4_ASAP7_75t_R FILLER_308_887 ();
 FILLER_ASAP7_75t_R FILLER_308_897 ();
 DECAPx10_ASAP7_75t_R FILLER_309_2 ();
 DECAPx10_ASAP7_75t_R FILLER_309_24 ();
 DECAPx10_ASAP7_75t_R FILLER_309_46 ();
 DECAPx2_ASAP7_75t_R FILLER_309_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_74 ();
 FILLER_ASAP7_75t_R FILLER_309_83 ();
 DECAPx2_ASAP7_75t_R FILLER_309_88 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_106 ();
 DECAPx6_ASAP7_75t_R FILLER_309_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_181 ();
 DECAPx1_ASAP7_75t_R FILLER_309_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_247 ();
 DECAPx10_ASAP7_75t_R FILLER_309_254 ();
 DECAPx2_ASAP7_75t_R FILLER_309_276 ();
 FILLER_ASAP7_75t_R FILLER_309_288 ();
 DECAPx4_ASAP7_75t_R FILLER_309_293 ();
 FILLER_ASAP7_75t_R FILLER_309_303 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_325 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_343 ();
 DECAPx4_ASAP7_75t_R FILLER_309_350 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_360 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_372 ();
 DECAPx10_ASAP7_75t_R FILLER_309_396 ();
 DECAPx4_ASAP7_75t_R FILLER_309_418 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_436 ();
 FILLER_ASAP7_75t_R FILLER_309_471 ();
 DECAPx1_ASAP7_75t_R FILLER_309_481 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_485 ();
 DECAPx2_ASAP7_75t_R FILLER_309_526 ();
 DECAPx4_ASAP7_75t_R FILLER_309_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_545 ();
 DECAPx4_ASAP7_75t_R FILLER_309_563 ();
 FILLER_ASAP7_75t_R FILLER_309_573 ();
 DECAPx2_ASAP7_75t_R FILLER_309_578 ();
 FILLER_ASAP7_75t_R FILLER_309_584 ();
 DECAPx2_ASAP7_75t_R FILLER_309_589 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_595 ();
 DECAPx10_ASAP7_75t_R FILLER_309_610 ();
 DECAPx10_ASAP7_75t_R FILLER_309_632 ();
 DECAPx10_ASAP7_75t_R FILLER_309_654 ();
 DECAPx2_ASAP7_75t_R FILLER_309_676 ();
 DECAPx6_ASAP7_75t_R FILLER_309_696 ();
 DECAPx2_ASAP7_75t_R FILLER_309_710 ();
 FILLER_ASAP7_75t_R FILLER_309_728 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_746 ();
 FILLERxp5_ASAP7_75t_R FILLER_309_756 ();
 DECAPx2_ASAP7_75t_R FILLER_309_790 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_309_796 ();
 FILLER_ASAP7_75t_R FILLER_309_809 ();
 DECAPx2_ASAP7_75t_R FILLER_309_820 ();
 FILLER_ASAP7_75t_R FILLER_309_826 ();
 DECAPx10_ASAP7_75t_R FILLER_309_843 ();
 DECAPx10_ASAP7_75t_R FILLER_309_865 ();
 DECAPx10_ASAP7_75t_R FILLER_309_887 ();
 DECAPx6_ASAP7_75t_R FILLER_309_909 ();
 FILLER_ASAP7_75t_R FILLER_309_923 ();
 DECAPx1_ASAP7_75t_R FILLER_309_930 ();
 DECAPx10_ASAP7_75t_R FILLER_310_2 ();
 DECAPx10_ASAP7_75t_R FILLER_310_24 ();
 DECAPx10_ASAP7_75t_R FILLER_310_46 ();
 DECAPx10_ASAP7_75t_R FILLER_310_68 ();
 DECAPx10_ASAP7_75t_R FILLER_310_90 ();
 FILLER_ASAP7_75t_R FILLER_310_112 ();
 DECAPx2_ASAP7_75t_R FILLER_310_129 ();
 DECAPx4_ASAP7_75t_R FILLER_310_173 ();
 FILLER_ASAP7_75t_R FILLER_310_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_228 ();
 DECAPx10_ASAP7_75t_R FILLER_310_257 ();
 DECAPx6_ASAP7_75t_R FILLER_310_279 ();
 DECAPx2_ASAP7_75t_R FILLER_310_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_299 ();
 DECAPx4_ASAP7_75t_R FILLER_310_380 ();
 DECAPx2_ASAP7_75t_R FILLER_310_402 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_414 ();
 DECAPx1_ASAP7_75t_R FILLER_310_421 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_425 ();
 FILLER_ASAP7_75t_R FILLER_310_460 ();
 DECAPx1_ASAP7_75t_R FILLER_310_485 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_498 ();
 DECAPx10_ASAP7_75t_R FILLER_310_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_536 ();
 DECAPx4_ASAP7_75t_R FILLER_310_540 ();
 FILLER_ASAP7_75t_R FILLER_310_556 ();
 DECAPx10_ASAP7_75t_R FILLER_310_563 ();
 DECAPx2_ASAP7_75t_R FILLER_310_585 ();
 FILLER_ASAP7_75t_R FILLER_310_591 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_639 ();
 DECAPx4_ASAP7_75t_R FILLER_310_656 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_666 ();
 DECAPx4_ASAP7_75t_R FILLER_310_672 ();
 FILLER_ASAP7_75t_R FILLER_310_682 ();
 DECAPx10_ASAP7_75t_R FILLER_310_696 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_718 ();
 DECAPx4_ASAP7_75t_R FILLER_310_724 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_734 ();
 DECAPx6_ASAP7_75t_R FILLER_310_740 ();
 FILLER_ASAP7_75t_R FILLER_310_754 ();
 FILLER_ASAP7_75t_R FILLER_310_779 ();
 DECAPx4_ASAP7_75t_R FILLER_310_791 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_801 ();
 DECAPx10_ASAP7_75t_R FILLER_310_807 ();
 FILLER_ASAP7_75t_R FILLER_310_829 ();
 DECAPx1_ASAP7_75t_R FILLER_310_834 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_310_844 ();
 DECAPx6_ASAP7_75t_R FILLER_310_875 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_889 ();
 DECAPx2_ASAP7_75t_R FILLER_310_901 ();
 FILLERxp5_ASAP7_75t_R FILLER_310_907 ();
 DECAPx10_ASAP7_75t_R FILLER_311_2 ();
 DECAPx10_ASAP7_75t_R FILLER_311_24 ();
 DECAPx10_ASAP7_75t_R FILLER_311_46 ();
 DECAPx4_ASAP7_75t_R FILLER_311_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_78 ();
 DECAPx4_ASAP7_75t_R FILLER_311_85 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_101 ();
 DECAPx10_ASAP7_75t_R FILLER_311_115 ();
 FILLER_ASAP7_75t_R FILLER_311_137 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_154 ();
 DECAPx2_ASAP7_75t_R FILLER_311_164 ();
 FILLER_ASAP7_75t_R FILLER_311_170 ();
 DECAPx1_ASAP7_75t_R FILLER_311_198 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_311_220 ();
 DECAPx1_ASAP7_75t_R FILLER_311_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_233 ();
 FILLER_ASAP7_75t_R FILLER_311_252 ();
 FILLER_ASAP7_75t_R FILLER_311_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_268 ();
 DECAPx10_ASAP7_75t_R FILLER_311_272 ();
 DECAPx1_ASAP7_75t_R FILLER_311_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_304 ();
 DECAPx10_ASAP7_75t_R FILLER_311_331 ();
 DECAPx2_ASAP7_75t_R FILLER_311_379 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_311_385 ();
 DECAPx1_ASAP7_75t_R FILLER_311_422 ();
 DECAPx4_ASAP7_75t_R FILLER_311_434 ();
 FILLER_ASAP7_75t_R FILLER_311_466 ();
 DECAPx6_ASAP7_75t_R FILLER_311_480 ();
 DECAPx2_ASAP7_75t_R FILLER_311_494 ();
 DECAPx10_ASAP7_75t_R FILLER_311_505 ();
 DECAPx6_ASAP7_75t_R FILLER_311_527 ();
 FILLER_ASAP7_75t_R FILLER_311_541 ();
 DECAPx2_ASAP7_75t_R FILLER_311_555 ();
 DECAPx6_ASAP7_75t_R FILLER_311_579 ();
 DECAPx2_ASAP7_75t_R FILLER_311_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_599 ();
 DECAPx2_ASAP7_75t_R FILLER_311_612 ();
 FILLER_ASAP7_75t_R FILLER_311_618 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_311_634 ();
 DECAPx10_ASAP7_75t_R FILLER_311_680 ();
 DECAPx10_ASAP7_75t_R FILLER_311_702 ();
 DECAPx10_ASAP7_75t_R FILLER_311_724 ();
 DECAPx10_ASAP7_75t_R FILLER_311_746 ();
 DECAPx4_ASAP7_75t_R FILLER_311_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_778 ();
 DECAPx6_ASAP7_75t_R FILLER_311_782 ();
 DECAPx1_ASAP7_75t_R FILLER_311_796 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_800 ();
 DECAPx6_ASAP7_75t_R FILLER_311_807 ();
 DECAPx1_ASAP7_75t_R FILLER_311_821 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_835 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_311_842 ();
 DECAPx2_ASAP7_75t_R FILLER_311_918 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_924 ();
 DECAPx2_ASAP7_75t_R FILLER_311_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_311_933 ();
 DECAPx10_ASAP7_75t_R FILLER_312_2 ();
 DECAPx10_ASAP7_75t_R FILLER_312_24 ();
 DECAPx6_ASAP7_75t_R FILLER_312_46 ();
 DECAPx2_ASAP7_75t_R FILLER_312_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_66 ();
 DECAPx1_ASAP7_75t_R FILLER_312_93 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_97 ();
 DECAPx10_ASAP7_75t_R FILLER_312_106 ();
 DECAPx10_ASAP7_75t_R FILLER_312_128 ();
 DECAPx10_ASAP7_75t_R FILLER_312_150 ();
 DECAPx2_ASAP7_75t_R FILLER_312_172 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_197 ();
 DECAPx1_ASAP7_75t_R FILLER_312_230 ();
 DECAPx2_ASAP7_75t_R FILLER_312_240 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_312_246 ();
 DECAPx1_ASAP7_75t_R FILLER_312_307 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_311 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_318 ();
 DECAPx10_ASAP7_75t_R FILLER_312_325 ();
 DECAPx6_ASAP7_75t_R FILLER_312_347 ();
 DECAPx2_ASAP7_75t_R FILLER_312_361 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_367 ();
 DECAPx10_ASAP7_75t_R FILLER_312_371 ();
 DECAPx2_ASAP7_75t_R FILLER_312_393 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_312_399 ();
 DECAPx10_ASAP7_75t_R FILLER_312_405 ();
 DECAPx2_ASAP7_75t_R FILLER_312_430 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_451 ();
 DECAPx6_ASAP7_75t_R FILLER_312_464 ();
 FILLER_ASAP7_75t_R FILLER_312_478 ();
 DECAPx10_ASAP7_75t_R FILLER_312_494 ();
 DECAPx2_ASAP7_75t_R FILLER_312_516 ();
 FILLER_ASAP7_75t_R FILLER_312_522 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_529 ();
 FILLER_ASAP7_75t_R FILLER_312_541 ();
 FILLER_ASAP7_75t_R FILLER_312_569 ();
 DECAPx6_ASAP7_75t_R FILLER_312_586 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_312_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_615 ();
 DECAPx2_ASAP7_75t_R FILLER_312_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_639 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_647 ();
 FILLER_ASAP7_75t_R FILLER_312_656 ();
 DECAPx10_ASAP7_75t_R FILLER_312_675 ();
 DECAPx10_ASAP7_75t_R FILLER_312_697 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_719 ();
 FILLER_ASAP7_75t_R FILLER_312_728 ();
 DECAPx2_ASAP7_75t_R FILLER_312_733 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_312_739 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_748 ();
 DECAPx10_ASAP7_75t_R FILLER_312_755 ();
 DECAPx1_ASAP7_75t_R FILLER_312_777 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_781 ();
 DECAPx10_ASAP7_75t_R FILLER_312_796 ();
 DECAPx1_ASAP7_75t_R FILLER_312_818 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_822 ();
 DECAPx1_ASAP7_75t_R FILLER_312_826 ();
 DECAPx10_ASAP7_75t_R FILLER_312_833 ();
 DECAPx1_ASAP7_75t_R FILLER_312_855 ();
 DECAPx1_ASAP7_75t_R FILLER_312_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_312_933 ();
 DECAPx10_ASAP7_75t_R FILLER_313_2 ();
 DECAPx10_ASAP7_75t_R FILLER_313_24 ();
 DECAPx6_ASAP7_75t_R FILLER_313_46 ();
 DECAPx2_ASAP7_75t_R FILLER_313_60 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_98 ();
 DECAPx1_ASAP7_75t_R FILLER_313_107 ();
 DECAPx2_ASAP7_75t_R FILLER_313_137 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_143 ();
 DECAPx4_ASAP7_75t_R FILLER_313_149 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_159 ();
 DECAPx6_ASAP7_75t_R FILLER_313_171 ();
 FILLER_ASAP7_75t_R FILLER_313_185 ();
 FILLER_ASAP7_75t_R FILLER_313_201 ();
 DECAPx10_ASAP7_75t_R FILLER_313_218 ();
 DECAPx10_ASAP7_75t_R FILLER_313_240 ();
 FILLER_ASAP7_75t_R FILLER_313_262 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_267 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_282 ();
 FILLER_ASAP7_75t_R FILLER_313_330 ();
 DECAPx4_ASAP7_75t_R FILLER_313_358 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_374 ();
 DECAPx10_ASAP7_75t_R FILLER_313_380 ();
 FILLER_ASAP7_75t_R FILLER_313_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_410 ();
 DECAPx1_ASAP7_75t_R FILLER_313_417 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_421 ();
 DECAPx1_ASAP7_75t_R FILLER_313_428 ();
 DECAPx6_ASAP7_75t_R FILLER_313_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_467 ();
 DECAPx4_ASAP7_75t_R FILLER_313_493 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_511 ();
 DECAPx1_ASAP7_75t_R FILLER_313_548 ();
 DECAPx1_ASAP7_75t_R FILLER_313_576 ();
 DECAPx10_ASAP7_75t_R FILLER_313_604 ();
 DECAPx1_ASAP7_75t_R FILLER_313_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_630 ();
 DECAPx6_ASAP7_75t_R FILLER_313_634 ();
 DECAPx2_ASAP7_75t_R FILLER_313_648 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_654 ();
 DECAPx1_ASAP7_75t_R FILLER_313_658 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_662 ();
 DECAPx2_ASAP7_75t_R FILLER_313_666 ();
 FILLER_ASAP7_75t_R FILLER_313_672 ();
 DECAPx2_ASAP7_75t_R FILLER_313_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_686 ();
 DECAPx10_ASAP7_75t_R FILLER_313_690 ();
 DECAPx1_ASAP7_75t_R FILLER_313_712 ();
 FILLER_ASAP7_75t_R FILLER_313_742 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_752 ();
 FILLER_ASAP7_75t_R FILLER_313_763 ();
 FILLER_ASAP7_75t_R FILLER_313_775 ();
 DECAPx1_ASAP7_75t_R FILLER_313_810 ();
 DECAPx10_ASAP7_75t_R FILLER_313_835 ();
 DECAPx1_ASAP7_75t_R FILLER_313_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_861 ();
 DECAPx4_ASAP7_75t_R FILLER_313_886 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_896 ();
 DECAPx4_ASAP7_75t_R FILLER_313_900 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_313_910 ();
 DECAPx1_ASAP7_75t_R FILLER_313_921 ();
 DECAPx2_ASAP7_75t_R FILLER_313_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_313_933 ();
 DECAPx10_ASAP7_75t_R FILLER_314_2 ();
 DECAPx10_ASAP7_75t_R FILLER_314_24 ();
 DECAPx10_ASAP7_75t_R FILLER_314_46 ();
 DECAPx4_ASAP7_75t_R FILLER_314_68 ();
 FILLER_ASAP7_75t_R FILLER_314_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_101 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_314_142 ();
 DECAPx4_ASAP7_75t_R FILLER_314_151 ();
 FILLER_ASAP7_75t_R FILLER_314_161 ();
 DECAPx4_ASAP7_75t_R FILLER_314_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_188 ();
 FILLER_ASAP7_75t_R FILLER_314_197 ();
 DECAPx6_ASAP7_75t_R FILLER_314_205 ();
 DECAPx2_ASAP7_75t_R FILLER_314_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_225 ();
 DECAPx4_ASAP7_75t_R FILLER_314_232 ();
 DECAPx10_ASAP7_75t_R FILLER_314_250 ();
 DECAPx1_ASAP7_75t_R FILLER_314_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_284 ();
 DECAPx1_ASAP7_75t_R FILLER_314_291 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_304 ();
 DECAPx10_ASAP7_75t_R FILLER_314_308 ();
 DECAPx2_ASAP7_75t_R FILLER_314_330 ();
 FILLER_ASAP7_75t_R FILLER_314_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_388 ();
 DECAPx1_ASAP7_75t_R FILLER_314_395 ();
 DECAPx10_ASAP7_75t_R FILLER_314_440 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_314_464 ();
 DECAPx4_ASAP7_75t_R FILLER_314_470 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_314_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_498 ();
 FILLER_ASAP7_75t_R FILLER_314_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_548 ();
 DECAPx4_ASAP7_75t_R FILLER_314_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_579 ();
 DECAPx4_ASAP7_75t_R FILLER_314_608 ();
 FILLER_ASAP7_75t_R FILLER_314_618 ();
 DECAPx10_ASAP7_75t_R FILLER_314_623 ();
 DECAPx6_ASAP7_75t_R FILLER_314_645 ();
 DECAPx2_ASAP7_75t_R FILLER_314_659 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_665 ();
 DECAPx4_ASAP7_75t_R FILLER_314_703 ();
 FILLER_ASAP7_75t_R FILLER_314_713 ();
 FILLER_ASAP7_75t_R FILLER_314_729 ();
 DECAPx2_ASAP7_75t_R FILLER_314_790 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_796 ();
 DECAPx4_ASAP7_75t_R FILLER_314_808 ();
 FILLER_ASAP7_75t_R FILLER_314_828 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_833 ();
 FILLER_ASAP7_75t_R FILLER_314_844 ();
 DECAPx4_ASAP7_75t_R FILLER_314_861 ();
 FILLER_ASAP7_75t_R FILLER_314_871 ();
 DECAPx10_ASAP7_75t_R FILLER_314_879 ();
 DECAPx10_ASAP7_75t_R FILLER_314_901 ();
 DECAPx4_ASAP7_75t_R FILLER_314_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_314_933 ();
 DECAPx10_ASAP7_75t_R FILLER_315_2 ();
 DECAPx10_ASAP7_75t_R FILLER_315_24 ();
 DECAPx10_ASAP7_75t_R FILLER_315_46 ();
 DECAPx4_ASAP7_75t_R FILLER_315_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_78 ();
 FILLER_ASAP7_75t_R FILLER_315_84 ();
 DECAPx10_ASAP7_75t_R FILLER_315_89 ();
 DECAPx4_ASAP7_75t_R FILLER_315_111 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_121 ();
 FILLER_ASAP7_75t_R FILLER_315_125 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_133 ();
 DECAPx10_ASAP7_75t_R FILLER_315_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_184 ();
 DECAPx10_ASAP7_75t_R FILLER_315_197 ();
 FILLER_ASAP7_75t_R FILLER_315_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_234 ();
 DECAPx4_ASAP7_75t_R FILLER_315_242 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_252 ();
 DECAPx10_ASAP7_75t_R FILLER_315_264 ();
 DECAPx10_ASAP7_75t_R FILLER_315_286 ();
 DECAPx6_ASAP7_75t_R FILLER_315_308 ();
 DECAPx10_ASAP7_75t_R FILLER_315_340 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_362 ();
 DECAPx4_ASAP7_75t_R FILLER_315_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_413 ();
 DECAPx10_ASAP7_75t_R FILLER_315_417 ();
 DECAPx2_ASAP7_75t_R FILLER_315_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_456 ();
 DECAPx4_ASAP7_75t_R FILLER_315_479 ();
 FILLER_ASAP7_75t_R FILLER_315_489 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_511 ();
 DECAPx6_ASAP7_75t_R FILLER_315_531 ();
 FILLER_ASAP7_75t_R FILLER_315_545 ();
 DECAPx4_ASAP7_75t_R FILLER_315_557 ();
 DECAPx4_ASAP7_75t_R FILLER_315_573 ();
 DECAPx1_ASAP7_75t_R FILLER_315_589 ();
 DECAPx4_ASAP7_75t_R FILLER_315_599 ();
 DECAPx2_ASAP7_75t_R FILLER_315_623 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_646 ();
 DECAPx6_ASAP7_75t_R FILLER_315_663 ();
 DECAPx2_ASAP7_75t_R FILLER_315_677 ();
 DECAPx10_ASAP7_75t_R FILLER_315_697 ();
 DECAPx2_ASAP7_75t_R FILLER_315_719 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_766 ();
 DECAPx4_ASAP7_75t_R FILLER_315_772 ();
 FILLER_ASAP7_75t_R FILLER_315_782 ();
 FILLER_ASAP7_75t_R FILLER_315_794 ();
 DECAPx10_ASAP7_75t_R FILLER_315_864 ();
 FILLER_ASAP7_75t_R FILLER_315_886 ();
 FILLER_ASAP7_75t_R FILLER_315_894 ();
 DECAPx6_ASAP7_75t_R FILLER_315_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_315_922 ();
 DECAPx2_ASAP7_75t_R FILLER_315_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_315_933 ();
 DECAPx10_ASAP7_75t_R FILLER_316_2 ();
 DECAPx10_ASAP7_75t_R FILLER_316_24 ();
 DECAPx10_ASAP7_75t_R FILLER_316_46 ();
 DECAPx10_ASAP7_75t_R FILLER_316_68 ();
 DECAPx10_ASAP7_75t_R FILLER_316_90 ();
 DECAPx10_ASAP7_75t_R FILLER_316_112 ();
 DECAPx2_ASAP7_75t_R FILLER_316_134 ();
 DECAPx1_ASAP7_75t_R FILLER_316_146 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_150 ();
 DECAPx10_ASAP7_75t_R FILLER_316_154 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_176 ();
 DECAPx10_ASAP7_75t_R FILLER_316_185 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_213 ();
 DECAPx6_ASAP7_75t_R FILLER_316_275 ();
 DECAPx1_ASAP7_75t_R FILLER_316_289 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_300 ();
 DECAPx10_ASAP7_75t_R FILLER_316_307 ();
 DECAPx10_ASAP7_75t_R FILLER_316_329 ();
 DECAPx10_ASAP7_75t_R FILLER_316_351 ();
 DECAPx1_ASAP7_75t_R FILLER_316_373 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_383 ();
 FILLER_ASAP7_75t_R FILLER_316_389 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_408 ();
 DECAPx10_ASAP7_75t_R FILLER_316_423 ();
 DECAPx4_ASAP7_75t_R FILLER_316_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_455 ();
 DECAPx6_ASAP7_75t_R FILLER_316_484 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_518 ();
 DECAPx10_ASAP7_75t_R FILLER_316_526 ();
 DECAPx6_ASAP7_75t_R FILLER_316_548 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_562 ();
 DECAPx10_ASAP7_75t_R FILLER_316_579 ();
 DECAPx2_ASAP7_75t_R FILLER_316_601 ();
 DECAPx1_ASAP7_75t_R FILLER_316_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_628 ();
 FILLER_ASAP7_75t_R FILLER_316_649 ();
 DECAPx6_ASAP7_75t_R FILLER_316_665 ();
 FILLER_ASAP7_75t_R FILLER_316_679 ();
 DECAPx10_ASAP7_75t_R FILLER_316_687 ();
 DECAPx10_ASAP7_75t_R FILLER_316_709 ();
 DECAPx10_ASAP7_75t_R FILLER_316_731 ();
 DECAPx2_ASAP7_75t_R FILLER_316_753 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_759 ();
 DECAPx10_ASAP7_75t_R FILLER_316_767 ();
 DECAPx4_ASAP7_75t_R FILLER_316_789 ();
 FILLERxp5_ASAP7_75t_R FILLER_316_799 ();
 DECAPx10_ASAP7_75t_R FILLER_316_816 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_838 ();
 DECAPx6_ASAP7_75t_R FILLER_316_867 ();
 DECAPx1_ASAP7_75t_R FILLER_316_881 ();
 FILLER_ASAP7_75t_R FILLER_316_911 ();
 DECAPx2_ASAP7_75t_R FILLER_316_925 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_316_931 ();
 DECAPx10_ASAP7_75t_R FILLER_317_2 ();
 DECAPx10_ASAP7_75t_R FILLER_317_24 ();
 DECAPx10_ASAP7_75t_R FILLER_317_46 ();
 DECAPx10_ASAP7_75t_R FILLER_317_68 ();
 DECAPx6_ASAP7_75t_R FILLER_317_90 ();
 DECAPx1_ASAP7_75t_R FILLER_317_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_108 ();
 DECAPx10_ASAP7_75t_R FILLER_317_121 ();
 DECAPx2_ASAP7_75t_R FILLER_317_143 ();
 FILLER_ASAP7_75t_R FILLER_317_149 ();
 DECAPx1_ASAP7_75t_R FILLER_317_163 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_167 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_317_194 ();
 DECAPx1_ASAP7_75t_R FILLER_317_230 ();
 DECAPx2_ASAP7_75t_R FILLER_317_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_288 ();
 DECAPx1_ASAP7_75t_R FILLER_317_318 ();
 DECAPx6_ASAP7_75t_R FILLER_317_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_342 ();
 DECAPx10_ASAP7_75t_R FILLER_317_365 ();
 DECAPx10_ASAP7_75t_R FILLER_317_387 ();
 DECAPx4_ASAP7_75t_R FILLER_317_415 ();
 DECAPx10_ASAP7_75t_R FILLER_317_447 ();
 DECAPx4_ASAP7_75t_R FILLER_317_469 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_317_479 ();
 DECAPx10_ASAP7_75t_R FILLER_317_490 ();
 DECAPx6_ASAP7_75t_R FILLER_317_512 ();
 DECAPx2_ASAP7_75t_R FILLER_317_526 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_532 ();
 FILLER_ASAP7_75t_R FILLER_317_536 ();
 DECAPx4_ASAP7_75t_R FILLER_317_541 ();
 FILLER_ASAP7_75t_R FILLER_317_551 ();
 DECAPx10_ASAP7_75t_R FILLER_317_556 ();
 DECAPx10_ASAP7_75t_R FILLER_317_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_600 ();
 DECAPx2_ASAP7_75t_R FILLER_317_613 ();
 DECAPx1_ASAP7_75t_R FILLER_317_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_640 ();
 DECAPx10_ASAP7_75t_R FILLER_317_658 ();
 DECAPx10_ASAP7_75t_R FILLER_317_680 ();
 DECAPx10_ASAP7_75t_R FILLER_317_702 ();
 DECAPx10_ASAP7_75t_R FILLER_317_724 ();
 DECAPx10_ASAP7_75t_R FILLER_317_746 ();
 DECAPx1_ASAP7_75t_R FILLER_317_768 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_772 ();
 DECAPx10_ASAP7_75t_R FILLER_317_781 ();
 DECAPx2_ASAP7_75t_R FILLER_317_803 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_809 ();
 DECAPx10_ASAP7_75t_R FILLER_317_820 ();
 DECAPx4_ASAP7_75t_R FILLER_317_842 ();
 DECAPx4_ASAP7_75t_R FILLER_317_883 ();
 FILLERxp5_ASAP7_75t_R FILLER_317_906 ();
 FILLER_ASAP7_75t_R FILLER_317_923 ();
 DECAPx1_ASAP7_75t_R FILLER_317_930 ();
 DECAPx10_ASAP7_75t_R FILLER_318_2 ();
 DECAPx10_ASAP7_75t_R FILLER_318_24 ();
 DECAPx10_ASAP7_75t_R FILLER_318_46 ();
 DECAPx2_ASAP7_75t_R FILLER_318_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_74 ();
 FILLER_ASAP7_75t_R FILLER_318_89 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_101 ();
 DECAPx2_ASAP7_75t_R FILLER_318_128 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_134 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_143 ();
 FILLER_ASAP7_75t_R FILLER_318_181 ();
 DECAPx6_ASAP7_75t_R FILLER_318_186 ();
 DECAPx1_ASAP7_75t_R FILLER_318_200 ();
 FILLER_ASAP7_75t_R FILLER_318_210 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_215 ();
 DECAPx2_ASAP7_75t_R FILLER_318_219 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_225 ();
 DECAPx1_ASAP7_75t_R FILLER_318_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_245 ();
 DECAPx4_ASAP7_75t_R FILLER_318_254 ();
 FILLER_ASAP7_75t_R FILLER_318_264 ();
 FILLER_ASAP7_75t_R FILLER_318_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_300 ();
 FILLER_ASAP7_75t_R FILLER_318_307 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_323 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_346 ();
 DECAPx2_ASAP7_75t_R FILLER_318_375 ();
 FILLER_ASAP7_75t_R FILLER_318_381 ();
 DECAPx10_ASAP7_75t_R FILLER_318_389 ();
 DECAPx4_ASAP7_75t_R FILLER_318_411 ();
 FILLER_ASAP7_75t_R FILLER_318_421 ();
 DECAPx1_ASAP7_75t_R FILLER_318_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_433 ();
 DECAPx2_ASAP7_75t_R FILLER_318_446 ();
 FILLER_ASAP7_75t_R FILLER_318_452 ();
 FILLER_ASAP7_75t_R FILLER_318_460 ();
 DECAPx6_ASAP7_75t_R FILLER_318_464 ();
 DECAPx2_ASAP7_75t_R FILLER_318_478 ();
 DECAPx10_ASAP7_75t_R FILLER_318_492 ();
 DECAPx2_ASAP7_75t_R FILLER_318_514 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_520 ();
 FILLER_ASAP7_75t_R FILLER_318_530 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_535 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_564 ();
 DECAPx2_ASAP7_75t_R FILLER_318_584 ();
 FILLER_ASAP7_75t_R FILLER_318_590 ();
 DECAPx4_ASAP7_75t_R FILLER_318_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_605 ();
 DECAPx4_ASAP7_75t_R FILLER_318_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_628 ();
 DECAPx10_ASAP7_75t_R FILLER_318_632 ();
 DECAPx4_ASAP7_75t_R FILLER_318_654 ();
 FILLER_ASAP7_75t_R FILLER_318_664 ();
 DECAPx10_ASAP7_75t_R FILLER_318_688 ();
 DECAPx10_ASAP7_75t_R FILLER_318_710 ();
 DECAPx1_ASAP7_75t_R FILLER_318_732 ();
 DECAPx4_ASAP7_75t_R FILLER_318_748 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_758 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_769 ();
 FILLER_ASAP7_75t_R FILLER_318_782 ();
 DECAPx10_ASAP7_75t_R FILLER_318_797 ();
 DECAPx10_ASAP7_75t_R FILLER_318_819 ();
 DECAPx10_ASAP7_75t_R FILLER_318_841 ();
 DECAPx4_ASAP7_75t_R FILLER_318_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_318_873 ();
 DECAPx6_ASAP7_75t_R FILLER_318_877 ();
 FILLER_ASAP7_75t_R FILLER_318_891 ();
 DECAPx2_ASAP7_75t_R FILLER_318_899 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_318_905 ();
 DECAPx10_ASAP7_75t_R FILLER_319_2 ();
 DECAPx10_ASAP7_75t_R FILLER_319_24 ();
 DECAPx10_ASAP7_75t_R FILLER_319_46 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_68 ();
 FILLER_ASAP7_75t_R FILLER_319_95 ();
 DECAPx1_ASAP7_75t_R FILLER_319_120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_319_127 ();
 DECAPx10_ASAP7_75t_R FILLER_319_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_160 ();
 DECAPx10_ASAP7_75t_R FILLER_319_164 ();
 FILLER_ASAP7_75t_R FILLER_319_186 ();
 DECAPx10_ASAP7_75t_R FILLER_319_204 ();
 DECAPx10_ASAP7_75t_R FILLER_319_226 ();
 DECAPx4_ASAP7_75t_R FILLER_319_248 ();
 DECAPx4_ASAP7_75t_R FILLER_319_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_321 ();
 FILLER_ASAP7_75t_R FILLER_319_354 ();
 DECAPx2_ASAP7_75t_R FILLER_319_396 ();
 DECAPx6_ASAP7_75t_R FILLER_319_408 ();
 FILLER_ASAP7_75t_R FILLER_319_422 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_430 ();
 FILLER_ASAP7_75t_R FILLER_319_457 ();
 DECAPx1_ASAP7_75t_R FILLER_319_465 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_477 ();
 DECAPx4_ASAP7_75t_R FILLER_319_484 ();
 FILLER_ASAP7_75t_R FILLER_319_494 ();
 FILLER_ASAP7_75t_R FILLER_319_524 ();
 FILLER_ASAP7_75t_R FILLER_319_582 ();
 DECAPx4_ASAP7_75t_R FILLER_319_598 ();
 DECAPx2_ASAP7_75t_R FILLER_319_632 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_319_638 ();
 DECAPx4_ASAP7_75t_R FILLER_319_644 ();
 FILLER_ASAP7_75t_R FILLER_319_654 ();
 DECAPx6_ASAP7_75t_R FILLER_319_704 ();
 DECAPx2_ASAP7_75t_R FILLER_319_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_768 ();
 DECAPx10_ASAP7_75t_R FILLER_319_795 ();
 DECAPx2_ASAP7_75t_R FILLER_319_817 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_319_823 ();
 DECAPx10_ASAP7_75t_R FILLER_319_842 ();
 DECAPx2_ASAP7_75t_R FILLER_319_864 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_319_870 ();
 DECAPx1_ASAP7_75t_R FILLER_319_882 ();
 DECAPx10_ASAP7_75t_R FILLER_319_892 ();
 DECAPx4_ASAP7_75t_R FILLER_319_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_924 ();
 DECAPx2_ASAP7_75t_R FILLER_319_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_319_933 ();
 DECAPx10_ASAP7_75t_R FILLER_320_2 ();
 DECAPx10_ASAP7_75t_R FILLER_320_24 ();
 DECAPx10_ASAP7_75t_R FILLER_320_46 ();
 DECAPx6_ASAP7_75t_R FILLER_320_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_91 ();
 DECAPx1_ASAP7_75t_R FILLER_320_106 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_110 ();
 DECAPx6_ASAP7_75t_R FILLER_320_143 ();
 DECAPx1_ASAP7_75t_R FILLER_320_157 ();
 DECAPx2_ASAP7_75t_R FILLER_320_181 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_187 ();
 DECAPx10_ASAP7_75t_R FILLER_320_202 ();
 DECAPx10_ASAP7_75t_R FILLER_320_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_261 ();
 DECAPx1_ASAP7_75t_R FILLER_320_268 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_272 ();
 DECAPx10_ASAP7_75t_R FILLER_320_279 ();
 FILLER_ASAP7_75t_R FILLER_320_301 ();
 FILLER_ASAP7_75t_R FILLER_320_309 ();
 DECAPx6_ASAP7_75t_R FILLER_320_317 ();
 DECAPx10_ASAP7_75t_R FILLER_320_340 ();
 FILLER_ASAP7_75t_R FILLER_320_389 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_401 ();
 FILLER_ASAP7_75t_R FILLER_320_418 ();
 DECAPx6_ASAP7_75t_R FILLER_320_432 ();
 DECAPx1_ASAP7_75t_R FILLER_320_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_450 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_459 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_464 ();
 DECAPx2_ASAP7_75t_R FILLER_320_471 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_477 ();
 DECAPx6_ASAP7_75t_R FILLER_320_486 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_500 ();
 DECAPx2_ASAP7_75t_R FILLER_320_523 ();
 DECAPx1_ASAP7_75t_R FILLER_320_532 ();
 DECAPx4_ASAP7_75t_R FILLER_320_539 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_549 ();
 DECAPx1_ASAP7_75t_R FILLER_320_555 ();
 DECAPx2_ASAP7_75t_R FILLER_320_562 ();
 FILLER_ASAP7_75t_R FILLER_320_568 ();
 DECAPx2_ASAP7_75t_R FILLER_320_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_579 ();
 DECAPx2_ASAP7_75t_R FILLER_320_586 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_592 ();
 DECAPx2_ASAP7_75t_R FILLER_320_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_604 ();
 DECAPx2_ASAP7_75t_R FILLER_320_617 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_320_623 ();
 DECAPx6_ASAP7_75t_R FILLER_320_640 ();
 FILLER_ASAP7_75t_R FILLER_320_668 ();
 FILLER_ASAP7_75t_R FILLER_320_681 ();
 DECAPx10_ASAP7_75t_R FILLER_320_691 ();
 FILLER_ASAP7_75t_R FILLER_320_713 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_742 ();
 DECAPx2_ASAP7_75t_R FILLER_320_746 ();
 FILLER_ASAP7_75t_R FILLER_320_752 ();
 DECAPx1_ASAP7_75t_R FILLER_320_763 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_767 ();
 DECAPx6_ASAP7_75t_R FILLER_320_780 ();
 FILLER_ASAP7_75t_R FILLER_320_794 ();
 DECAPx2_ASAP7_75t_R FILLER_320_811 ();
 DECAPx10_ASAP7_75t_R FILLER_320_849 ();
 FILLER_ASAP7_75t_R FILLER_320_871 ();
 DECAPx10_ASAP7_75t_R FILLER_320_905 ();
 DECAPx2_ASAP7_75t_R FILLER_320_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_320_933 ();
 DECAPx10_ASAP7_75t_R FILLER_321_2 ();
 DECAPx10_ASAP7_75t_R FILLER_321_24 ();
 DECAPx10_ASAP7_75t_R FILLER_321_46 ();
 FILLER_ASAP7_75t_R FILLER_321_68 ();
 DECAPx4_ASAP7_75t_R FILLER_321_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_106 ();
 DECAPx1_ASAP7_75t_R FILLER_321_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_137 ();
 DECAPx4_ASAP7_75t_R FILLER_321_152 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_162 ();
 DECAPx6_ASAP7_75t_R FILLER_321_195 ();
 DECAPx1_ASAP7_75t_R FILLER_321_209 ();
 DECAPx1_ASAP7_75t_R FILLER_321_221 ();
 FILLER_ASAP7_75t_R FILLER_321_237 ();
 DECAPx10_ASAP7_75t_R FILLER_321_271 ();
 DECAPx10_ASAP7_75t_R FILLER_321_293 ();
 DECAPx10_ASAP7_75t_R FILLER_321_315 ();
 DECAPx10_ASAP7_75t_R FILLER_321_337 ();
 DECAPx1_ASAP7_75t_R FILLER_321_359 ();
 FILLER_ASAP7_75t_R FILLER_321_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_321_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_443 ();
 DECAPx4_ASAP7_75t_R FILLER_321_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_459 ();
 DECAPx4_ASAP7_75t_R FILLER_321_466 ();
 FILLER_ASAP7_75t_R FILLER_321_476 ();
 DECAPx4_ASAP7_75t_R FILLER_321_498 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_321_508 ();
 DECAPx10_ASAP7_75t_R FILLER_321_517 ();
 DECAPx6_ASAP7_75t_R FILLER_321_539 ();
 FILLER_ASAP7_75t_R FILLER_321_553 ();
 DECAPx2_ASAP7_75t_R FILLER_321_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_321_575 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_321_598 ();
 DECAPx10_ASAP7_75t_R FILLER_321_613 ();
 FILLER_ASAP7_75t_R FILLER_321_635 ();
 DECAPx4_ASAP7_75t_R FILLER_321_666 ();
 DECAPx10_ASAP7_75t_R FILLER_321_682 ();
 DECAPx6_ASAP7_75t_R FILLER_321_704 ();
 DECAPx10_ASAP7_75t_R FILLER_321_744 ();
 DECAPx4_ASAP7_75t_R FILLER_321_766 ();
 FILLER_ASAP7_75t_R FILLER_321_776 ();
 DECAPx1_ASAP7_75t_R FILLER_321_799 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_803 ();
 DECAPx2_ASAP7_75t_R FILLER_321_820 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_321_826 ();
 DECAPx6_ASAP7_75t_R FILLER_321_845 ();
 DECAPx1_ASAP7_75t_R FILLER_321_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_863 ();
 DECAPx6_ASAP7_75t_R FILLER_321_890 ();
 FILLER_ASAP7_75t_R FILLER_321_904 ();
 DECAPx4_ASAP7_75t_R FILLER_321_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_924 ();
 DECAPx2_ASAP7_75t_R FILLER_321_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_321_933 ();
 DECAPx10_ASAP7_75t_R FILLER_322_2 ();
 DECAPx10_ASAP7_75t_R FILLER_322_24 ();
 DECAPx10_ASAP7_75t_R FILLER_322_46 ();
 DECAPx2_ASAP7_75t_R FILLER_322_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_74 ();
 FILLER_ASAP7_75t_R FILLER_322_83 ();
 DECAPx10_ASAP7_75t_R FILLER_322_88 ();
 DECAPx4_ASAP7_75t_R FILLER_322_110 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_120 ();
 DECAPx4_ASAP7_75t_R FILLER_322_124 ();
 FILLER_ASAP7_75t_R FILLER_322_134 ();
 DECAPx4_ASAP7_75t_R FILLER_322_162 ();
 FILLER_ASAP7_75t_R FILLER_322_172 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_223 ();
 DECAPx1_ASAP7_75t_R FILLER_322_246 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_250 ();
 FILLER_ASAP7_75t_R FILLER_322_257 ();
 DECAPx6_ASAP7_75t_R FILLER_322_262 ();
 DECAPx2_ASAP7_75t_R FILLER_322_276 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_288 ();
 DECAPx10_ASAP7_75t_R FILLER_322_294 ();
 DECAPx6_ASAP7_75t_R FILLER_322_316 ();
 DECAPx2_ASAP7_75t_R FILLER_322_330 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_336 ();
 DECAPx4_ASAP7_75t_R FILLER_322_344 ();
 FILLER_ASAP7_75t_R FILLER_322_354 ();
 DECAPx6_ASAP7_75t_R FILLER_322_382 ();
 FILLER_ASAP7_75t_R FILLER_322_396 ();
 DECAPx4_ASAP7_75t_R FILLER_322_406 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_416 ();
 DECAPx10_ASAP7_75t_R FILLER_322_436 ();
 DECAPx1_ASAP7_75t_R FILLER_322_458 ();
 DECAPx4_ASAP7_75t_R FILLER_322_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_474 ();
 DECAPx6_ASAP7_75t_R FILLER_322_495 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_518 ();
 DECAPx10_ASAP7_75t_R FILLER_322_543 ();
 DECAPx1_ASAP7_75t_R FILLER_322_565 ();
 DECAPx2_ASAP7_75t_R FILLER_322_575 ();
 FILLER_ASAP7_75t_R FILLER_322_581 ();
 DECAPx2_ASAP7_75t_R FILLER_322_589 ();
 DECAPx6_ASAP7_75t_R FILLER_322_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_615 ();
 FILLER_ASAP7_75t_R FILLER_322_627 ();
 FILLER_ASAP7_75t_R FILLER_322_633 ();
 DECAPx10_ASAP7_75t_R FILLER_322_642 ();
 DECAPx4_ASAP7_75t_R FILLER_322_664 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_674 ();
 DECAPx10_ASAP7_75t_R FILLER_322_692 ();
 DECAPx6_ASAP7_75t_R FILLER_322_714 ();
 DECAPx1_ASAP7_75t_R FILLER_322_728 ();
 DECAPx10_ASAP7_75t_R FILLER_322_735 ();
 DECAPx10_ASAP7_75t_R FILLER_322_757 ();
 DECAPx10_ASAP7_75t_R FILLER_322_779 ();
 DECAPx4_ASAP7_75t_R FILLER_322_833 ();
 DECAPx4_ASAP7_75t_R FILLER_322_867 ();
 FILLERxp5_ASAP7_75t_R FILLER_322_877 ();
 DECAPx6_ASAP7_75t_R FILLER_322_881 ();
 FILLER_ASAP7_75t_R FILLER_322_895 ();
 DECAPx2_ASAP7_75t_R FILLER_322_925 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_322_931 ();
 DECAPx10_ASAP7_75t_R FILLER_323_2 ();
 DECAPx10_ASAP7_75t_R FILLER_323_24 ();
 DECAPx10_ASAP7_75t_R FILLER_323_46 ();
 DECAPx10_ASAP7_75t_R FILLER_323_68 ();
 DECAPx10_ASAP7_75t_R FILLER_323_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_112 ();
 DECAPx10_ASAP7_75t_R FILLER_323_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_144 ();
 DECAPx2_ASAP7_75t_R FILLER_323_173 ();
 DECAPx1_ASAP7_75t_R FILLER_323_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_224 ();
 DECAPx2_ASAP7_75t_R FILLER_323_231 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_237 ();
 DECAPx10_ASAP7_75t_R FILLER_323_246 ();
 DECAPx2_ASAP7_75t_R FILLER_323_268 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_274 ();
 DECAPx1_ASAP7_75t_R FILLER_323_306 ();
 DECAPx1_ASAP7_75t_R FILLER_323_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_320 ();
 DECAPx1_ASAP7_75t_R FILLER_323_332 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_348 ();
 DECAPx1_ASAP7_75t_R FILLER_323_357 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_367 ();
 DECAPx10_ASAP7_75t_R FILLER_323_373 ();
 DECAPx4_ASAP7_75t_R FILLER_323_405 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_415 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_430 ();
 DECAPx4_ASAP7_75t_R FILLER_323_434 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_444 ();
 DECAPx10_ASAP7_75t_R FILLER_323_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_492 ();
 DECAPx1_ASAP7_75t_R FILLER_323_496 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_517 ();
 DECAPx2_ASAP7_75t_R FILLER_323_534 ();
 FILLER_ASAP7_75t_R FILLER_323_540 ();
 DECAPx1_ASAP7_75t_R FILLER_323_545 ();
 DECAPx1_ASAP7_75t_R FILLER_323_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_556 ();
 DECAPx4_ASAP7_75t_R FILLER_323_560 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_570 ();
 DECAPx2_ASAP7_75t_R FILLER_323_577 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_583 ();
 DECAPx2_ASAP7_75t_R FILLER_323_611 ();
 FILLER_ASAP7_75t_R FILLER_323_617 ();
 DECAPx2_ASAP7_75t_R FILLER_323_649 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_655 ();
 DECAPx10_ASAP7_75t_R FILLER_323_661 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_683 ();
 DECAPx10_ASAP7_75t_R FILLER_323_687 ();
 DECAPx10_ASAP7_75t_R FILLER_323_709 ();
 DECAPx10_ASAP7_75t_R FILLER_323_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_753 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_760 ();
 DECAPx6_ASAP7_75t_R FILLER_323_769 ();
 FILLER_ASAP7_75t_R FILLER_323_783 ();
 DECAPx1_ASAP7_75t_R FILLER_323_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_801 ();
 DECAPx2_ASAP7_75t_R FILLER_323_828 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_323_834 ();
 FILLER_ASAP7_75t_R FILLER_323_849 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_863 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_877 ();
 DECAPx2_ASAP7_75t_R FILLER_323_885 ();
 FILLER_ASAP7_75t_R FILLER_323_891 ();
 FILLER_ASAP7_75t_R FILLER_323_908 ();
 DECAPx2_ASAP7_75t_R FILLER_323_919 ();
 DECAPx2_ASAP7_75t_R FILLER_323_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_323_933 ();
 DECAPx10_ASAP7_75t_R FILLER_324_2 ();
 DECAPx10_ASAP7_75t_R FILLER_324_24 ();
 DECAPx10_ASAP7_75t_R FILLER_324_46 ();
 DECAPx10_ASAP7_75t_R FILLER_324_68 ();
 DECAPx2_ASAP7_75t_R FILLER_324_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_96 ();
 DECAPx4_ASAP7_75t_R FILLER_324_134 ();
 FILLER_ASAP7_75t_R FILLER_324_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_155 ();
 DECAPx10_ASAP7_75t_R FILLER_324_162 ();
 FILLER_ASAP7_75t_R FILLER_324_184 ();
 DECAPx1_ASAP7_75t_R FILLER_324_196 ();
 DECAPx1_ASAP7_75t_R FILLER_324_215 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_219 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_324_226 ();
 DECAPx6_ASAP7_75t_R FILLER_324_256 ();
 DECAPx1_ASAP7_75t_R FILLER_324_270 ();
 DECAPx1_ASAP7_75t_R FILLER_324_294 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_325 ();
 FILLER_ASAP7_75t_R FILLER_324_334 ();
 DECAPx10_ASAP7_75t_R FILLER_324_356 ();
 DECAPx6_ASAP7_75t_R FILLER_324_378 ();
 DECAPx4_ASAP7_75t_R FILLER_324_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_435 ();
 DECAPx6_ASAP7_75t_R FILLER_324_479 ();
 FILLER_ASAP7_75t_R FILLER_324_521 ();
 DECAPx4_ASAP7_75t_R FILLER_324_529 ();
 FILLER_ASAP7_75t_R FILLER_324_539 ();
 DECAPx2_ASAP7_75t_R FILLER_324_558 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_324_564 ();
 DECAPx6_ASAP7_75t_R FILLER_324_581 ();
 FILLER_ASAP7_75t_R FILLER_324_595 ();
 DECAPx10_ASAP7_75t_R FILLER_324_603 ();
 DECAPx10_ASAP7_75t_R FILLER_324_625 ();
 DECAPx10_ASAP7_75t_R FILLER_324_647 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_669 ();
 DECAPx2_ASAP7_75t_R FILLER_324_673 ();
 DECAPx10_ASAP7_75t_R FILLER_324_688 ();
 DECAPx6_ASAP7_75t_R FILLER_324_710 ();
 DECAPx1_ASAP7_75t_R FILLER_324_724 ();
 DECAPx2_ASAP7_75t_R FILLER_324_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_760 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_771 ();
 DECAPx1_ASAP7_75t_R FILLER_324_782 ();
 DECAPx4_ASAP7_75t_R FILLER_324_804 ();
 FILLER_ASAP7_75t_R FILLER_324_814 ();
 DECAPx2_ASAP7_75t_R FILLER_324_825 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_831 ();
 DECAPx2_ASAP7_75t_R FILLER_324_844 ();
 FILLER_ASAP7_75t_R FILLER_324_861 ();
 DECAPx10_ASAP7_75t_R FILLER_324_889 ();
 DECAPx10_ASAP7_75t_R FILLER_324_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_324_933 ();
 DECAPx10_ASAP7_75t_R FILLER_325_2 ();
 DECAPx10_ASAP7_75t_R FILLER_325_24 ();
 DECAPx10_ASAP7_75t_R FILLER_325_46 ();
 DECAPx10_ASAP7_75t_R FILLER_325_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_90 ();
 FILLER_ASAP7_75t_R FILLER_325_107 ();
 DECAPx10_ASAP7_75t_R FILLER_325_115 ();
 DECAPx10_ASAP7_75t_R FILLER_325_137 ();
 DECAPx10_ASAP7_75t_R FILLER_325_159 ();
 DECAPx2_ASAP7_75t_R FILLER_325_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_187 ();
 DECAPx10_ASAP7_75t_R FILLER_325_199 ();
 DECAPx6_ASAP7_75t_R FILLER_325_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_235 ();
 DECAPx2_ASAP7_75t_R FILLER_325_250 ();
 FILLER_ASAP7_75t_R FILLER_325_265 ();
 FILLER_ASAP7_75t_R FILLER_325_278 ();
 FILLER_ASAP7_75t_R FILLER_325_286 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_311 ();
 DECAPx4_ASAP7_75t_R FILLER_325_351 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_361 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_370 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_390 ();
 DECAPx4_ASAP7_75t_R FILLER_325_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_415 ();
 DECAPx2_ASAP7_75t_R FILLER_325_435 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_441 ();
 DECAPx6_ASAP7_75t_R FILLER_325_464 ();
 DECAPx1_ASAP7_75t_R FILLER_325_478 ();
 DECAPx1_ASAP7_75t_R FILLER_325_496 ();
 FILLER_ASAP7_75t_R FILLER_325_506 ();
 DECAPx10_ASAP7_75t_R FILLER_325_511 ();
 FILLER_ASAP7_75t_R FILLER_325_533 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_538 ();
 DECAPx1_ASAP7_75t_R FILLER_325_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_548 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_552 ();
 DECAPx6_ASAP7_75t_R FILLER_325_556 ();
 FILLER_ASAP7_75t_R FILLER_325_570 ();
 DECAPx6_ASAP7_75t_R FILLER_325_575 ();
 FILLER_ASAP7_75t_R FILLER_325_589 ();
 DECAPx6_ASAP7_75t_R FILLER_325_594 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_608 ();
 DECAPx6_ASAP7_75t_R FILLER_325_620 ();
 DECAPx2_ASAP7_75t_R FILLER_325_634 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_647 ();
 DECAPx6_ASAP7_75t_R FILLER_325_664 ();
 DECAPx1_ASAP7_75t_R FILLER_325_678 ();
 DECAPx10_ASAP7_75t_R FILLER_325_696 ();
 DECAPx1_ASAP7_75t_R FILLER_325_718 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_757 ();
 DECAPx6_ASAP7_75t_R FILLER_325_784 ();
 DECAPx10_ASAP7_75t_R FILLER_325_808 ();
 DECAPx10_ASAP7_75t_R FILLER_325_838 ();
 DECAPx2_ASAP7_75t_R FILLER_325_860 ();
 DECAPx2_ASAP7_75t_R FILLER_325_872 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_881 ();
 DECAPx2_ASAP7_75t_R FILLER_325_892 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_325_907 ();
 DECAPx2_ASAP7_75t_R FILLER_325_917 ();
 FILLER_ASAP7_75t_R FILLER_325_923 ();
 DECAPx2_ASAP7_75t_R FILLER_325_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_325_933 ();
 DECAPx10_ASAP7_75t_R FILLER_326_2 ();
 DECAPx10_ASAP7_75t_R FILLER_326_24 ();
 DECAPx10_ASAP7_75t_R FILLER_326_46 ();
 DECAPx4_ASAP7_75t_R FILLER_326_68 ();
 FILLER_ASAP7_75t_R FILLER_326_78 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_92 ();
 DECAPx10_ASAP7_75t_R FILLER_326_104 ();
 DECAPx10_ASAP7_75t_R FILLER_326_126 ();
 DECAPx10_ASAP7_75t_R FILLER_326_148 ();
 DECAPx2_ASAP7_75t_R FILLER_326_170 ();
 FILLER_ASAP7_75t_R FILLER_326_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_204 ();
 DECAPx4_ASAP7_75t_R FILLER_326_211 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_221 ();
 DECAPx10_ASAP7_75t_R FILLER_326_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_247 ();
 DECAPx2_ASAP7_75t_R FILLER_326_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_288 ();
 DECAPx4_ASAP7_75t_R FILLER_326_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_305 ();
 DECAPx6_ASAP7_75t_R FILLER_326_318 ();
 DECAPx6_ASAP7_75t_R FILLER_326_338 ();
 DECAPx1_ASAP7_75t_R FILLER_326_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_356 ();
 DECAPx4_ASAP7_75t_R FILLER_326_419 ();
 FILLER_ASAP7_75t_R FILLER_326_429 ();
 DECAPx1_ASAP7_75t_R FILLER_326_441 ();
 DECAPx4_ASAP7_75t_R FILLER_326_450 ();
 FILLER_ASAP7_75t_R FILLER_326_460 ();
 DECAPx2_ASAP7_75t_R FILLER_326_464 ();
 FILLER_ASAP7_75t_R FILLER_326_470 ();
 DECAPx10_ASAP7_75t_R FILLER_326_482 ();
 DECAPx10_ASAP7_75t_R FILLER_326_504 ();
 FILLER_ASAP7_75t_R FILLER_326_529 ();
 DECAPx6_ASAP7_75t_R FILLER_326_534 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_548 ();
 DECAPx2_ASAP7_75t_R FILLER_326_563 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_569 ();
 DECAPx2_ASAP7_75t_R FILLER_326_575 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_581 ();
 DECAPx10_ASAP7_75t_R FILLER_326_590 ();
 DECAPx6_ASAP7_75t_R FILLER_326_612 ();
 FILLER_ASAP7_75t_R FILLER_326_626 ();
 DECAPx2_ASAP7_75t_R FILLER_326_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_655 ();
 DECAPx4_ASAP7_75t_R FILLER_326_673 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_689 ();
 DECAPx10_ASAP7_75t_R FILLER_326_695 ();
 DECAPx2_ASAP7_75t_R FILLER_326_717 ();
 FILLER_ASAP7_75t_R FILLER_326_758 ();
 FILLER_ASAP7_75t_R FILLER_326_781 ();
 DECAPx10_ASAP7_75t_R FILLER_326_809 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_831 ();
 DECAPx2_ASAP7_75t_R FILLER_326_840 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_326_846 ();
 DECAPx10_ASAP7_75t_R FILLER_326_862 ();
 DECAPx6_ASAP7_75t_R FILLER_326_884 ();
 FILLERxp5_ASAP7_75t_R FILLER_326_901 ();
 DECAPx10_ASAP7_75t_R FILLER_327_2 ();
 DECAPx10_ASAP7_75t_R FILLER_327_24 ();
 DECAPx10_ASAP7_75t_R FILLER_327_46 ();
 DECAPx1_ASAP7_75t_R FILLER_327_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_72 ();
 DECAPx6_ASAP7_75t_R FILLER_327_99 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_113 ();
 FILLER_ASAP7_75t_R FILLER_327_122 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_152 ();
 DECAPx1_ASAP7_75t_R FILLER_327_158 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_180 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_189 ();
 DECAPx4_ASAP7_75t_R FILLER_327_221 ();
 DECAPx2_ASAP7_75t_R FILLER_327_243 ();
 FILLER_ASAP7_75t_R FILLER_327_249 ();
 DECAPx1_ASAP7_75t_R FILLER_327_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_261 ();
 DECAPx1_ASAP7_75t_R FILLER_327_296 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_300 ();
 DECAPx4_ASAP7_75t_R FILLER_327_327 ();
 DECAPx1_ASAP7_75t_R FILLER_327_343 ();
 FILLER_ASAP7_75t_R FILLER_327_350 ();
 DECAPx2_ASAP7_75t_R FILLER_327_355 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_367 ();
 FILLER_ASAP7_75t_R FILLER_327_387 ();
 DECAPx6_ASAP7_75t_R FILLER_327_415 ();
 DECAPx1_ASAP7_75t_R FILLER_327_429 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_433 ();
 DECAPx10_ASAP7_75t_R FILLER_327_446 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_468 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_490 ();
 FILLER_ASAP7_75t_R FILLER_327_504 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_509 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_518 ();
 DECAPx2_ASAP7_75t_R FILLER_327_552 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_558 ();
 FILLER_ASAP7_75t_R FILLER_327_564 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_580 ();
 DECAPx6_ASAP7_75t_R FILLER_327_595 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_609 ();
 DECAPx4_ASAP7_75t_R FILLER_327_624 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_634 ();
 DECAPx6_ASAP7_75t_R FILLER_327_644 ();
 FILLER_ASAP7_75t_R FILLER_327_658 ();
 DECAPx10_ASAP7_75t_R FILLER_327_674 ();
 DECAPx10_ASAP7_75t_R FILLER_327_696 ();
 DECAPx2_ASAP7_75t_R FILLER_327_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_724 ();
 DECAPx10_ASAP7_75t_R FILLER_327_757 ();
 DECAPx6_ASAP7_75t_R FILLER_327_779 ();
 DECAPx1_ASAP7_75t_R FILLER_327_793 ();
 DECAPx10_ASAP7_75t_R FILLER_327_800 ();
 DECAPx2_ASAP7_75t_R FILLER_327_822 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_828 ();
 FILLER_ASAP7_75t_R FILLER_327_838 ();
 DECAPx1_ASAP7_75t_R FILLER_327_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_327_854 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_327_864 ();
 DECAPx4_ASAP7_75t_R FILLER_327_877 ();
 FILLER_ASAP7_75t_R FILLER_327_887 ();
 DECAPx1_ASAP7_75t_R FILLER_327_930 ();
 DECAPx10_ASAP7_75t_R FILLER_328_2 ();
 DECAPx10_ASAP7_75t_R FILLER_328_24 ();
 DECAPx10_ASAP7_75t_R FILLER_328_46 ();
 DECAPx6_ASAP7_75t_R FILLER_328_68 ();
 DECAPx2_ASAP7_75t_R FILLER_328_82 ();
 DECAPx6_ASAP7_75t_R FILLER_328_91 ();
 DECAPx2_ASAP7_75t_R FILLER_328_105 ();
 DECAPx1_ASAP7_75t_R FILLER_328_127 ();
 FILLER_ASAP7_75t_R FILLER_328_137 ();
 DECAPx6_ASAP7_75t_R FILLER_328_179 ();
 DECAPx2_ASAP7_75t_R FILLER_328_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_199 ();
 DECAPx1_ASAP7_75t_R FILLER_328_206 ();
 FILLER_ASAP7_75t_R FILLER_328_213 ();
 DECAPx1_ASAP7_75t_R FILLER_328_223 ();
 DECAPx1_ASAP7_75t_R FILLER_328_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_237 ();
 DECAPx1_ASAP7_75t_R FILLER_328_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_256 ();
 DECAPx6_ASAP7_75t_R FILLER_328_266 ();
 DECAPx1_ASAP7_75t_R FILLER_328_280 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_290 ();
 DECAPx6_ASAP7_75t_R FILLER_328_300 ();
 FILLER_ASAP7_75t_R FILLER_328_314 ();
 DECAPx2_ASAP7_75t_R FILLER_328_319 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_325 ();
 DECAPx10_ASAP7_75t_R FILLER_328_358 ();
 DECAPx4_ASAP7_75t_R FILLER_328_380 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_328_390 ();
 DECAPx6_ASAP7_75t_R FILLER_328_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_422 ();
 DECAPx6_ASAP7_75t_R FILLER_328_443 ();
 DECAPx1_ASAP7_75t_R FILLER_328_457 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_461 ();
 FILLER_ASAP7_75t_R FILLER_328_479 ();
 DECAPx4_ASAP7_75t_R FILLER_328_491 ();
 FILLER_ASAP7_75t_R FILLER_328_501 ();
 DECAPx10_ASAP7_75t_R FILLER_328_523 ();
 DECAPx2_ASAP7_75t_R FILLER_328_545 ();
 DECAPx4_ASAP7_75t_R FILLER_328_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_581 ();
 DECAPx1_ASAP7_75t_R FILLER_328_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_595 ();
 DECAPx2_ASAP7_75t_R FILLER_328_607 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_328_613 ();
 DECAPx1_ASAP7_75t_R FILLER_328_625 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_629 ();
 DECAPx2_ASAP7_75t_R FILLER_328_653 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_659 ();
 DECAPx2_ASAP7_75t_R FILLER_328_683 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_328_689 ();
 DECAPx10_ASAP7_75t_R FILLER_328_695 ();
 DECAPx6_ASAP7_75t_R FILLER_328_717 ();
 DECAPx2_ASAP7_75t_R FILLER_328_731 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_737 ();
 DECAPx10_ASAP7_75t_R FILLER_328_741 ();
 DECAPx4_ASAP7_75t_R FILLER_328_763 ();
 DECAPx10_ASAP7_75t_R FILLER_328_779 ();
 DECAPx4_ASAP7_75t_R FILLER_328_801 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_328_811 ();
 DECAPx1_ASAP7_75t_R FILLER_328_824 ();
 FILLER_ASAP7_75t_R FILLER_328_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_328_882 ();
 DECAPx6_ASAP7_75t_R FILLER_328_897 ();
 DECAPx1_ASAP7_75t_R FILLER_328_911 ();
 DECAPx6_ASAP7_75t_R FILLER_328_918 ();
 FILLER_ASAP7_75t_R FILLER_328_932 ();
 DECAPx10_ASAP7_75t_R FILLER_329_2 ();
 DECAPx10_ASAP7_75t_R FILLER_329_24 ();
 DECAPx10_ASAP7_75t_R FILLER_329_46 ();
 DECAPx10_ASAP7_75t_R FILLER_329_68 ();
 DECAPx6_ASAP7_75t_R FILLER_329_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_113 ();
 FILLER_ASAP7_75t_R FILLER_329_123 ();
 DECAPx2_ASAP7_75t_R FILLER_329_137 ();
 DECAPx1_ASAP7_75t_R FILLER_329_149 ();
 DECAPx10_ASAP7_75t_R FILLER_329_164 ();
 DECAPx2_ASAP7_75t_R FILLER_329_186 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_192 ();
 DECAPx2_ASAP7_75t_R FILLER_329_205 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_211 ();
 DECAPx1_ASAP7_75t_R FILLER_329_275 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_279 ();
 DECAPx1_ASAP7_75t_R FILLER_329_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_310 ();
 DECAPx6_ASAP7_75t_R FILLER_329_317 ();
 DECAPx1_ASAP7_75t_R FILLER_329_331 ();
 FILLER_ASAP7_75t_R FILLER_329_361 ();
 DECAPx10_ASAP7_75t_R FILLER_329_369 ();
 DECAPx6_ASAP7_75t_R FILLER_329_391 ();
 DECAPx1_ASAP7_75t_R FILLER_329_405 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_409 ();
 DECAPx1_ASAP7_75t_R FILLER_329_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_443 ();
 DECAPx10_ASAP7_75t_R FILLER_329_480 ();
 DECAPx4_ASAP7_75t_R FILLER_329_502 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_512 ();
 DECAPx2_ASAP7_75t_R FILLER_329_528 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_329_537 ();
 DECAPx6_ASAP7_75t_R FILLER_329_543 ();
 DECAPx1_ASAP7_75t_R FILLER_329_557 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_561 ();
 DECAPx10_ASAP7_75t_R FILLER_329_565 ();
 DECAPx6_ASAP7_75t_R FILLER_329_587 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_329_601 ();
 FILLER_ASAP7_75t_R FILLER_329_626 ();
 DECAPx4_ASAP7_75t_R FILLER_329_638 ();
 FILLER_ASAP7_75t_R FILLER_329_648 ();
 DECAPx2_ASAP7_75t_R FILLER_329_664 ();
 FILLER_ASAP7_75t_R FILLER_329_684 ();
 DECAPx10_ASAP7_75t_R FILLER_329_703 ();
 DECAPx10_ASAP7_75t_R FILLER_329_725 ();
 DECAPx10_ASAP7_75t_R FILLER_329_747 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_769 ();
 DECAPx1_ASAP7_75t_R FILLER_329_787 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_791 ();
 FILLER_ASAP7_75t_R FILLER_329_804 ();
 DECAPx1_ASAP7_75t_R FILLER_329_832 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_842 ();
 DECAPx4_ASAP7_75t_R FILLER_329_846 ();
 DECAPx1_ASAP7_75t_R FILLER_329_859 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_869 ();
 FILLER_ASAP7_75t_R FILLER_329_879 ();
 DECAPx6_ASAP7_75t_R FILLER_329_907 ();
 DECAPx1_ASAP7_75t_R FILLER_329_921 ();
 DECAPx2_ASAP7_75t_R FILLER_329_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_329_933 ();
 DECAPx10_ASAP7_75t_R FILLER_330_2 ();
 DECAPx10_ASAP7_75t_R FILLER_330_24 ();
 DECAPx10_ASAP7_75t_R FILLER_330_46 ();
 DECAPx6_ASAP7_75t_R FILLER_330_68 ();
 FILLER_ASAP7_75t_R FILLER_330_82 ();
 DECAPx10_ASAP7_75t_R FILLER_330_116 ();
 DECAPx6_ASAP7_75t_R FILLER_330_138 ();
 FILLER_ASAP7_75t_R FILLER_330_152 ();
 DECAPx10_ASAP7_75t_R FILLER_330_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_188 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_215 ();
 DECAPx1_ASAP7_75t_R FILLER_330_228 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_232 ();
 DECAPx1_ASAP7_75t_R FILLER_330_248 ();
 DECAPx10_ASAP7_75t_R FILLER_330_258 ();
 DECAPx6_ASAP7_75t_R FILLER_330_280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_330_294 ();
 DECAPx2_ASAP7_75t_R FILLER_330_334 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_356 ();
 DECAPx1_ASAP7_75t_R FILLER_330_389 ();
 DECAPx2_ASAP7_75t_R FILLER_330_396 ();
 FILLER_ASAP7_75t_R FILLER_330_402 ();
 FILLER_ASAP7_75t_R FILLER_330_410 ();
 DECAPx4_ASAP7_75t_R FILLER_330_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_467 ();
 DECAPx10_ASAP7_75t_R FILLER_330_503 ();
 DECAPx1_ASAP7_75t_R FILLER_330_525 ();
 DECAPx10_ASAP7_75t_R FILLER_330_562 ();
 DECAPx4_ASAP7_75t_R FILLER_330_584 ();
 FILLER_ASAP7_75t_R FILLER_330_608 ();
 DECAPx10_ASAP7_75t_R FILLER_330_622 ();
 DECAPx6_ASAP7_75t_R FILLER_330_644 ();
 FILLER_ASAP7_75t_R FILLER_330_658 ();
 DECAPx10_ASAP7_75t_R FILLER_330_663 ();
 FILLER_ASAP7_75t_R FILLER_330_685 ();
 DECAPx10_ASAP7_75t_R FILLER_330_704 ();
 DECAPx10_ASAP7_75t_R FILLER_330_726 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_330_748 ();
 DECAPx6_ASAP7_75t_R FILLER_330_757 ();
 DECAPx2_ASAP7_75t_R FILLER_330_771 ();
 FILLERxp5_ASAP7_75t_R FILLER_330_777 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_330_810 ();
 DECAPx10_ASAP7_75t_R FILLER_330_831 ();
 DECAPx10_ASAP7_75t_R FILLER_330_853 ();
 DECAPx4_ASAP7_75t_R FILLER_330_875 ();
 FILLER_ASAP7_75t_R FILLER_330_885 ();
 DECAPx10_ASAP7_75t_R FILLER_330_909 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_330_931 ();
 DECAPx10_ASAP7_75t_R FILLER_331_2 ();
 DECAPx10_ASAP7_75t_R FILLER_331_24 ();
 DECAPx10_ASAP7_75t_R FILLER_331_46 ();
 DECAPx4_ASAP7_75t_R FILLER_331_68 ();
 DECAPx1_ASAP7_75t_R FILLER_331_110 ();
 DECAPx6_ASAP7_75t_R FILLER_331_126 ();
 DECAPx2_ASAP7_75t_R FILLER_331_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_146 ();
 DECAPx2_ASAP7_75t_R FILLER_331_159 ();
 FILLER_ASAP7_75t_R FILLER_331_165 ();
 DECAPx4_ASAP7_75t_R FILLER_331_193 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_203 ();
 DECAPx10_ASAP7_75t_R FILLER_331_207 ();
 DECAPx10_ASAP7_75t_R FILLER_331_229 ();
 DECAPx2_ASAP7_75t_R FILLER_331_251 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_257 ();
 DECAPx6_ASAP7_75t_R FILLER_331_266 ();
 FILLER_ASAP7_75t_R FILLER_331_280 ();
 DECAPx6_ASAP7_75t_R FILLER_331_288 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_302 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_309 ();
 DECAPx4_ASAP7_75t_R FILLER_331_315 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_325 ();
 DECAPx10_ASAP7_75t_R FILLER_331_336 ();
 FILLER_ASAP7_75t_R FILLER_331_358 ();
 FILLER_ASAP7_75t_R FILLER_331_366 ();
 DECAPx6_ASAP7_75t_R FILLER_331_430 ();
 DECAPx2_ASAP7_75t_R FILLER_331_444 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_450 ();
 DECAPx2_ASAP7_75t_R FILLER_331_469 ();
 DECAPx6_ASAP7_75t_R FILLER_331_495 ();
 DECAPx4_ASAP7_75t_R FILLER_331_523 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_533 ();
 DECAPx2_ASAP7_75t_R FILLER_331_537 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_543 ();
 DECAPx6_ASAP7_75t_R FILLER_331_558 ();
 DECAPx1_ASAP7_75t_R FILLER_331_572 ();
 DECAPx10_ASAP7_75t_R FILLER_331_579 ();
 DECAPx6_ASAP7_75t_R FILLER_331_615 ();
 FILLER_ASAP7_75t_R FILLER_331_629 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_640 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_657 ();
 DECAPx1_ASAP7_75t_R FILLER_331_685 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_689 ();
 DECAPx10_ASAP7_75t_R FILLER_331_696 ();
 DECAPx1_ASAP7_75t_R FILLER_331_718 ();
 FILLER_ASAP7_75t_R FILLER_331_754 ();
 DECAPx4_ASAP7_75t_R FILLER_331_772 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_331_782 ();
 DECAPx6_ASAP7_75t_R FILLER_331_807 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_824 ();
 DECAPx10_ASAP7_75t_R FILLER_331_828 ();
 DECAPx2_ASAP7_75t_R FILLER_331_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_856 ();
 DECAPx10_ASAP7_75t_R FILLER_331_863 ();
 DECAPx4_ASAP7_75t_R FILLER_331_885 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_895 ();
 DECAPx10_ASAP7_75t_R FILLER_331_899 ();
 DECAPx1_ASAP7_75t_R FILLER_331_921 ();
 DECAPx2_ASAP7_75t_R FILLER_331_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_331_933 ();
 DECAPx10_ASAP7_75t_R FILLER_332_2 ();
 DECAPx10_ASAP7_75t_R FILLER_332_24 ();
 DECAPx10_ASAP7_75t_R FILLER_332_46 ();
 DECAPx6_ASAP7_75t_R FILLER_332_68 ();
 DECAPx2_ASAP7_75t_R FILLER_332_82 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_88 ();
 DECAPx4_ASAP7_75t_R FILLER_332_98 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_108 ();
 DECAPx1_ASAP7_75t_R FILLER_332_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_139 ();
 DECAPx1_ASAP7_75t_R FILLER_332_195 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_199 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_206 ();
 DECAPx10_ASAP7_75t_R FILLER_332_213 ();
 DECAPx6_ASAP7_75t_R FILLER_332_235 ();
 FILLER_ASAP7_75t_R FILLER_332_249 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_306 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_315 ();
 DECAPx1_ASAP7_75t_R FILLER_332_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_326 ();
 DECAPx10_ASAP7_75t_R FILLER_332_339 ();
 DECAPx4_ASAP7_75t_R FILLER_332_361 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_380 ();
 DECAPx6_ASAP7_75t_R FILLER_332_386 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_400 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_407 ();
 DECAPx4_ASAP7_75t_R FILLER_332_411 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_421 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_427 ();
 DECAPx6_ASAP7_75t_R FILLER_332_433 ();
 DECAPx1_ASAP7_75t_R FILLER_332_447 ();
 DECAPx2_ASAP7_75t_R FILLER_332_456 ();
 DECAPx6_ASAP7_75t_R FILLER_332_464 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_486 ();
 DECAPx4_ASAP7_75t_R FILLER_332_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_506 ();
 DECAPx10_ASAP7_75t_R FILLER_332_521 ();
 DECAPx6_ASAP7_75t_R FILLER_332_543 ();
 DECAPx1_ASAP7_75t_R FILLER_332_569 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_573 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_588 ();
 DECAPx10_ASAP7_75t_R FILLER_332_616 ();
 DECAPx6_ASAP7_75t_R FILLER_332_638 ();
 DECAPx1_ASAP7_75t_R FILLER_332_669 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_673 ();
 DECAPx10_ASAP7_75t_R FILLER_332_694 ();
 DECAPx6_ASAP7_75t_R FILLER_332_716 ();
 DECAPx2_ASAP7_75t_R FILLER_332_730 ();
 FILLER_ASAP7_75t_R FILLER_332_739 ();
 DECAPx10_ASAP7_75t_R FILLER_332_777 ();
 DECAPx4_ASAP7_75t_R FILLER_332_799 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_809 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_332_821 ();
 DECAPx2_ASAP7_75t_R FILLER_332_833 ();
 DECAPx1_ASAP7_75t_R FILLER_332_871 ();
 FILLERxp5_ASAP7_75t_R FILLER_332_875 ();
 DECAPx10_ASAP7_75t_R FILLER_332_882 ();
 DECAPx10_ASAP7_75t_R FILLER_332_904 ();
 DECAPx2_ASAP7_75t_R FILLER_332_926 ();
 FILLER_ASAP7_75t_R FILLER_332_932 ();
 DECAPx10_ASAP7_75t_R FILLER_333_2 ();
 DECAPx10_ASAP7_75t_R FILLER_333_24 ();
 DECAPx10_ASAP7_75t_R FILLER_333_46 ();
 DECAPx10_ASAP7_75t_R FILLER_333_68 ();
 DECAPx6_ASAP7_75t_R FILLER_333_90 ();
 DECAPx6_ASAP7_75t_R FILLER_333_110 ();
 DECAPx1_ASAP7_75t_R FILLER_333_153 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_157 ();
 DECAPx4_ASAP7_75t_R FILLER_333_161 ();
 FILLER_ASAP7_75t_R FILLER_333_171 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_179 ();
 DECAPx4_ASAP7_75t_R FILLER_333_183 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_333_193 ();
 DECAPx1_ASAP7_75t_R FILLER_333_222 ();
 DECAPx2_ASAP7_75t_R FILLER_333_252 ();
 DECAPx2_ASAP7_75t_R FILLER_333_261 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_267 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_333_277 ();
 DECAPx2_ASAP7_75t_R FILLER_333_286 ();
 DECAPx4_ASAP7_75t_R FILLER_333_295 ();
 DECAPx4_ASAP7_75t_R FILLER_333_331 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_333_341 ();
 DECAPx10_ASAP7_75t_R FILLER_333_360 ();
 DECAPx10_ASAP7_75t_R FILLER_333_382 ();
 DECAPx1_ASAP7_75t_R FILLER_333_404 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_443 ();
 DECAPx10_ASAP7_75t_R FILLER_333_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_472 ();
 DECAPx4_ASAP7_75t_R FILLER_333_516 ();
 DECAPx10_ASAP7_75t_R FILLER_333_535 ();
 FILLER_ASAP7_75t_R FILLER_333_568 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_576 ();
 DECAPx2_ASAP7_75t_R FILLER_333_621 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_627 ();
 DECAPx10_ASAP7_75t_R FILLER_333_631 ();
 DECAPx10_ASAP7_75t_R FILLER_333_653 ();
 DECAPx1_ASAP7_75t_R FILLER_333_675 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_679 ();
 DECAPx10_ASAP7_75t_R FILLER_333_686 ();
 DECAPx10_ASAP7_75t_R FILLER_333_708 ();
 DECAPx6_ASAP7_75t_R FILLER_333_730 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_756 ();
 DECAPx4_ASAP7_75t_R FILLER_333_772 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_782 ();
 DECAPx6_ASAP7_75t_R FILLER_333_786 ();
 DECAPx1_ASAP7_75t_R FILLER_333_800 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_804 ();
 DECAPx10_ASAP7_75t_R FILLER_333_811 ();
 DECAPx1_ASAP7_75t_R FILLER_333_833 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_837 ();
 DECAPx1_ASAP7_75t_R FILLER_333_861 ();
 DECAPx10_ASAP7_75t_R FILLER_333_893 ();
 DECAPx4_ASAP7_75t_R FILLER_333_915 ();
 DECAPx2_ASAP7_75t_R FILLER_333_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_333_933 ();
 DECAPx10_ASAP7_75t_R FILLER_334_2 ();
 DECAPx10_ASAP7_75t_R FILLER_334_24 ();
 DECAPx10_ASAP7_75t_R FILLER_334_46 ();
 DECAPx10_ASAP7_75t_R FILLER_334_68 ();
 DECAPx1_ASAP7_75t_R FILLER_334_90 ();
 DECAPx4_ASAP7_75t_R FILLER_334_120 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_130 ();
 DECAPx10_ASAP7_75t_R FILLER_334_151 ();
 DECAPx6_ASAP7_75t_R FILLER_334_173 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_187 ();
 DECAPx6_ASAP7_75t_R FILLER_334_194 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_208 ();
 DECAPx2_ASAP7_75t_R FILLER_334_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_220 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_228 ();
 DECAPx10_ASAP7_75t_R FILLER_334_269 ();
 DECAPx10_ASAP7_75t_R FILLER_334_291 ();
 DECAPx2_ASAP7_75t_R FILLER_334_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_319 ();
 DECAPx6_ASAP7_75t_R FILLER_334_323 ();
 FILLER_ASAP7_75t_R FILLER_334_337 ();
 DECAPx2_ASAP7_75t_R FILLER_334_365 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_371 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_380 ();
 DECAPx10_ASAP7_75t_R FILLER_334_387 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_409 ();
 DECAPx2_ASAP7_75t_R FILLER_334_453 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_459 ();
 DECAPx4_ASAP7_75t_R FILLER_334_464 ();
 FILLER_ASAP7_75t_R FILLER_334_474 ();
 FILLER_ASAP7_75t_R FILLER_334_493 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_513 ();
 DECAPx4_ASAP7_75t_R FILLER_334_522 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_532 ();
 DECAPx2_ASAP7_75t_R FILLER_334_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_593 ();
 DECAPx1_ASAP7_75t_R FILLER_334_603 ();
 FILLER_ASAP7_75t_R FILLER_334_630 ();
 DECAPx10_ASAP7_75t_R FILLER_334_646 ();
 DECAPx10_ASAP7_75t_R FILLER_334_671 ();
 DECAPx10_ASAP7_75t_R FILLER_334_693 ();
 DECAPx10_ASAP7_75t_R FILLER_334_715 ();
 DECAPx10_ASAP7_75t_R FILLER_334_737 ();
 DECAPx4_ASAP7_75t_R FILLER_334_759 ();
 DECAPx6_ASAP7_75t_R FILLER_334_795 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_809 ();
 FILLER_ASAP7_75t_R FILLER_334_829 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_839 ();
 DECAPx10_ASAP7_75t_R FILLER_334_848 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_334_870 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_885 ();
 DECAPx1_ASAP7_75t_R FILLER_334_904 ();
 FILLERxp5_ASAP7_75t_R FILLER_334_908 ();
 DECAPx10_ASAP7_75t_R FILLER_334_912 ();
 DECAPx10_ASAP7_75t_R FILLER_335_2 ();
 DECAPx10_ASAP7_75t_R FILLER_335_24 ();
 DECAPx10_ASAP7_75t_R FILLER_335_46 ();
 DECAPx10_ASAP7_75t_R FILLER_335_68 ();
 DECAPx2_ASAP7_75t_R FILLER_335_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_335_96 ();
 DECAPx1_ASAP7_75t_R FILLER_335_105 ();
 DECAPx10_ASAP7_75t_R FILLER_335_112 ();
 DECAPx10_ASAP7_75t_R FILLER_335_134 ();
 DECAPx10_ASAP7_75t_R FILLER_335_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_335_178 ();
 DECAPx4_ASAP7_75t_R FILLER_335_207 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_217 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_250 ();
 DECAPx6_ASAP7_75t_R FILLER_335_257 ();
 DECAPx2_ASAP7_75t_R FILLER_335_271 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_277 ();
 DECAPx2_ASAP7_75t_R FILLER_335_290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_335_296 ();
 FILLER_ASAP7_75t_R FILLER_335_305 ();
 DECAPx6_ASAP7_75t_R FILLER_335_310 ();
 DECAPx1_ASAP7_75t_R FILLER_335_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_328 ();
 DECAPx2_ASAP7_75t_R FILLER_335_364 ();
 DECAPx2_ASAP7_75t_R FILLER_335_396 ();
 DECAPx2_ASAP7_75t_R FILLER_335_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_414 ();
 FILLER_ASAP7_75t_R FILLER_335_431 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_454 ();
 FILLER_ASAP7_75t_R FILLER_335_461 ();
 FILLER_ASAP7_75t_R FILLER_335_466 ();
 DECAPx2_ASAP7_75t_R FILLER_335_529 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_535 ();
 DECAPx10_ASAP7_75t_R FILLER_335_579 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_601 ();
 DECAPx2_ASAP7_75t_R FILLER_335_608 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_634 ();
 DECAPx2_ASAP7_75t_R FILLER_335_658 ();
 DECAPx2_ASAP7_75t_R FILLER_335_686 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_692 ();
 DECAPx10_ASAP7_75t_R FILLER_335_696 ();
 DECAPx10_ASAP7_75t_R FILLER_335_718 ();
 DECAPx10_ASAP7_75t_R FILLER_335_740 ();
 DECAPx4_ASAP7_75t_R FILLER_335_762 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_772 ();
 DECAPx2_ASAP7_75t_R FILLER_335_789 ();
 DECAPx1_ASAP7_75t_R FILLER_335_801 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_805 ();
 DECAPx6_ASAP7_75t_R FILLER_335_840 ();
 DECAPx1_ASAP7_75t_R FILLER_335_854 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_858 ();
 FILLER_ASAP7_75t_R FILLER_335_887 ();
 DECAPx1_ASAP7_75t_R FILLER_335_921 ();
 DECAPx2_ASAP7_75t_R FILLER_335_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_335_933 ();
 DECAPx10_ASAP7_75t_R FILLER_336_2 ();
 DECAPx10_ASAP7_75t_R FILLER_336_24 ();
 DECAPx10_ASAP7_75t_R FILLER_336_46 ();
 DECAPx10_ASAP7_75t_R FILLER_336_68 ();
 DECAPx10_ASAP7_75t_R FILLER_336_90 ();
 DECAPx10_ASAP7_75t_R FILLER_336_112 ();
 DECAPx6_ASAP7_75t_R FILLER_336_134 ();
 DECAPx2_ASAP7_75t_R FILLER_336_148 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_154 ();
 DECAPx1_ASAP7_75t_R FILLER_336_167 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_171 ();
 DECAPx4_ASAP7_75t_R FILLER_336_175 ();
 DECAPx1_ASAP7_75t_R FILLER_336_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_195 ();
 DECAPx10_ASAP7_75t_R FILLER_336_199 ();
 DECAPx1_ASAP7_75t_R FILLER_336_221 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_225 ();
 DECAPx6_ASAP7_75t_R FILLER_336_235 ();
 DECAPx1_ASAP7_75t_R FILLER_336_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_253 ();
 DECAPx2_ASAP7_75t_R FILLER_336_257 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_263 ();
 DECAPx2_ASAP7_75t_R FILLER_336_270 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_336_290 ();
 DECAPx6_ASAP7_75t_R FILLER_336_319 ();
 DECAPx2_ASAP7_75t_R FILLER_336_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_339 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_336_346 ();
 DECAPx4_ASAP7_75t_R FILLER_336_352 ();
 DECAPx4_ASAP7_75t_R FILLER_336_374 ();
 FILLER_ASAP7_75t_R FILLER_336_387 ();
 DECAPx1_ASAP7_75t_R FILLER_336_404 ();
 DECAPx2_ASAP7_75t_R FILLER_336_414 ();
 FILLER_ASAP7_75t_R FILLER_336_420 ();
 DECAPx6_ASAP7_75t_R FILLER_336_433 ();
 DECAPx2_ASAP7_75t_R FILLER_336_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_453 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_461 ();
 DECAPx10_ASAP7_75t_R FILLER_336_496 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_527 ();
 DECAPx4_ASAP7_75t_R FILLER_336_551 ();
 FILLER_ASAP7_75t_R FILLER_336_561 ();
 DECAPx10_ASAP7_75t_R FILLER_336_569 ();
 DECAPx6_ASAP7_75t_R FILLER_336_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_605 ();
 FILLER_ASAP7_75t_R FILLER_336_634 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_678 ();
 DECAPx10_ASAP7_75t_R FILLER_336_691 ();
 DECAPx10_ASAP7_75t_R FILLER_336_713 ();
 DECAPx10_ASAP7_75t_R FILLER_336_735 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_757 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_336_766 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_772 ();
 DECAPx4_ASAP7_75t_R FILLER_336_785 ();
 DECAPx2_ASAP7_75t_R FILLER_336_811 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_817 ();
 DECAPx2_ASAP7_75t_R FILLER_336_844 ();
 DECAPx2_ASAP7_75t_R FILLER_336_885 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_336_891 ();
 DECAPx10_ASAP7_75t_R FILLER_336_901 ();
 DECAPx4_ASAP7_75t_R FILLER_336_923 ();
 FILLERxp5_ASAP7_75t_R FILLER_336_933 ();
 DECAPx10_ASAP7_75t_R FILLER_337_2 ();
 DECAPx10_ASAP7_75t_R FILLER_337_24 ();
 DECAPx10_ASAP7_75t_R FILLER_337_46 ();
 DECAPx10_ASAP7_75t_R FILLER_337_68 ();
 DECAPx6_ASAP7_75t_R FILLER_337_90 ();
 FILLER_ASAP7_75t_R FILLER_337_104 ();
 FILLER_ASAP7_75t_R FILLER_337_141 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_149 ();
 DECAPx4_ASAP7_75t_R FILLER_337_190 ();
 DECAPx10_ASAP7_75t_R FILLER_337_209 ();
 DECAPx10_ASAP7_75t_R FILLER_337_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_337_253 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_264 ();
 FILLER_ASAP7_75t_R FILLER_337_271 ();
 DECAPx2_ASAP7_75t_R FILLER_337_279 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_285 ();
 FILLER_ASAP7_75t_R FILLER_337_294 ();
 DECAPx2_ASAP7_75t_R FILLER_337_302 ();
 FILLER_ASAP7_75t_R FILLER_337_308 ();
 FILLER_ASAP7_75t_R FILLER_337_316 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_324 ();
 DECAPx10_ASAP7_75t_R FILLER_337_331 ();
 DECAPx2_ASAP7_75t_R FILLER_337_353 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_337_402 ();
 DECAPx10_ASAP7_75t_R FILLER_337_421 ();
 DECAPx1_ASAP7_75t_R FILLER_337_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_447 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_474 ();
 DECAPx10_ASAP7_75t_R FILLER_337_485 ();
 DECAPx4_ASAP7_75t_R FILLER_337_507 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_337_517 ();
 DECAPx10_ASAP7_75t_R FILLER_337_534 ();
 DECAPx6_ASAP7_75t_R FILLER_337_556 ();
 FILLER_ASAP7_75t_R FILLER_337_570 ();
 DECAPx2_ASAP7_75t_R FILLER_337_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_584 ();
 DECAPx10_ASAP7_75t_R FILLER_337_597 ();
 DECAPx10_ASAP7_75t_R FILLER_337_619 ();
 DECAPx2_ASAP7_75t_R FILLER_337_641 ();
 DECAPx1_ASAP7_75t_R FILLER_337_661 ();
 DECAPx1_ASAP7_75t_R FILLER_337_678 ();
 DECAPx10_ASAP7_75t_R FILLER_337_696 ();
 DECAPx10_ASAP7_75t_R FILLER_337_718 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_337_740 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_337_784 ();
 DECAPx6_ASAP7_75t_R FILLER_337_813 ();
 DECAPx1_ASAP7_75t_R FILLER_337_827 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_831 ();
 DECAPx10_ASAP7_75t_R FILLER_337_835 ();
 DECAPx1_ASAP7_75t_R FILLER_337_857 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_861 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_874 ();
 DECAPx10_ASAP7_75t_R FILLER_337_885 ();
 DECAPx6_ASAP7_75t_R FILLER_337_907 ();
 DECAPx1_ASAP7_75t_R FILLER_337_921 ();
 DECAPx2_ASAP7_75t_R FILLER_337_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_337_933 ();
 DECAPx10_ASAP7_75t_R FILLER_338_2 ();
 DECAPx10_ASAP7_75t_R FILLER_338_24 ();
 DECAPx10_ASAP7_75t_R FILLER_338_46 ();
 DECAPx10_ASAP7_75t_R FILLER_338_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_338_90 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_181 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_190 ();
 DECAPx1_ASAP7_75t_R FILLER_338_220 ();
 DECAPx2_ASAP7_75t_R FILLER_338_230 ();
 DECAPx2_ASAP7_75t_R FILLER_338_242 ();
 FILLER_ASAP7_75t_R FILLER_338_248 ();
 DECAPx4_ASAP7_75t_R FILLER_338_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_266 ();
 DECAPx6_ASAP7_75t_R FILLER_338_275 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_338_289 ();
 DECAPx2_ASAP7_75t_R FILLER_338_298 ();
 FILLER_ASAP7_75t_R FILLER_338_304 ();
 DECAPx2_ASAP7_75t_R FILLER_338_338 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_344 ();
 DECAPx10_ASAP7_75t_R FILLER_338_351 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_373 ();
 DECAPx1_ASAP7_75t_R FILLER_338_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_381 ();
 DECAPx6_ASAP7_75t_R FILLER_338_388 ();
 DECAPx2_ASAP7_75t_R FILLER_338_402 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_338_415 ();
 DECAPx4_ASAP7_75t_R FILLER_338_440 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_461 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_464 ();
 DECAPx4_ASAP7_75t_R FILLER_338_477 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_487 ();
 DECAPx2_ASAP7_75t_R FILLER_338_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_338_500 ();
 DECAPx10_ASAP7_75t_R FILLER_338_518 ();
 DECAPx4_ASAP7_75t_R FILLER_338_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_550 ();
 DECAPx6_ASAP7_75t_R FILLER_338_554 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_568 ();
 DECAPx1_ASAP7_75t_R FILLER_338_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_593 ();
 DECAPx10_ASAP7_75t_R FILLER_338_608 ();
 DECAPx10_ASAP7_75t_R FILLER_338_630 ();
 DECAPx6_ASAP7_75t_R FILLER_338_652 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_338_666 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_674 ();
 DECAPx2_ASAP7_75t_R FILLER_338_678 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_690 ();
 DECAPx10_ASAP7_75t_R FILLER_338_694 ();
 DECAPx10_ASAP7_75t_R FILLER_338_716 ();
 DECAPx6_ASAP7_75t_R FILLER_338_738 ();
 DECAPx2_ASAP7_75t_R FILLER_338_752 ();
 DECAPx10_ASAP7_75t_R FILLER_338_769 ();
 DECAPx1_ASAP7_75t_R FILLER_338_791 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_795 ();
 DECAPx10_ASAP7_75t_R FILLER_338_811 ();
 DECAPx4_ASAP7_75t_R FILLER_338_833 ();
 FILLER_ASAP7_75t_R FILLER_338_843 ();
 DECAPx10_ASAP7_75t_R FILLER_338_851 ();
 DECAPx1_ASAP7_75t_R FILLER_338_873 ();
 FILLERxp5_ASAP7_75t_R FILLER_338_877 ();
 DECAPx10_ASAP7_75t_R FILLER_338_904 ();
 DECAPx2_ASAP7_75t_R FILLER_338_926 ();
 FILLER_ASAP7_75t_R FILLER_338_932 ();
 DECAPx10_ASAP7_75t_R FILLER_339_2 ();
 DECAPx10_ASAP7_75t_R FILLER_339_24 ();
 DECAPx10_ASAP7_75t_R FILLER_339_46 ();
 DECAPx6_ASAP7_75t_R FILLER_339_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_82 ();
 FILLER_ASAP7_75t_R FILLER_339_114 ();
 FILLER_ASAP7_75t_R FILLER_339_130 ();
 DECAPx1_ASAP7_75t_R FILLER_339_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_142 ();
 FILLER_ASAP7_75t_R FILLER_339_152 ();
 DECAPx4_ASAP7_75t_R FILLER_339_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_167 ();
 DECAPx2_ASAP7_75t_R FILLER_339_187 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_193 ();
 DECAPx4_ASAP7_75t_R FILLER_339_202 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_271 ();
 DECAPx4_ASAP7_75t_R FILLER_339_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_292 ();
 DECAPx6_ASAP7_75t_R FILLER_339_299 ();
 DECAPx2_ASAP7_75t_R FILLER_339_313 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_319 ();
 DECAPx2_ASAP7_75t_R FILLER_339_323 ();
 FILLER_ASAP7_75t_R FILLER_339_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_367 ();
 DECAPx2_ASAP7_75t_R FILLER_339_376 ();
 FILLER_ASAP7_75t_R FILLER_339_382 ();
 DECAPx6_ASAP7_75t_R FILLER_339_400 ();
 DECAPx1_ASAP7_75t_R FILLER_339_414 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_418 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_456 ();
 DECAPx4_ASAP7_75t_R FILLER_339_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_479 ();
 DECAPx10_ASAP7_75t_R FILLER_339_519 ();
 DECAPx4_ASAP7_75t_R FILLER_339_541 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_551 ();
 DECAPx6_ASAP7_75t_R FILLER_339_555 ();
 DECAPx1_ASAP7_75t_R FILLER_339_569 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_579 ();
 FILLER_ASAP7_75t_R FILLER_339_596 ();
 FILLER_ASAP7_75t_R FILLER_339_601 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_339_623 ();
 DECAPx1_ASAP7_75t_R FILLER_339_632 ();
 DECAPx6_ASAP7_75t_R FILLER_339_639 ();
 FILLER_ASAP7_75t_R FILLER_339_653 ();
 DECAPx10_ASAP7_75t_R FILLER_339_658 ();
 DECAPx1_ASAP7_75t_R FILLER_339_680 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_684 ();
 DECAPx10_ASAP7_75t_R FILLER_339_702 ();
 DECAPx10_ASAP7_75t_R FILLER_339_724 ();
 DECAPx10_ASAP7_75t_R FILLER_339_746 ();
 DECAPx4_ASAP7_75t_R FILLER_339_768 ();
 FILLER_ASAP7_75t_R FILLER_339_778 ();
 DECAPx10_ASAP7_75t_R FILLER_339_786 ();
 DECAPx4_ASAP7_75t_R FILLER_339_808 ();
 DECAPx1_ASAP7_75t_R FILLER_339_824 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_828 ();
 DECAPx10_ASAP7_75t_R FILLER_339_860 ();
 DECAPx4_ASAP7_75t_R FILLER_339_882 ();
 DECAPx10_ASAP7_75t_R FILLER_339_895 ();
 DECAPx2_ASAP7_75t_R FILLER_339_917 ();
 FILLER_ASAP7_75t_R FILLER_339_923 ();
 DECAPx2_ASAP7_75t_R FILLER_339_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_339_933 ();
 DECAPx10_ASAP7_75t_R FILLER_340_2 ();
 DECAPx10_ASAP7_75t_R FILLER_340_24 ();
 DECAPx10_ASAP7_75t_R FILLER_340_46 ();
 DECAPx10_ASAP7_75t_R FILLER_340_68 ();
 DECAPx2_ASAP7_75t_R FILLER_340_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_96 ();
 DECAPx10_ASAP7_75t_R FILLER_340_108 ();
 DECAPx10_ASAP7_75t_R FILLER_340_130 ();
 DECAPx6_ASAP7_75t_R FILLER_340_152 ();
 DECAPx2_ASAP7_75t_R FILLER_340_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_172 ();
 DECAPx4_ASAP7_75t_R FILLER_340_179 ();
 FILLER_ASAP7_75t_R FILLER_340_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_197 ();
 DECAPx1_ASAP7_75t_R FILLER_340_204 ();
 DECAPx1_ASAP7_75t_R FILLER_340_222 ();
 DECAPx2_ASAP7_75t_R FILLER_340_232 ();
 FILLER_ASAP7_75t_R FILLER_340_244 ();
 DECAPx1_ASAP7_75t_R FILLER_340_252 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_256 ();
 DECAPx2_ASAP7_75t_R FILLER_340_268 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_274 ();
 DECAPx2_ASAP7_75t_R FILLER_340_283 ();
 DECAPx2_ASAP7_75t_R FILLER_340_297 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_303 ();
 FILLER_ASAP7_75t_R FILLER_340_310 ();
 DECAPx2_ASAP7_75t_R FILLER_340_318 ();
 FILLER_ASAP7_75t_R FILLER_340_324 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_362 ();
 DECAPx10_ASAP7_75t_R FILLER_340_389 ();
 DECAPx10_ASAP7_75t_R FILLER_340_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_433 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_476 ();
 DECAPx1_ASAP7_75t_R FILLER_340_484 ();
 DECAPx2_ASAP7_75t_R FILLER_340_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_509 ();
 DECAPx1_ASAP7_75t_R FILLER_340_513 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_517 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_544 ();
 DECAPx1_ASAP7_75t_R FILLER_340_564 ();
 DECAPx6_ASAP7_75t_R FILLER_340_571 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_585 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_591 ();
 DECAPx2_ASAP7_75t_R FILLER_340_597 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_620 ();
 DECAPx2_ASAP7_75t_R FILLER_340_668 ();
 DECAPx10_ASAP7_75t_R FILLER_340_677 ();
 DECAPx10_ASAP7_75t_R FILLER_340_699 ();
 DECAPx10_ASAP7_75t_R FILLER_340_721 ();
 DECAPx10_ASAP7_75t_R FILLER_340_743 ();
 DECAPx4_ASAP7_75t_R FILLER_340_765 ();
 DECAPx1_ASAP7_75t_R FILLER_340_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_340_785 ();
 DECAPx6_ASAP7_75t_R FILLER_340_794 ();
 FILLER_ASAP7_75t_R FILLER_340_823 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_340_837 ();
 DECAPx4_ASAP7_75t_R FILLER_340_869 ();
 FILLER_ASAP7_75t_R FILLER_340_895 ();
 DECAPx10_ASAP7_75t_R FILLER_340_900 ();
 DECAPx4_ASAP7_75t_R FILLER_340_922 ();
 FILLER_ASAP7_75t_R FILLER_340_932 ();
 DECAPx10_ASAP7_75t_R FILLER_341_2 ();
 DECAPx10_ASAP7_75t_R FILLER_341_24 ();
 DECAPx10_ASAP7_75t_R FILLER_341_46 ();
 DECAPx10_ASAP7_75t_R FILLER_341_68 ();
 DECAPx10_ASAP7_75t_R FILLER_341_90 ();
 DECAPx2_ASAP7_75t_R FILLER_341_112 ();
 FILLER_ASAP7_75t_R FILLER_341_118 ();
 DECAPx4_ASAP7_75t_R FILLER_341_126 ();
 DECAPx6_ASAP7_75t_R FILLER_341_142 ();
 DECAPx1_ASAP7_75t_R FILLER_341_156 ();
 FILLER_ASAP7_75t_R FILLER_341_166 ();
 DECAPx4_ASAP7_75t_R FILLER_341_174 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_184 ();
 DECAPx1_ASAP7_75t_R FILLER_341_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_217 ();
 DECAPx4_ASAP7_75t_R FILLER_341_224 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_234 ();
 DECAPx10_ASAP7_75t_R FILLER_341_247 ();
 DECAPx6_ASAP7_75t_R FILLER_341_269 ();
 DECAPx1_ASAP7_75t_R FILLER_341_295 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_328 ();
 DECAPx6_ASAP7_75t_R FILLER_341_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_366 ();
 DECAPx1_ASAP7_75t_R FILLER_341_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_377 ();
 DECAPx10_ASAP7_75t_R FILLER_341_381 ();
 DECAPx1_ASAP7_75t_R FILLER_341_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_407 ();
 DECAPx4_ASAP7_75t_R FILLER_341_427 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_437 ();
 DECAPx1_ASAP7_75t_R FILLER_341_448 ();
 DECAPx6_ASAP7_75t_R FILLER_341_494 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_508 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_531 ();
 DECAPx10_ASAP7_75t_R FILLER_341_574 ();
 DECAPx4_ASAP7_75t_R FILLER_341_596 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_606 ();
 DECAPx2_ASAP7_75t_R FILLER_341_622 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_628 ();
 DECAPx1_ASAP7_75t_R FILLER_341_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_645 ();
 FILLER_ASAP7_75t_R FILLER_341_663 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_671 ();
 DECAPx4_ASAP7_75t_R FILLER_341_677 ();
 FILLER_ASAP7_75t_R FILLER_341_687 ();
 DECAPx10_ASAP7_75t_R FILLER_341_695 ();
 DECAPx10_ASAP7_75t_R FILLER_341_717 ();
 DECAPx6_ASAP7_75t_R FILLER_341_739 ();
 DECAPx1_ASAP7_75t_R FILLER_341_753 ();
 DECAPx2_ASAP7_75t_R FILLER_341_773 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_779 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_803 ();
 DECAPx2_ASAP7_75t_R FILLER_341_810 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_816 ();
 DECAPx10_ASAP7_75t_R FILLER_341_825 ();
 DECAPx2_ASAP7_75t_R FILLER_341_847 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_853 ();
 DECAPx2_ASAP7_75t_R FILLER_341_857 ();
 FILLER_ASAP7_75t_R FILLER_341_880 ();
 DECAPx6_ASAP7_75t_R FILLER_341_908 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_341_922 ();
 DECAPx2_ASAP7_75t_R FILLER_341_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_341_933 ();
 DECAPx10_ASAP7_75t_R FILLER_342_2 ();
 DECAPx10_ASAP7_75t_R FILLER_342_24 ();
 DECAPx10_ASAP7_75t_R FILLER_342_46 ();
 DECAPx10_ASAP7_75t_R FILLER_342_68 ();
 DECAPx10_ASAP7_75t_R FILLER_342_90 ();
 DECAPx2_ASAP7_75t_R FILLER_342_112 ();
 FILLER_ASAP7_75t_R FILLER_342_118 ();
 DECAPx2_ASAP7_75t_R FILLER_342_133 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_139 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_154 ();
 DECAPx6_ASAP7_75t_R FILLER_342_181 ();
 DECAPx2_ASAP7_75t_R FILLER_342_195 ();
 DECAPx1_ASAP7_75t_R FILLER_342_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_208 ();
 DECAPx10_ASAP7_75t_R FILLER_342_215 ();
 DECAPx6_ASAP7_75t_R FILLER_342_237 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_342_251 ();
 DECAPx10_ASAP7_75t_R FILLER_342_260 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_282 ();
 DECAPx6_ASAP7_75t_R FILLER_342_291 ();
 FILLER_ASAP7_75t_R FILLER_342_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_313 ();
 DECAPx4_ASAP7_75t_R FILLER_342_317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_342_327 ();
 DECAPx10_ASAP7_75t_R FILLER_342_338 ();
 DECAPx10_ASAP7_75t_R FILLER_342_360 ();
 DECAPx6_ASAP7_75t_R FILLER_342_382 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_416 ();
 FILLER_ASAP7_75t_R FILLER_342_430 ();
 DECAPx2_ASAP7_75t_R FILLER_342_445 ();
 FILLER_ASAP7_75t_R FILLER_342_451 ();
 DECAPx1_ASAP7_75t_R FILLER_342_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_474 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_342_486 ();
 DECAPx6_ASAP7_75t_R FILLER_342_497 ();
 DECAPx2_ASAP7_75t_R FILLER_342_511 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_517 ();
 FILLER_ASAP7_75t_R FILLER_342_530 ();
 DECAPx2_ASAP7_75t_R FILLER_342_546 ();
 DECAPx2_ASAP7_75t_R FILLER_342_566 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_342_572 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_578 ();
 DECAPx4_ASAP7_75t_R FILLER_342_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_603 ();
 DECAPx6_ASAP7_75t_R FILLER_342_630 ();
 DECAPx1_ASAP7_75t_R FILLER_342_644 ();
 DECAPx10_ASAP7_75t_R FILLER_342_690 ();
 DECAPx10_ASAP7_75t_R FILLER_342_712 ();
 DECAPx6_ASAP7_75t_R FILLER_342_734 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_342_748 ();
 DECAPx1_ASAP7_75t_R FILLER_342_777 ();
 DECAPx2_ASAP7_75t_R FILLER_342_807 ();
 DECAPx6_ASAP7_75t_R FILLER_342_816 ();
 FILLER_ASAP7_75t_R FILLER_342_830 ();
 DECAPx10_ASAP7_75t_R FILLER_342_838 ();
 DECAPx2_ASAP7_75t_R FILLER_342_860 ();
 FILLERxp5_ASAP7_75t_R FILLER_342_866 ();
 DECAPx10_ASAP7_75t_R FILLER_342_870 ();
 DECAPx10_ASAP7_75t_R FILLER_342_892 ();
 DECAPx6_ASAP7_75t_R FILLER_342_914 ();
 DECAPx2_ASAP7_75t_R FILLER_342_928 ();
 DECAPx10_ASAP7_75t_R FILLER_343_2 ();
 DECAPx10_ASAP7_75t_R FILLER_343_24 ();
 DECAPx10_ASAP7_75t_R FILLER_343_46 ();
 DECAPx10_ASAP7_75t_R FILLER_343_68 ();
 DECAPx4_ASAP7_75t_R FILLER_343_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_100 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_134 ();
 DECAPx6_ASAP7_75t_R FILLER_343_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_187 ();
 DECAPx10_ASAP7_75t_R FILLER_343_196 ();
 DECAPx1_ASAP7_75t_R FILLER_343_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_222 ();
 DECAPx4_ASAP7_75t_R FILLER_343_229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_239 ();
 DECAPx1_ASAP7_75t_R FILLER_343_254 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_258 ();
 DECAPx1_ASAP7_75t_R FILLER_343_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_275 ();
 DECAPx6_ASAP7_75t_R FILLER_343_284 ();
 DECAPx1_ASAP7_75t_R FILLER_343_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_331 ();
 DECAPx10_ASAP7_75t_R FILLER_343_340 ();
 DECAPx4_ASAP7_75t_R FILLER_343_362 ();
 FILLER_ASAP7_75t_R FILLER_343_372 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_383 ();
 DECAPx6_ASAP7_75t_R FILLER_343_397 ();
 DECAPx1_ASAP7_75t_R FILLER_343_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_446 ();
 DECAPx2_ASAP7_75t_R FILLER_343_462 ();
 FILLER_ASAP7_75t_R FILLER_343_468 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_475 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_482 ();
 DECAPx10_ASAP7_75t_R FILLER_343_488 ();
 DECAPx10_ASAP7_75t_R FILLER_343_510 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_532 ();
 DECAPx6_ASAP7_75t_R FILLER_343_538 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_552 ();
 DECAPx10_ASAP7_75t_R FILLER_343_558 ();
 DECAPx1_ASAP7_75t_R FILLER_343_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_584 ();
 DECAPx10_ASAP7_75t_R FILLER_343_619 ();
 DECAPx6_ASAP7_75t_R FILLER_343_641 ();
 DECAPx2_ASAP7_75t_R FILLER_343_655 ();
 DECAPx4_ASAP7_75t_R FILLER_343_667 ();
 DECAPx10_ASAP7_75t_R FILLER_343_697 ();
 DECAPx10_ASAP7_75t_R FILLER_343_719 ();
 DECAPx6_ASAP7_75t_R FILLER_343_741 ();
 DECAPx1_ASAP7_75t_R FILLER_343_755 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_774 ();
 DECAPx6_ASAP7_75t_R FILLER_343_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_795 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_799 ();
 DECAPx2_ASAP7_75t_R FILLER_343_819 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_343_825 ();
 DECAPx1_ASAP7_75t_R FILLER_343_850 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_854 ();
 DECAPx10_ASAP7_75t_R FILLER_343_885 ();
 DECAPx6_ASAP7_75t_R FILLER_343_907 ();
 DECAPx1_ASAP7_75t_R FILLER_343_921 ();
 DECAPx2_ASAP7_75t_R FILLER_343_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_343_933 ();
 DECAPx10_ASAP7_75t_R FILLER_344_2 ();
 DECAPx10_ASAP7_75t_R FILLER_344_24 ();
 DECAPx10_ASAP7_75t_R FILLER_344_46 ();
 DECAPx6_ASAP7_75t_R FILLER_344_68 ();
 DECAPx1_ASAP7_75t_R FILLER_344_82 ();
 DECAPx1_ASAP7_75t_R FILLER_344_120 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_124 ();
 DECAPx1_ASAP7_75t_R FILLER_344_147 ();
 DECAPx6_ASAP7_75t_R FILLER_344_166 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_180 ();
 DECAPx6_ASAP7_75t_R FILLER_344_218 ();
 DECAPx2_ASAP7_75t_R FILLER_344_232 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_238 ();
 DECAPx10_ASAP7_75t_R FILLER_344_277 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_299 ();
 DECAPx1_ASAP7_75t_R FILLER_344_308 ();
 DECAPx6_ASAP7_75t_R FILLER_344_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_329 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_342 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_397 ();
 DECAPx1_ASAP7_75t_R FILLER_344_406 ();
 DECAPx2_ASAP7_75t_R FILLER_344_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_451 ();
 DECAPx6_ASAP7_75t_R FILLER_344_464 ();
 DECAPx2_ASAP7_75t_R FILLER_344_478 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_484 ();
 DECAPx1_ASAP7_75t_R FILLER_344_490 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_502 ();
 DECAPx2_ASAP7_75t_R FILLER_344_513 ();
 FILLER_ASAP7_75t_R FILLER_344_519 ();
 DECAPx10_ASAP7_75t_R FILLER_344_526 ();
 DECAPx10_ASAP7_75t_R FILLER_344_548 ();
 DECAPx1_ASAP7_75t_R FILLER_344_570 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_577 ();
 DECAPx4_ASAP7_75t_R FILLER_344_583 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_613 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_624 ();
 FILLER_ASAP7_75t_R FILLER_344_633 ();
 DECAPx2_ASAP7_75t_R FILLER_344_649 ();
 FILLER_ASAP7_75t_R FILLER_344_655 ();
 DECAPx10_ASAP7_75t_R FILLER_344_662 ();
 DECAPx10_ASAP7_75t_R FILLER_344_684 ();
 DECAPx10_ASAP7_75t_R FILLER_344_706 ();
 DECAPx10_ASAP7_75t_R FILLER_344_728 ();
 DECAPx6_ASAP7_75t_R FILLER_344_750 ();
 FILLER_ASAP7_75t_R FILLER_344_764 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_769 ();
 DECAPx10_ASAP7_75t_R FILLER_344_778 ();
 DECAPx4_ASAP7_75t_R FILLER_344_800 ();
 FILLER_ASAP7_75t_R FILLER_344_810 ();
 DECAPx1_ASAP7_75t_R FILLER_344_815 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_819 ();
 DECAPx2_ASAP7_75t_R FILLER_344_858 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_344_864 ();
 DECAPx10_ASAP7_75t_R FILLER_344_893 ();
 DECAPx6_ASAP7_75t_R FILLER_344_915 ();
 DECAPx1_ASAP7_75t_R FILLER_344_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_344_933 ();
 DECAPx10_ASAP7_75t_R FILLER_345_2 ();
 DECAPx10_ASAP7_75t_R FILLER_345_24 ();
 DECAPx10_ASAP7_75t_R FILLER_345_46 ();
 DECAPx10_ASAP7_75t_R FILLER_345_68 ();
 DECAPx2_ASAP7_75t_R FILLER_345_90 ();
 FILLER_ASAP7_75t_R FILLER_345_96 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_107 ();
 DECAPx10_ASAP7_75t_R FILLER_345_140 ();
 DECAPx10_ASAP7_75t_R FILLER_345_162 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_184 ();
 DECAPx1_ASAP7_75t_R FILLER_345_191 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_195 ();
 DECAPx4_ASAP7_75t_R FILLER_345_199 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_345_209 ();
 DECAPx1_ASAP7_75t_R FILLER_345_220 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_224 ();
 DECAPx2_ASAP7_75t_R FILLER_345_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_271 ();
 DECAPx2_ASAP7_75t_R FILLER_345_278 ();
 FILLER_ASAP7_75t_R FILLER_345_284 ();
 DECAPx10_ASAP7_75t_R FILLER_345_289 ();
 DECAPx1_ASAP7_75t_R FILLER_345_311 ();
 DECAPx2_ASAP7_75t_R FILLER_345_327 ();
 FILLER_ASAP7_75t_R FILLER_345_368 ();
 DECAPx4_ASAP7_75t_R FILLER_345_376 ();
 FILLER_ASAP7_75t_R FILLER_345_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_420 ();
 DECAPx2_ASAP7_75t_R FILLER_345_436 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_453 ();
 FILLER_ASAP7_75t_R FILLER_345_468 ();
 DECAPx2_ASAP7_75t_R FILLER_345_476 ();
 DECAPx1_ASAP7_75t_R FILLER_345_501 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_345_515 ();
 DECAPx10_ASAP7_75t_R FILLER_345_521 ();
 DECAPx2_ASAP7_75t_R FILLER_345_543 ();
 DECAPx2_ASAP7_75t_R FILLER_345_552 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_345_558 ();
 DECAPx2_ASAP7_75t_R FILLER_345_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_587 ();
 DECAPx4_ASAP7_75t_R FILLER_345_597 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_607 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_611 ();
 DECAPx4_ASAP7_75t_R FILLER_345_638 ();
 FILLER_ASAP7_75t_R FILLER_345_648 ();
 DECAPx10_ASAP7_75t_R FILLER_345_662 ();
 DECAPx10_ASAP7_75t_R FILLER_345_684 ();
 DECAPx10_ASAP7_75t_R FILLER_345_706 ();
 DECAPx10_ASAP7_75t_R FILLER_345_728 ();
 DECAPx6_ASAP7_75t_R FILLER_345_750 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_764 ();
 DECAPx4_ASAP7_75t_R FILLER_345_781 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_791 ();
 DECAPx2_ASAP7_75t_R FILLER_345_810 ();
 FILLER_ASAP7_75t_R FILLER_345_816 ();
 DECAPx10_ASAP7_75t_R FILLER_345_824 ();
 DECAPx10_ASAP7_75t_R FILLER_345_849 ();
 DECAPx4_ASAP7_75t_R FILLER_345_871 ();
 DECAPx10_ASAP7_75t_R FILLER_345_884 ();
 DECAPx6_ASAP7_75t_R FILLER_345_906 ();
 DECAPx1_ASAP7_75t_R FILLER_345_920 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_924 ();
 DECAPx2_ASAP7_75t_R FILLER_345_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_345_933 ();
 DECAPx10_ASAP7_75t_R FILLER_346_2 ();
 DECAPx10_ASAP7_75t_R FILLER_346_24 ();
 DECAPx10_ASAP7_75t_R FILLER_346_46 ();
 DECAPx10_ASAP7_75t_R FILLER_346_68 ();
 DECAPx10_ASAP7_75t_R FILLER_346_90 ();
 DECAPx4_ASAP7_75t_R FILLER_346_112 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_122 ();
 DECAPx10_ASAP7_75t_R FILLER_346_129 ();
 DECAPx6_ASAP7_75t_R FILLER_346_151 ();
 DECAPx2_ASAP7_75t_R FILLER_346_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_171 ();
 DECAPx6_ASAP7_75t_R FILLER_346_178 ();
 DECAPx1_ASAP7_75t_R FILLER_346_204 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_208 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_221 ();
 DECAPx2_ASAP7_75t_R FILLER_346_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_250 ();
 DECAPx1_ASAP7_75t_R FILLER_346_256 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_263 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_292 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_299 ();
 DECAPx1_ASAP7_75t_R FILLER_346_306 ();
 DECAPx2_ASAP7_75t_R FILLER_346_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_342 ();
 DECAPx4_ASAP7_75t_R FILLER_346_364 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_374 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_383 ();
 DECAPx1_ASAP7_75t_R FILLER_346_392 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_396 ();
 DECAPx1_ASAP7_75t_R FILLER_346_403 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_407 ();
 DECAPx2_ASAP7_75t_R FILLER_346_411 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_417 ();
 DECAPx10_ASAP7_75t_R FILLER_346_426 ();
 DECAPx1_ASAP7_75t_R FILLER_346_448 ();
 FILLER_ASAP7_75t_R FILLER_346_460 ();
 DECAPx6_ASAP7_75t_R FILLER_346_483 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_497 ();
 FILLER_ASAP7_75t_R FILLER_346_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_528 ();
 DECAPx2_ASAP7_75t_R FILLER_346_554 ();
 FILLER_ASAP7_75t_R FILLER_346_560 ();
 DECAPx1_ASAP7_75t_R FILLER_346_565 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_586 ();
 DECAPx4_ASAP7_75t_R FILLER_346_606 ();
 DECAPx1_ASAP7_75t_R FILLER_346_678 ();
 DECAPx10_ASAP7_75t_R FILLER_346_685 ();
 DECAPx10_ASAP7_75t_R FILLER_346_707 ();
 DECAPx10_ASAP7_75t_R FILLER_346_729 ();
 DECAPx6_ASAP7_75t_R FILLER_346_751 ();
 FILLERxp5_ASAP7_75t_R FILLER_346_791 ();
 FILLER_ASAP7_75t_R FILLER_346_805 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_346_815 ();
 DECAPx10_ASAP7_75t_R FILLER_346_828 ();
 DECAPx10_ASAP7_75t_R FILLER_346_850 ();
 DECAPx10_ASAP7_75t_R FILLER_346_872 ();
 DECAPx10_ASAP7_75t_R FILLER_346_894 ();
 DECAPx6_ASAP7_75t_R FILLER_346_916 ();
 DECAPx1_ASAP7_75t_R FILLER_346_930 ();
 DECAPx10_ASAP7_75t_R FILLER_347_2 ();
 DECAPx10_ASAP7_75t_R FILLER_347_24 ();
 DECAPx10_ASAP7_75t_R FILLER_347_46 ();
 DECAPx10_ASAP7_75t_R FILLER_347_68 ();
 DECAPx10_ASAP7_75t_R FILLER_347_90 ();
 DECAPx2_ASAP7_75t_R FILLER_347_112 ();
 FILLER_ASAP7_75t_R FILLER_347_118 ();
 DECAPx6_ASAP7_75t_R FILLER_347_126 ();
 DECAPx2_ASAP7_75t_R FILLER_347_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_146 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_347_167 ();
 DECAPx4_ASAP7_75t_R FILLER_347_176 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_186 ();
 DECAPx4_ASAP7_75t_R FILLER_347_213 ();
 DECAPx10_ASAP7_75t_R FILLER_347_229 ();
 DECAPx6_ASAP7_75t_R FILLER_347_251 ();
 DECAPx1_ASAP7_75t_R FILLER_347_265 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_309 ();
 DECAPx2_ASAP7_75t_R FILLER_347_316 ();
 FILLER_ASAP7_75t_R FILLER_347_322 ();
 DECAPx10_ASAP7_75t_R FILLER_347_327 ();
 DECAPx6_ASAP7_75t_R FILLER_347_349 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_347_363 ();
 DECAPx4_ASAP7_75t_R FILLER_347_392 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_347_402 ();
 DECAPx4_ASAP7_75t_R FILLER_347_411 ();
 FILLER_ASAP7_75t_R FILLER_347_421 ();
 DECAPx6_ASAP7_75t_R FILLER_347_428 ();
 DECAPx1_ASAP7_75t_R FILLER_347_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_446 ();
 DECAPx1_ASAP7_75t_R FILLER_347_452 ();
 DECAPx4_ASAP7_75t_R FILLER_347_461 ();
 DECAPx6_ASAP7_75t_R FILLER_347_489 ();
 FILLER_ASAP7_75t_R FILLER_347_509 ();
 FILLER_ASAP7_75t_R FILLER_347_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_560 ();
 DECAPx4_ASAP7_75t_R FILLER_347_575 ();
 FILLER_ASAP7_75t_R FILLER_347_585 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_590 ();
 DECAPx10_ASAP7_75t_R FILLER_347_608 ();
 DECAPx4_ASAP7_75t_R FILLER_347_630 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_347_640 ();
 DECAPx4_ASAP7_75t_R FILLER_347_652 ();
 FILLER_ASAP7_75t_R FILLER_347_679 ();
 DECAPx10_ASAP7_75t_R FILLER_347_687 ();
 DECAPx10_ASAP7_75t_R FILLER_347_709 ();
 DECAPx10_ASAP7_75t_R FILLER_347_731 ();
 DECAPx10_ASAP7_75t_R FILLER_347_753 ();
 DECAPx1_ASAP7_75t_R FILLER_347_775 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_347_782 ();
 DECAPx10_ASAP7_75t_R FILLER_347_837 ();
 DECAPx10_ASAP7_75t_R FILLER_347_859 ();
 DECAPx10_ASAP7_75t_R FILLER_347_881 ();
 DECAPx10_ASAP7_75t_R FILLER_347_903 ();
 DECAPx2_ASAP7_75t_R FILLER_347_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_347_933 ();
 DECAPx10_ASAP7_75t_R FILLER_348_2 ();
 DECAPx10_ASAP7_75t_R FILLER_348_24 ();
 DECAPx10_ASAP7_75t_R FILLER_348_46 ();
 DECAPx10_ASAP7_75t_R FILLER_348_68 ();
 DECAPx2_ASAP7_75t_R FILLER_348_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_96 ();
 DECAPx2_ASAP7_75t_R FILLER_348_111 ();
 FILLER_ASAP7_75t_R FILLER_348_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_125 ();
 DECAPx1_ASAP7_75t_R FILLER_348_132 ();
 DECAPx1_ASAP7_75t_R FILLER_348_176 ();
 DECAPx4_ASAP7_75t_R FILLER_348_192 ();
 DECAPx2_ASAP7_75t_R FILLER_348_205 ();
 FILLER_ASAP7_75t_R FILLER_348_211 ();
 DECAPx10_ASAP7_75t_R FILLER_348_239 ();
 DECAPx6_ASAP7_75t_R FILLER_348_261 ();
 FILLER_ASAP7_75t_R FILLER_348_275 ();
 DECAPx10_ASAP7_75t_R FILLER_348_295 ();
 DECAPx10_ASAP7_75t_R FILLER_348_317 ();
 DECAPx6_ASAP7_75t_R FILLER_348_339 ();
 FILLER_ASAP7_75t_R FILLER_348_359 ();
 DECAPx2_ASAP7_75t_R FILLER_348_364 ();
 FILLER_ASAP7_75t_R FILLER_348_370 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_378 ();
 DECAPx2_ASAP7_75t_R FILLER_348_384 ();
 FILLER_ASAP7_75t_R FILLER_348_390 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_418 ();
 DECAPx2_ASAP7_75t_R FILLER_348_428 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_434 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_440 ();
 DECAPx2_ASAP7_75t_R FILLER_348_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_456 ();
 DECAPx1_ASAP7_75t_R FILLER_348_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_468 ();
 DECAPx2_ASAP7_75t_R FILLER_348_495 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_501 ();
 DECAPx2_ASAP7_75t_R FILLER_348_509 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_515 ();
 FILLERxp5_ASAP7_75t_R FILLER_348_519 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_534 ();
 DECAPx10_ASAP7_75t_R FILLER_348_551 ();
 DECAPx10_ASAP7_75t_R FILLER_348_573 ();
 DECAPx4_ASAP7_75t_R FILLER_348_595 ();
 FILLER_ASAP7_75t_R FILLER_348_605 ();
 DECAPx10_ASAP7_75t_R FILLER_348_613 ();
 DECAPx2_ASAP7_75t_R FILLER_348_635 ();
 DECAPx6_ASAP7_75t_R FILLER_348_655 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_669 ();
 DECAPx10_ASAP7_75t_R FILLER_348_695 ();
 DECAPx10_ASAP7_75t_R FILLER_348_717 ();
 DECAPx10_ASAP7_75t_R FILLER_348_739 ();
 DECAPx10_ASAP7_75t_R FILLER_348_761 ();
 DECAPx6_ASAP7_75t_R FILLER_348_783 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_348_797 ();
 DECAPx10_ASAP7_75t_R FILLER_348_826 ();
 DECAPx10_ASAP7_75t_R FILLER_348_848 ();
 DECAPx10_ASAP7_75t_R FILLER_348_870 ();
 DECAPx10_ASAP7_75t_R FILLER_348_892 ();
 DECAPx6_ASAP7_75t_R FILLER_348_914 ();
 DECAPx2_ASAP7_75t_R FILLER_348_928 ();
 DECAPx10_ASAP7_75t_R FILLER_349_2 ();
 DECAPx10_ASAP7_75t_R FILLER_349_24 ();
 DECAPx10_ASAP7_75t_R FILLER_349_46 ();
 DECAPx10_ASAP7_75t_R FILLER_349_68 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_90 ();
 FILLER_ASAP7_75t_R FILLER_349_149 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_154 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_161 ();
 DECAPx10_ASAP7_75t_R FILLER_349_196 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_349_224 ();
 DECAPx2_ASAP7_75t_R FILLER_349_230 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_236 ();
 DECAPx10_ASAP7_75t_R FILLER_349_263 ();
 DECAPx4_ASAP7_75t_R FILLER_349_285 ();
 FILLER_ASAP7_75t_R FILLER_349_295 ();
 DECAPx2_ASAP7_75t_R FILLER_349_303 ();
 FILLER_ASAP7_75t_R FILLER_349_309 ();
 DECAPx2_ASAP7_75t_R FILLER_349_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_346 ();
 DECAPx10_ASAP7_75t_R FILLER_349_373 ();
 DECAPx1_ASAP7_75t_R FILLER_349_427 ();
 DECAPx1_ASAP7_75t_R FILLER_349_452 ();
 DECAPx6_ASAP7_75t_R FILLER_349_463 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_349_477 ();
 DECAPx6_ASAP7_75t_R FILLER_349_491 ();
 DECAPx2_ASAP7_75t_R FILLER_349_505 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_511 ();
 DECAPx10_ASAP7_75t_R FILLER_349_553 ();
 DECAPx6_ASAP7_75t_R FILLER_349_575 ();
 DECAPx2_ASAP7_75t_R FILLER_349_589 ();
 DECAPx2_ASAP7_75t_R FILLER_349_598 ();
 DECAPx2_ASAP7_75t_R FILLER_349_624 ();
 FILLER_ASAP7_75t_R FILLER_349_630 ();
 DECAPx10_ASAP7_75t_R FILLER_349_635 ();
 FILLER_ASAP7_75t_R FILLER_349_657 ();
 DECAPx1_ASAP7_75t_R FILLER_349_662 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_666 ();
 DECAPx2_ASAP7_75t_R FILLER_349_670 ();
 DECAPx10_ASAP7_75t_R FILLER_349_682 ();
 DECAPx10_ASAP7_75t_R FILLER_349_704 ();
 DECAPx10_ASAP7_75t_R FILLER_349_726 ();
 DECAPx10_ASAP7_75t_R FILLER_349_748 ();
 DECAPx10_ASAP7_75t_R FILLER_349_770 ();
 DECAPx10_ASAP7_75t_R FILLER_349_792 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_814 ();
 DECAPx2_ASAP7_75t_R FILLER_349_818 ();
 FILLER_ASAP7_75t_R FILLER_349_824 ();
 DECAPx10_ASAP7_75t_R FILLER_349_829 ();
 DECAPx10_ASAP7_75t_R FILLER_349_851 ();
 DECAPx10_ASAP7_75t_R FILLER_349_873 ();
 DECAPx10_ASAP7_75t_R FILLER_349_895 ();
 DECAPx2_ASAP7_75t_R FILLER_349_917 ();
 FILLER_ASAP7_75t_R FILLER_349_923 ();
 DECAPx2_ASAP7_75t_R FILLER_349_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_349_933 ();
 DECAPx10_ASAP7_75t_R FILLER_350_2 ();
 DECAPx10_ASAP7_75t_R FILLER_350_24 ();
 DECAPx10_ASAP7_75t_R FILLER_350_46 ();
 DECAPx10_ASAP7_75t_R FILLER_350_68 ();
 DECAPx6_ASAP7_75t_R FILLER_350_90 ();
 FILLER_ASAP7_75t_R FILLER_350_104 ();
 DECAPx1_ASAP7_75t_R FILLER_350_109 ();
 DECAPx10_ASAP7_75t_R FILLER_350_142 ();
 DECAPx2_ASAP7_75t_R FILLER_350_164 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_184 ();
 DECAPx10_ASAP7_75t_R FILLER_350_188 ();
 DECAPx10_ASAP7_75t_R FILLER_350_210 ();
 DECAPx4_ASAP7_75t_R FILLER_350_232 ();
 DECAPx6_ASAP7_75t_R FILLER_350_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_280 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_290 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_296 ();
 DECAPx4_ASAP7_75t_R FILLER_350_305 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_315 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_330 ();
 DECAPx1_ASAP7_75t_R FILLER_350_345 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_349 ();
 DECAPx4_ASAP7_75t_R FILLER_350_356 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_366 ();
 DECAPx10_ASAP7_75t_R FILLER_350_376 ();
 DECAPx2_ASAP7_75t_R FILLER_350_398 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_427 ();
 FILLER_ASAP7_75t_R FILLER_350_436 ();
 DECAPx1_ASAP7_75t_R FILLER_350_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_477 ();
 DECAPx1_ASAP7_75t_R FILLER_350_486 ();
 DECAPx10_ASAP7_75t_R FILLER_350_498 ();
 DECAPx1_ASAP7_75t_R FILLER_350_520 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_524 ();
 FILLER_ASAP7_75t_R FILLER_350_534 ();
 DECAPx4_ASAP7_75t_R FILLER_350_545 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_555 ();
 DECAPx1_ASAP7_75t_R FILLER_350_567 ();
 DECAPx1_ASAP7_75t_R FILLER_350_585 ();
 DECAPx6_ASAP7_75t_R FILLER_350_592 ();
 FILLER_ASAP7_75t_R FILLER_350_606 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_350_618 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_624 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_628 ();
 DECAPx4_ASAP7_75t_R FILLER_350_643 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_653 ();
 DECAPx10_ASAP7_75t_R FILLER_350_671 ();
 DECAPx10_ASAP7_75t_R FILLER_350_693 ();
 DECAPx10_ASAP7_75t_R FILLER_350_715 ();
 DECAPx10_ASAP7_75t_R FILLER_350_737 ();
 DECAPx10_ASAP7_75t_R FILLER_350_759 ();
 DECAPx10_ASAP7_75t_R FILLER_350_781 ();
 DECAPx10_ASAP7_75t_R FILLER_350_803 ();
 DECAPx10_ASAP7_75t_R FILLER_350_825 ();
 DECAPx10_ASAP7_75t_R FILLER_350_847 ();
 DECAPx10_ASAP7_75t_R FILLER_350_869 ();
 DECAPx10_ASAP7_75t_R FILLER_350_891 ();
 DECAPx6_ASAP7_75t_R FILLER_350_913 ();
 DECAPx2_ASAP7_75t_R FILLER_350_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_350_933 ();
 DECAPx10_ASAP7_75t_R FILLER_351_2 ();
 DECAPx10_ASAP7_75t_R FILLER_351_24 ();
 DECAPx10_ASAP7_75t_R FILLER_351_46 ();
 DECAPx10_ASAP7_75t_R FILLER_351_68 ();
 DECAPx10_ASAP7_75t_R FILLER_351_90 ();
 DECAPx6_ASAP7_75t_R FILLER_351_112 ();
 FILLER_ASAP7_75t_R FILLER_351_126 ();
 DECAPx10_ASAP7_75t_R FILLER_351_134 ();
 DECAPx10_ASAP7_75t_R FILLER_351_156 ();
 DECAPx10_ASAP7_75t_R FILLER_351_178 ();
 DECAPx2_ASAP7_75t_R FILLER_351_200 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_206 ();
 DECAPx1_ASAP7_75t_R FILLER_351_213 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_217 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_351_224 ();
 DECAPx6_ASAP7_75t_R FILLER_351_233 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_247 ();
 FILLER_ASAP7_75t_R FILLER_351_256 ();
 DECAPx2_ASAP7_75t_R FILLER_351_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_272 ();
 DECAPx1_ASAP7_75t_R FILLER_351_299 ();
 DECAPx2_ASAP7_75t_R FILLER_351_311 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_351_317 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_337 ();
 DECAPx2_ASAP7_75t_R FILLER_351_352 ();
 DECAPx10_ASAP7_75t_R FILLER_351_387 ();
 DECAPx1_ASAP7_75t_R FILLER_351_424 ();
 DECAPx6_ASAP7_75t_R FILLER_351_436 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_351_450 ();
 DECAPx2_ASAP7_75t_R FILLER_351_458 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_351_464 ();
 DECAPx1_ASAP7_75t_R FILLER_351_473 ();
 FILLER_ASAP7_75t_R FILLER_351_483 ();
 DECAPx6_ASAP7_75t_R FILLER_351_513 ();
 DECAPx1_ASAP7_75t_R FILLER_351_527 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_531 ();
 DECAPx2_ASAP7_75t_R FILLER_351_535 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_541 ();
 DECAPx4_ASAP7_75t_R FILLER_351_593 ();
 FILLER_ASAP7_75t_R FILLER_351_603 ();
 DECAPx2_ASAP7_75t_R FILLER_351_608 ();
 DECAPx1_ASAP7_75t_R FILLER_351_645 ();
 DECAPx10_ASAP7_75t_R FILLER_351_652 ();
 DECAPx10_ASAP7_75t_R FILLER_351_674 ();
 DECAPx10_ASAP7_75t_R FILLER_351_696 ();
 DECAPx10_ASAP7_75t_R FILLER_351_718 ();
 DECAPx10_ASAP7_75t_R FILLER_351_740 ();
 DECAPx10_ASAP7_75t_R FILLER_351_762 ();
 DECAPx10_ASAP7_75t_R FILLER_351_784 ();
 DECAPx10_ASAP7_75t_R FILLER_351_806 ();
 DECAPx10_ASAP7_75t_R FILLER_351_828 ();
 DECAPx10_ASAP7_75t_R FILLER_351_850 ();
 DECAPx10_ASAP7_75t_R FILLER_351_872 ();
 DECAPx10_ASAP7_75t_R FILLER_351_894 ();
 DECAPx2_ASAP7_75t_R FILLER_351_916 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_351_922 ();
 DECAPx2_ASAP7_75t_R FILLER_351_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_351_933 ();
 DECAPx10_ASAP7_75t_R FILLER_352_2 ();
 DECAPx10_ASAP7_75t_R FILLER_352_24 ();
 DECAPx10_ASAP7_75t_R FILLER_352_46 ();
 DECAPx10_ASAP7_75t_R FILLER_352_68 ();
 DECAPx10_ASAP7_75t_R FILLER_352_90 ();
 DECAPx10_ASAP7_75t_R FILLER_352_112 ();
 FILLER_ASAP7_75t_R FILLER_352_160 ();
 DECAPx10_ASAP7_75t_R FILLER_352_165 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_187 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_352_197 ();
 FILLER_ASAP7_75t_R FILLER_352_211 ();
 DECAPx2_ASAP7_75t_R FILLER_352_239 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_245 ();
 FILLER_ASAP7_75t_R FILLER_352_252 ();
 DECAPx1_ASAP7_75t_R FILLER_352_260 ();
 DECAPx2_ASAP7_75t_R FILLER_352_283 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_289 ();
 DECAPx4_ASAP7_75t_R FILLER_352_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_303 ();
 DECAPx6_ASAP7_75t_R FILLER_352_345 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_352_359 ();
 DECAPx2_ASAP7_75t_R FILLER_352_368 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_374 ();
 FILLER_ASAP7_75t_R FILLER_352_387 ();
 DECAPx10_ASAP7_75t_R FILLER_352_401 ();
 DECAPx10_ASAP7_75t_R FILLER_352_423 ();
 DECAPx1_ASAP7_75t_R FILLER_352_445 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_449 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_453 ();
 DECAPx1_ASAP7_75t_R FILLER_352_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_468 ();
 DECAPx2_ASAP7_75t_R FILLER_352_479 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_485 ();
 DECAPx2_ASAP7_75t_R FILLER_352_491 ();
 FILLER_ASAP7_75t_R FILLER_352_497 ();
 DECAPx10_ASAP7_75t_R FILLER_352_519 ();
 DECAPx4_ASAP7_75t_R FILLER_352_541 ();
 FILLER_ASAP7_75t_R FILLER_352_551 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_352_567 ();
 FILLER_ASAP7_75t_R FILLER_352_573 ();
 FILLER_ASAP7_75t_R FILLER_352_587 ();
 DECAPx10_ASAP7_75t_R FILLER_352_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_352_625 ();
 DECAPx4_ASAP7_75t_R FILLER_352_634 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_352_644 ();
 DECAPx4_ASAP7_75t_R FILLER_352_650 ();
 DECAPx1_ASAP7_75t_R FILLER_352_663 ();
 DECAPx10_ASAP7_75t_R FILLER_352_670 ();
 DECAPx10_ASAP7_75t_R FILLER_352_692 ();
 DECAPx10_ASAP7_75t_R FILLER_352_714 ();
 DECAPx10_ASAP7_75t_R FILLER_352_736 ();
 DECAPx10_ASAP7_75t_R FILLER_352_758 ();
 DECAPx10_ASAP7_75t_R FILLER_352_780 ();
 DECAPx10_ASAP7_75t_R FILLER_352_802 ();
 DECAPx10_ASAP7_75t_R FILLER_352_824 ();
 DECAPx10_ASAP7_75t_R FILLER_352_846 ();
 DECAPx10_ASAP7_75t_R FILLER_352_868 ();
 DECAPx10_ASAP7_75t_R FILLER_352_890 ();
 DECAPx10_ASAP7_75t_R FILLER_352_912 ();
 DECAPx10_ASAP7_75t_R FILLER_353_2 ();
 DECAPx10_ASAP7_75t_R FILLER_353_24 ();
 DECAPx10_ASAP7_75t_R FILLER_353_46 ();
 DECAPx10_ASAP7_75t_R FILLER_353_68 ();
 DECAPx4_ASAP7_75t_R FILLER_353_90 ();
 DECAPx6_ASAP7_75t_R FILLER_353_112 ();
 DECAPx2_ASAP7_75t_R FILLER_353_126 ();
 DECAPx2_ASAP7_75t_R FILLER_353_173 ();
 FILLER_ASAP7_75t_R FILLER_353_213 ();
 DECAPx10_ASAP7_75t_R FILLER_353_242 ();
 DECAPx10_ASAP7_75t_R FILLER_353_264 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_286 ();
 DECAPx4_ASAP7_75t_R FILLER_353_307 ();
 FILLER_ASAP7_75t_R FILLER_353_349 ();
 DECAPx1_ASAP7_75t_R FILLER_353_357 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_387 ();
 DECAPx1_ASAP7_75t_R FILLER_353_396 ();
 DECAPx6_ASAP7_75t_R FILLER_353_408 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_353_422 ();
 DECAPx10_ASAP7_75t_R FILLER_353_436 ();
 DECAPx6_ASAP7_75t_R FILLER_353_458 ();
 DECAPx1_ASAP7_75t_R FILLER_353_472 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_476 ();
 FILLER_ASAP7_75t_R FILLER_353_482 ();
 DECAPx6_ASAP7_75t_R FILLER_353_489 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_353_503 ();
 DECAPx10_ASAP7_75t_R FILLER_353_512 ();
 DECAPx2_ASAP7_75t_R FILLER_353_534 ();
 FILLER_ASAP7_75t_R FILLER_353_540 ();
 DECAPx10_ASAP7_75t_R FILLER_353_545 ();
 DECAPx10_ASAP7_75t_R FILLER_353_567 ();
 DECAPx1_ASAP7_75t_R FILLER_353_589 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_597 ();
 FILLER_ASAP7_75t_R FILLER_353_604 ();
 DECAPx4_ASAP7_75t_R FILLER_353_611 ();
 DECAPx10_ASAP7_75t_R FILLER_353_631 ();
 DECAPx2_ASAP7_75t_R FILLER_353_653 ();
 FILLER_ASAP7_75t_R FILLER_353_659 ();
 DECAPx10_ASAP7_75t_R FILLER_353_687 ();
 DECAPx10_ASAP7_75t_R FILLER_353_709 ();
 DECAPx10_ASAP7_75t_R FILLER_353_731 ();
 DECAPx10_ASAP7_75t_R FILLER_353_753 ();
 DECAPx10_ASAP7_75t_R FILLER_353_775 ();
 DECAPx10_ASAP7_75t_R FILLER_353_797 ();
 DECAPx10_ASAP7_75t_R FILLER_353_819 ();
 DECAPx10_ASAP7_75t_R FILLER_353_841 ();
 DECAPx10_ASAP7_75t_R FILLER_353_863 ();
 DECAPx10_ASAP7_75t_R FILLER_353_885 ();
 DECAPx6_ASAP7_75t_R FILLER_353_907 ();
 DECAPx1_ASAP7_75t_R FILLER_353_921 ();
 DECAPx2_ASAP7_75t_R FILLER_353_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_353_933 ();
 DECAPx10_ASAP7_75t_R FILLER_354_2 ();
 DECAPx10_ASAP7_75t_R FILLER_354_24 ();
 DECAPx10_ASAP7_75t_R FILLER_354_46 ();
 DECAPx10_ASAP7_75t_R FILLER_354_68 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_354_90 ();
 DECAPx1_ASAP7_75t_R FILLER_354_125 ();
 DECAPx2_ASAP7_75t_R FILLER_354_135 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_147 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_157 ();
 DECAPx6_ASAP7_75t_R FILLER_354_161 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_354_175 ();
 DECAPx2_ASAP7_75t_R FILLER_354_190 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_208 ();
 DECAPx2_ASAP7_75t_R FILLER_354_235 ();
 DECAPx6_ASAP7_75t_R FILLER_354_247 ();
 FILLER_ASAP7_75t_R FILLER_354_261 ();
 DECAPx4_ASAP7_75t_R FILLER_354_271 ();
 FILLER_ASAP7_75t_R FILLER_354_281 ();
 DECAPx6_ASAP7_75t_R FILLER_354_289 ();
 DECAPx2_ASAP7_75t_R FILLER_354_303 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_309 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_318 ();
 DECAPx10_ASAP7_75t_R FILLER_354_334 ();
 DECAPx2_ASAP7_75t_R FILLER_354_382 ();
 FILLER_ASAP7_75t_R FILLER_354_388 ();
 DECAPx1_ASAP7_75t_R FILLER_354_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_400 ();
 FILLER_ASAP7_75t_R FILLER_354_407 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_354_423 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_436 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_354_443 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_461 ();
 DECAPx1_ASAP7_75t_R FILLER_354_470 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_474 ();
 DECAPx1_ASAP7_75t_R FILLER_354_486 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_490 ();
 DECAPx6_ASAP7_75t_R FILLER_354_499 ();
 DECAPx2_ASAP7_75t_R FILLER_354_513 ();
 FILLER_ASAP7_75t_R FILLER_354_525 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_553 ();
 DECAPx1_ASAP7_75t_R FILLER_354_557 ();
 DECAPx6_ASAP7_75t_R FILLER_354_564 ();
 DECAPx2_ASAP7_75t_R FILLER_354_578 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_584 ();
 DECAPx6_ASAP7_75t_R FILLER_354_622 ();
 FILLERxp5_ASAP7_75t_R FILLER_354_636 ();
 DECAPx4_ASAP7_75t_R FILLER_354_663 ();
 DECAPx10_ASAP7_75t_R FILLER_354_696 ();
 DECAPx10_ASAP7_75t_R FILLER_354_718 ();
 DECAPx10_ASAP7_75t_R FILLER_354_740 ();
 DECAPx10_ASAP7_75t_R FILLER_354_762 ();
 DECAPx10_ASAP7_75t_R FILLER_354_784 ();
 DECAPx6_ASAP7_75t_R FILLER_354_806 ();
 DECAPx1_ASAP7_75t_R FILLER_354_820 ();
 DECAPx10_ASAP7_75t_R FILLER_354_829 ();
 DECAPx10_ASAP7_75t_R FILLER_354_851 ();
 DECAPx10_ASAP7_75t_R FILLER_354_873 ();
 DECAPx10_ASAP7_75t_R FILLER_354_895 ();
 DECAPx6_ASAP7_75t_R FILLER_354_917 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_354_931 ();
 DECAPx10_ASAP7_75t_R FILLER_355_2 ();
 DECAPx10_ASAP7_75t_R FILLER_355_24 ();
 DECAPx10_ASAP7_75t_R FILLER_355_46 ();
 DECAPx10_ASAP7_75t_R FILLER_355_68 ();
 DECAPx6_ASAP7_75t_R FILLER_355_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_355_104 ();
 FILLER_ASAP7_75t_R FILLER_355_110 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_355_124 ();
 DECAPx10_ASAP7_75t_R FILLER_355_133 ();
 DECAPx2_ASAP7_75t_R FILLER_355_155 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_355_161 ();
 DECAPx1_ASAP7_75t_R FILLER_355_170 ();
 DECAPx10_ASAP7_75t_R FILLER_355_200 ();
 DECAPx4_ASAP7_75t_R FILLER_355_222 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_355_258 ();
 DECAPx4_ASAP7_75t_R FILLER_355_301 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_311 ();
 DECAPx10_ASAP7_75t_R FILLER_355_318 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_340 ();
 DECAPx6_ASAP7_75t_R FILLER_355_354 ();
 FILLER_ASAP7_75t_R FILLER_355_368 ();
 DECAPx10_ASAP7_75t_R FILLER_355_373 ();
 DECAPx2_ASAP7_75t_R FILLER_355_395 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_401 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_408 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_451 ();
 DECAPx2_ASAP7_75t_R FILLER_355_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_470 ();
 DECAPx1_ASAP7_75t_R FILLER_355_488 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_492 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_355_501 ();
 DECAPx2_ASAP7_75t_R FILLER_355_545 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_551 ();
 DECAPx10_ASAP7_75t_R FILLER_355_569 ();
 DECAPx2_ASAP7_75t_R FILLER_355_591 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_597 ();
 DECAPx2_ASAP7_75t_R FILLER_355_601 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_607 ();
 DECAPx4_ASAP7_75t_R FILLER_355_622 ();
 FILLER_ASAP7_75t_R FILLER_355_632 ();
 DECAPx4_ASAP7_75t_R FILLER_355_640 ();
 FILLER_ASAP7_75t_R FILLER_355_650 ();
 DECAPx6_ASAP7_75t_R FILLER_355_666 ();
 DECAPx10_ASAP7_75t_R FILLER_355_691 ();
 DECAPx10_ASAP7_75t_R FILLER_355_713 ();
 DECAPx10_ASAP7_75t_R FILLER_355_735 ();
 DECAPx10_ASAP7_75t_R FILLER_355_757 ();
 DECAPx10_ASAP7_75t_R FILLER_355_779 ();
 DECAPx10_ASAP7_75t_R FILLER_355_801 ();
 DECAPx10_ASAP7_75t_R FILLER_355_823 ();
 DECAPx10_ASAP7_75t_R FILLER_355_845 ();
 DECAPx10_ASAP7_75t_R FILLER_355_867 ();
 DECAPx10_ASAP7_75t_R FILLER_355_889 ();
 DECAPx6_ASAP7_75t_R FILLER_355_911 ();
 DECAPx2_ASAP7_75t_R FILLER_355_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_355_933 ();
 DECAPx10_ASAP7_75t_R FILLER_356_2 ();
 DECAPx10_ASAP7_75t_R FILLER_356_24 ();
 DECAPx10_ASAP7_75t_R FILLER_356_46 ();
 DECAPx10_ASAP7_75t_R FILLER_356_68 ();
 DECAPx10_ASAP7_75t_R FILLER_356_90 ();
 FILLER_ASAP7_75t_R FILLER_356_112 ();
 DECAPx2_ASAP7_75t_R FILLER_356_120 ();
 DECAPx10_ASAP7_75t_R FILLER_356_134 ();
 DECAPx10_ASAP7_75t_R FILLER_356_156 ();
 DECAPx1_ASAP7_75t_R FILLER_356_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_182 ();
 DECAPx10_ASAP7_75t_R FILLER_356_192 ();
 FILLER_ASAP7_75t_R FILLER_356_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_222 ();
 DECAPx2_ASAP7_75t_R FILLER_356_229 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_235 ();
 DECAPx1_ASAP7_75t_R FILLER_356_242 ();
 DECAPx4_ASAP7_75t_R FILLER_356_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_259 ();
 DECAPx2_ASAP7_75t_R FILLER_356_272 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_278 ();
 DECAPx1_ASAP7_75t_R FILLER_356_285 ();
 DECAPx10_ASAP7_75t_R FILLER_356_292 ();
 DECAPx6_ASAP7_75t_R FILLER_356_314 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_356_328 ();
 DECAPx4_ASAP7_75t_R FILLER_356_339 ();
 FILLER_ASAP7_75t_R FILLER_356_349 ();
 DECAPx10_ASAP7_75t_R FILLER_356_357 ();
 DECAPx6_ASAP7_75t_R FILLER_356_379 ();
 DECAPx2_ASAP7_75t_R FILLER_356_393 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_447 ();
 DECAPx1_ASAP7_75t_R FILLER_356_458 ();
 FILLER_ASAP7_75t_R FILLER_356_470 ();
 DECAPx2_ASAP7_75t_R FILLER_356_482 ();
 DECAPx2_ASAP7_75t_R FILLER_356_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_506 ();
 DECAPx6_ASAP7_75t_R FILLER_356_513 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_356_527 ();
 DECAPx2_ASAP7_75t_R FILLER_356_544 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_356_550 ();
 DECAPx4_ASAP7_75t_R FILLER_356_556 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_566 ();
 DECAPx1_ASAP7_75t_R FILLER_356_570 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_574 ();
 DECAPx2_ASAP7_75t_R FILLER_356_581 ();
 DECAPx6_ASAP7_75t_R FILLER_356_590 ();
 DECAPx2_ASAP7_75t_R FILLER_356_604 ();
 DECAPx6_ASAP7_75t_R FILLER_356_627 ();
 DECAPx1_ASAP7_75t_R FILLER_356_641 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_645 ();
 DECAPx10_ASAP7_75t_R FILLER_356_663 ();
 DECAPx10_ASAP7_75t_R FILLER_356_685 ();
 DECAPx10_ASAP7_75t_R FILLER_356_707 ();
 DECAPx10_ASAP7_75t_R FILLER_356_729 ();
 DECAPx10_ASAP7_75t_R FILLER_356_751 ();
 DECAPx10_ASAP7_75t_R FILLER_356_773 ();
 DECAPx10_ASAP7_75t_R FILLER_356_795 ();
 DECAPx10_ASAP7_75t_R FILLER_356_817 ();
 DECAPx10_ASAP7_75t_R FILLER_356_839 ();
 DECAPx10_ASAP7_75t_R FILLER_356_861 ();
 DECAPx10_ASAP7_75t_R FILLER_356_883 ();
 DECAPx10_ASAP7_75t_R FILLER_356_905 ();
 DECAPx2_ASAP7_75t_R FILLER_356_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_356_933 ();
 DECAPx10_ASAP7_75t_R FILLER_357_2 ();
 DECAPx10_ASAP7_75t_R FILLER_357_24 ();
 DECAPx10_ASAP7_75t_R FILLER_357_46 ();
 DECAPx10_ASAP7_75t_R FILLER_357_68 ();
 DECAPx10_ASAP7_75t_R FILLER_357_90 ();
 DECAPx4_ASAP7_75t_R FILLER_357_112 ();
 FILLER_ASAP7_75t_R FILLER_357_122 ();
 DECAPx4_ASAP7_75t_R FILLER_357_138 ();
 FILLER_ASAP7_75t_R FILLER_357_148 ();
 DECAPx2_ASAP7_75t_R FILLER_357_156 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_162 ();
 DECAPx10_ASAP7_75t_R FILLER_357_179 ();
 DECAPx1_ASAP7_75t_R FILLER_357_201 ();
 DECAPx1_ASAP7_75t_R FILLER_357_219 ();
 DECAPx2_ASAP7_75t_R FILLER_357_229 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_235 ();
 DECAPx1_ASAP7_75t_R FILLER_357_244 ();
 DECAPx1_ASAP7_75t_R FILLER_357_256 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_260 ();
 DECAPx6_ASAP7_75t_R FILLER_357_267 ();
 DECAPx2_ASAP7_75t_R FILLER_357_281 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_287 ();
 DECAPx2_ASAP7_75t_R FILLER_357_294 ();
 FILLER_ASAP7_75t_R FILLER_357_300 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_310 ();
 DECAPx2_ASAP7_75t_R FILLER_357_317 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_323 ();
 DECAPx4_ASAP7_75t_R FILLER_357_340 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_350 ();
 DECAPx4_ASAP7_75t_R FILLER_357_365 ();
 FILLER_ASAP7_75t_R FILLER_357_398 ();
 FILLER_ASAP7_75t_R FILLER_357_426 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_447 ();
 DECAPx1_ASAP7_75t_R FILLER_357_458 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_462 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_471 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_485 ();
 DECAPx2_ASAP7_75t_R FILLER_357_496 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_502 ();
 DECAPx4_ASAP7_75t_R FILLER_357_522 ();
 DECAPx10_ASAP7_75t_R FILLER_357_538 ();
 DECAPx1_ASAP7_75t_R FILLER_357_560 ();
 FILLER_ASAP7_75t_R FILLER_357_567 ();
 DECAPx10_ASAP7_75t_R FILLER_357_583 ();
 DECAPx2_ASAP7_75t_R FILLER_357_605 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_611 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_357_617 ();
 DECAPx10_ASAP7_75t_R FILLER_357_632 ();
 DECAPx2_ASAP7_75t_R FILLER_357_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_660 ();
 DECAPx10_ASAP7_75t_R FILLER_357_681 ();
 DECAPx10_ASAP7_75t_R FILLER_357_703 ();
 DECAPx10_ASAP7_75t_R FILLER_357_725 ();
 DECAPx10_ASAP7_75t_R FILLER_357_747 ();
 DECAPx10_ASAP7_75t_R FILLER_357_769 ();
 DECAPx10_ASAP7_75t_R FILLER_357_791 ();
 DECAPx10_ASAP7_75t_R FILLER_357_813 ();
 DECAPx10_ASAP7_75t_R FILLER_357_835 ();
 DECAPx10_ASAP7_75t_R FILLER_357_857 ();
 DECAPx10_ASAP7_75t_R FILLER_357_879 ();
 DECAPx10_ASAP7_75t_R FILLER_357_901 ();
 FILLER_ASAP7_75t_R FILLER_357_923 ();
 DECAPx2_ASAP7_75t_R FILLER_357_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_357_933 ();
 DECAPx10_ASAP7_75t_R FILLER_358_2 ();
 DECAPx10_ASAP7_75t_R FILLER_358_24 ();
 DECAPx10_ASAP7_75t_R FILLER_358_46 ();
 DECAPx10_ASAP7_75t_R FILLER_358_68 ();
 DECAPx4_ASAP7_75t_R FILLER_358_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_358_100 ();
 DECAPx1_ASAP7_75t_R FILLER_358_109 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_113 ();
 DECAPx2_ASAP7_75t_R FILLER_358_117 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_123 ();
 DECAPx2_ASAP7_75t_R FILLER_358_130 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_358_136 ();
 DECAPx6_ASAP7_75t_R FILLER_358_168 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_358_182 ();
 DECAPx2_ASAP7_75t_R FILLER_358_191 ();
 FILLER_ASAP7_75t_R FILLER_358_197 ();
 DECAPx6_ASAP7_75t_R FILLER_358_263 ();
 FILLER_ASAP7_75t_R FILLER_358_317 ();
 DECAPx1_ASAP7_75t_R FILLER_358_325 ();
 DECAPx1_ASAP7_75t_R FILLER_358_335 ();
 DECAPx2_ASAP7_75t_R FILLER_358_346 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_352 ();
 DECAPx1_ASAP7_75t_R FILLER_358_361 ();
 FILLER_ASAP7_75t_R FILLER_358_377 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_439 ();
 FILLER_ASAP7_75t_R FILLER_358_455 ();
 DECAPx10_ASAP7_75t_R FILLER_358_464 ();
 DECAPx6_ASAP7_75t_R FILLER_358_486 ();
 DECAPx2_ASAP7_75t_R FILLER_358_500 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_506 ();
 DECAPx1_ASAP7_75t_R FILLER_358_519 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_523 ();
 DECAPx10_ASAP7_75t_R FILLER_358_535 ();
 DECAPx2_ASAP7_75t_R FILLER_358_557 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_358_563 ();
 FILLER_ASAP7_75t_R FILLER_358_580 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_596 ();
 DECAPx1_ASAP7_75t_R FILLER_358_600 ();
 DECAPx4_ASAP7_75t_R FILLER_358_610 ();
 FILLERxp5_ASAP7_75t_R FILLER_358_620 ();
 FILLER_ASAP7_75t_R FILLER_358_647 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_358_652 ();
 DECAPx2_ASAP7_75t_R FILLER_358_658 ();
 FILLER_ASAP7_75t_R FILLER_358_664 ();
 DECAPx10_ASAP7_75t_R FILLER_358_684 ();
 DECAPx10_ASAP7_75t_R FILLER_358_706 ();
 DECAPx10_ASAP7_75t_R FILLER_358_728 ();
 DECAPx10_ASAP7_75t_R FILLER_358_750 ();
 DECAPx10_ASAP7_75t_R FILLER_358_772 ();
 DECAPx10_ASAP7_75t_R FILLER_358_794 ();
 DECAPx10_ASAP7_75t_R FILLER_358_816 ();
 DECAPx10_ASAP7_75t_R FILLER_358_838 ();
 DECAPx10_ASAP7_75t_R FILLER_358_860 ();
 DECAPx10_ASAP7_75t_R FILLER_358_882 ();
 DECAPx10_ASAP7_75t_R FILLER_358_904 ();
 DECAPx2_ASAP7_75t_R FILLER_358_926 ();
 FILLER_ASAP7_75t_R FILLER_358_932 ();
 DECAPx10_ASAP7_75t_R FILLER_359_2 ();
 DECAPx10_ASAP7_75t_R FILLER_359_24 ();
 DECAPx10_ASAP7_75t_R FILLER_359_46 ();
 DECAPx10_ASAP7_75t_R FILLER_359_68 ();
 DECAPx6_ASAP7_75t_R FILLER_359_116 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_130 ();
 FILLER_ASAP7_75t_R FILLER_359_157 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_173 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_359_216 ();
 DECAPx2_ASAP7_75t_R FILLER_359_225 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_359_231 ();
 DECAPx1_ASAP7_75t_R FILLER_359_240 ();
 FILLER_ASAP7_75t_R FILLER_359_247 ();
 DECAPx2_ASAP7_75t_R FILLER_359_261 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_359_267 ();
 DECAPx1_ASAP7_75t_R FILLER_359_278 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_282 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_289 ();
 DECAPx1_ASAP7_75t_R FILLER_359_339 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_343 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_359_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_467 ();
 DECAPx2_ASAP7_75t_R FILLER_359_477 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_359_483 ();
 DECAPx6_ASAP7_75t_R FILLER_359_492 ();
 DECAPx1_ASAP7_75t_R FILLER_359_506 ();
 DECAPx2_ASAP7_75t_R FILLER_359_515 ();
 FILLER_ASAP7_75t_R FILLER_359_521 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_540 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_544 ();
 DECAPx4_ASAP7_75t_R FILLER_359_562 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_572 ();
 DECAPx1_ASAP7_75t_R FILLER_359_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_586 ();
 FILLER_ASAP7_75t_R FILLER_359_598 ();
 DECAPx6_ASAP7_75t_R FILLER_359_619 ();
 DECAPx2_ASAP7_75t_R FILLER_359_633 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_639 ();
 DECAPx10_ASAP7_75t_R FILLER_359_654 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_676 ();
 DECAPx10_ASAP7_75t_R FILLER_359_682 ();
 DECAPx10_ASAP7_75t_R FILLER_359_704 ();
 DECAPx10_ASAP7_75t_R FILLER_359_726 ();
 DECAPx10_ASAP7_75t_R FILLER_359_748 ();
 DECAPx10_ASAP7_75t_R FILLER_359_770 ();
 DECAPx10_ASAP7_75t_R FILLER_359_792 ();
 DECAPx10_ASAP7_75t_R FILLER_359_814 ();
 DECAPx10_ASAP7_75t_R FILLER_359_836 ();
 DECAPx10_ASAP7_75t_R FILLER_359_858 ();
 DECAPx10_ASAP7_75t_R FILLER_359_880 ();
 DECAPx10_ASAP7_75t_R FILLER_359_902 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_924 ();
 DECAPx2_ASAP7_75t_R FILLER_359_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_359_933 ();
 DECAPx10_ASAP7_75t_R FILLER_360_2 ();
 DECAPx10_ASAP7_75t_R FILLER_360_24 ();
 DECAPx10_ASAP7_75t_R FILLER_360_46 ();
 DECAPx10_ASAP7_75t_R FILLER_360_68 ();
 DECAPx2_ASAP7_75t_R FILLER_360_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_360_96 ();
 DECAPx2_ASAP7_75t_R FILLER_360_108 ();
 DECAPx6_ASAP7_75t_R FILLER_360_120 ();
 DECAPx2_ASAP7_75t_R FILLER_360_134 ();
 DECAPx1_ASAP7_75t_R FILLER_360_155 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_159 ();
 DECAPx6_ASAP7_75t_R FILLER_360_166 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_360_186 ();
 DECAPx10_ASAP7_75t_R FILLER_360_207 ();
 DECAPx10_ASAP7_75t_R FILLER_360_229 ();
 DECAPx6_ASAP7_75t_R FILLER_360_251 ();
 DECAPx10_ASAP7_75t_R FILLER_360_278 ();
 DECAPx10_ASAP7_75t_R FILLER_360_300 ();
 FILLER_ASAP7_75t_R FILLER_360_322 ();
 DECAPx2_ASAP7_75t_R FILLER_360_333 ();
 FILLER_ASAP7_75t_R FILLER_360_339 ();
 DECAPx1_ASAP7_75t_R FILLER_360_353 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_357 ();
 FILLER_ASAP7_75t_R FILLER_360_380 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_439 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_446 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_452 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_464 ();
 DECAPx1_ASAP7_75t_R FILLER_360_487 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_491 ();
 DECAPx6_ASAP7_75t_R FILLER_360_500 ();
 DECAPx2_ASAP7_75t_R FILLER_360_517 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_360_523 ();
 DECAPx2_ASAP7_75t_R FILLER_360_532 ();
 DECAPx6_ASAP7_75t_R FILLER_360_561 ();
 DECAPx2_ASAP7_75t_R FILLER_360_575 ();
 DECAPx10_ASAP7_75t_R FILLER_360_601 ();
 DECAPx6_ASAP7_75t_R FILLER_360_623 ();
 DECAPx2_ASAP7_75t_R FILLER_360_637 ();
 DECAPx10_ASAP7_75t_R FILLER_360_646 ();
 DECAPx10_ASAP7_75t_R FILLER_360_668 ();
 DECAPx10_ASAP7_75t_R FILLER_360_690 ();
 DECAPx10_ASAP7_75t_R FILLER_360_712 ();
 DECAPx10_ASAP7_75t_R FILLER_360_734 ();
 DECAPx10_ASAP7_75t_R FILLER_360_756 ();
 DECAPx10_ASAP7_75t_R FILLER_360_778 ();
 DECAPx6_ASAP7_75t_R FILLER_360_800 ();
 DECAPx1_ASAP7_75t_R FILLER_360_814 ();
 DECAPx10_ASAP7_75t_R FILLER_360_823 ();
 DECAPx10_ASAP7_75t_R FILLER_360_845 ();
 DECAPx10_ASAP7_75t_R FILLER_360_867 ();
 DECAPx10_ASAP7_75t_R FILLER_360_889 ();
 DECAPx10_ASAP7_75t_R FILLER_360_911 ();
 FILLERxp5_ASAP7_75t_R FILLER_360_933 ();
 DECAPx10_ASAP7_75t_R FILLER_361_2 ();
 DECAPx10_ASAP7_75t_R FILLER_361_24 ();
 DECAPx10_ASAP7_75t_R FILLER_361_46 ();
 DECAPx10_ASAP7_75t_R FILLER_361_68 ();
 DECAPx4_ASAP7_75t_R FILLER_361_90 ();
 FILLER_ASAP7_75t_R FILLER_361_100 ();
 DECAPx10_ASAP7_75t_R FILLER_361_131 ();
 DECAPx10_ASAP7_75t_R FILLER_361_153 ();
 DECAPx1_ASAP7_75t_R FILLER_361_175 ();
 DECAPx10_ASAP7_75t_R FILLER_361_191 ();
 DECAPx10_ASAP7_75t_R FILLER_361_213 ();
 FILLER_ASAP7_75t_R FILLER_361_235 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_361_243 ();
 DECAPx4_ASAP7_75t_R FILLER_361_249 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_259 ();
 FILLER_ASAP7_75t_R FILLER_361_266 ();
 DECAPx10_ASAP7_75t_R FILLER_361_277 ();
 DECAPx10_ASAP7_75t_R FILLER_361_299 ();
 DECAPx10_ASAP7_75t_R FILLER_361_321 ();
 DECAPx1_ASAP7_75t_R FILLER_361_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_389 ();
 FILLER_ASAP7_75t_R FILLER_361_442 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_481 ();
 FILLER_ASAP7_75t_R FILLER_361_507 ();
 DECAPx6_ASAP7_75t_R FILLER_361_524 ();
 DECAPx2_ASAP7_75t_R FILLER_361_538 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_544 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_557 ();
 DECAPx2_ASAP7_75t_R FILLER_361_561 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_567 ();
 DECAPx10_ASAP7_75t_R FILLER_361_571 ();
 DECAPx2_ASAP7_75t_R FILLER_361_593 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_599 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_361_603 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_609 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_361_613 ();
 DECAPx1_ASAP7_75t_R FILLER_361_619 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_626 ();
 DECAPx10_ASAP7_75t_R FILLER_361_647 ();
 DECAPx10_ASAP7_75t_R FILLER_361_669 ();
 DECAPx10_ASAP7_75t_R FILLER_361_691 ();
 DECAPx10_ASAP7_75t_R FILLER_361_713 ();
 DECAPx10_ASAP7_75t_R FILLER_361_735 ();
 DECAPx10_ASAP7_75t_R FILLER_361_757 ();
 DECAPx10_ASAP7_75t_R FILLER_361_779 ();
 DECAPx10_ASAP7_75t_R FILLER_361_801 ();
 DECAPx10_ASAP7_75t_R FILLER_361_823 ();
 DECAPx10_ASAP7_75t_R FILLER_361_845 ();
 DECAPx10_ASAP7_75t_R FILLER_361_867 ();
 DECAPx10_ASAP7_75t_R FILLER_361_889 ();
 DECAPx6_ASAP7_75t_R FILLER_361_911 ();
 DECAPx2_ASAP7_75t_R FILLER_361_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_361_933 ();
 DECAPx10_ASAP7_75t_R FILLER_362_2 ();
 DECAPx10_ASAP7_75t_R FILLER_362_24 ();
 DECAPx10_ASAP7_75t_R FILLER_362_46 ();
 DECAPx10_ASAP7_75t_R FILLER_362_68 ();
 DECAPx6_ASAP7_75t_R FILLER_362_90 ();
 DECAPx1_ASAP7_75t_R FILLER_362_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_108 ();
 FILLER_ASAP7_75t_R FILLER_362_115 ();
 DECAPx6_ASAP7_75t_R FILLER_362_120 ();
 DECAPx2_ASAP7_75t_R FILLER_362_134 ();
 FILLER_ASAP7_75t_R FILLER_362_146 ();
 DECAPx6_ASAP7_75t_R FILLER_362_151 ();
 DECAPx2_ASAP7_75t_R FILLER_362_165 ();
 DECAPx6_ASAP7_75t_R FILLER_362_197 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_211 ();
 DECAPx2_ASAP7_75t_R FILLER_362_218 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_224 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_362_251 ();
 FILLER_ASAP7_75t_R FILLER_362_280 ();
 DECAPx2_ASAP7_75t_R FILLER_362_297 ();
 DECAPx1_ASAP7_75t_R FILLER_362_312 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_322 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_329 ();
 FILLER_ASAP7_75t_R FILLER_362_333 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_355 ();
 FILLER_ASAP7_75t_R FILLER_362_396 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_435 ();
 FILLER_ASAP7_75t_R FILLER_362_450 ();
 FILLERxp5_ASAP7_75t_R FILLER_362_476 ();
 FILLER_ASAP7_75t_R FILLER_362_487 ();
 FILLER_ASAP7_75t_R FILLER_362_505 ();
 DECAPx10_ASAP7_75t_R FILLER_362_521 ();
 DECAPx6_ASAP7_75t_R FILLER_362_543 ();
 FILLER_ASAP7_75t_R FILLER_362_557 ();
 DECAPx10_ASAP7_75t_R FILLER_362_579 ();
 DECAPx2_ASAP7_75t_R FILLER_362_643 ();
 FILLER_ASAP7_75t_R FILLER_362_672 ();
 DECAPx10_ASAP7_75t_R FILLER_362_683 ();
 DECAPx10_ASAP7_75t_R FILLER_362_705 ();
 DECAPx10_ASAP7_75t_R FILLER_362_727 ();
 DECAPx10_ASAP7_75t_R FILLER_362_749 ();
 DECAPx10_ASAP7_75t_R FILLER_362_771 ();
 DECAPx10_ASAP7_75t_R FILLER_362_793 ();
 DECAPx10_ASAP7_75t_R FILLER_362_815 ();
 DECAPx10_ASAP7_75t_R FILLER_362_837 ();
 DECAPx10_ASAP7_75t_R FILLER_362_859 ();
 DECAPx10_ASAP7_75t_R FILLER_362_881 ();
 DECAPx10_ASAP7_75t_R FILLER_362_903 ();
 DECAPx2_ASAP7_75t_R FILLER_362_925 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_362_931 ();
 DECAPx10_ASAP7_75t_R FILLER_363_2 ();
 DECAPx10_ASAP7_75t_R FILLER_363_24 ();
 DECAPx10_ASAP7_75t_R FILLER_363_46 ();
 DECAPx10_ASAP7_75t_R FILLER_363_68 ();
 DECAPx10_ASAP7_75t_R FILLER_363_90 ();
 DECAPx2_ASAP7_75t_R FILLER_363_112 ();
 FILLER_ASAP7_75t_R FILLER_363_118 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_126 ();
 DECAPx6_ASAP7_75t_R FILLER_363_165 ();
 DECAPx2_ASAP7_75t_R FILLER_363_179 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_185 ();
 DECAPx6_ASAP7_75t_R FILLER_363_189 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_203 ();
 FILLER_ASAP7_75t_R FILLER_363_230 ();
 FILLER_ASAP7_75t_R FILLER_363_238 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_243 ();
 DECAPx1_ASAP7_75t_R FILLER_363_275 ();
 FILLER_ASAP7_75t_R FILLER_363_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_336 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_438 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_472 ();
 DECAPx6_ASAP7_75t_R FILLER_363_518 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_532 ();
 DECAPx1_ASAP7_75t_R FILLER_363_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_540 ();
 DECAPx6_ASAP7_75t_R FILLER_363_544 ();
 DECAPx2_ASAP7_75t_R FILLER_363_558 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_567 ();
 DECAPx10_ASAP7_75t_R FILLER_363_582 ();
 DECAPx2_ASAP7_75t_R FILLER_363_604 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_610 ();
 DECAPx2_ASAP7_75t_R FILLER_363_614 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_363_620 ();
 DECAPx4_ASAP7_75t_R FILLER_363_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_640 ();
 DECAPx1_ASAP7_75t_R FILLER_363_644 ();
 FILLER_ASAP7_75t_R FILLER_363_651 ();
 FILLER_ASAP7_75t_R FILLER_363_667 ();
 DECAPx10_ASAP7_75t_R FILLER_363_689 ();
 DECAPx10_ASAP7_75t_R FILLER_363_711 ();
 DECAPx10_ASAP7_75t_R FILLER_363_733 ();
 DECAPx10_ASAP7_75t_R FILLER_363_755 ();
 DECAPx10_ASAP7_75t_R FILLER_363_777 ();
 DECAPx10_ASAP7_75t_R FILLER_363_799 ();
 DECAPx10_ASAP7_75t_R FILLER_363_821 ();
 DECAPx10_ASAP7_75t_R FILLER_363_843 ();
 DECAPx10_ASAP7_75t_R FILLER_363_865 ();
 DECAPx10_ASAP7_75t_R FILLER_363_887 ();
 DECAPx6_ASAP7_75t_R FILLER_363_909 ();
 FILLER_ASAP7_75t_R FILLER_363_923 ();
 DECAPx2_ASAP7_75t_R FILLER_363_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_363_933 ();
 DECAPx10_ASAP7_75t_R FILLER_364_2 ();
 DECAPx10_ASAP7_75t_R FILLER_364_24 ();
 DECAPx10_ASAP7_75t_R FILLER_364_46 ();
 DECAPx10_ASAP7_75t_R FILLER_364_68 ();
 DECAPx6_ASAP7_75t_R FILLER_364_90 ();
 DECAPx1_ASAP7_75t_R FILLER_364_104 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_108 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_135 ();
 FILLER_ASAP7_75t_R FILLER_364_145 ();
 DECAPx10_ASAP7_75t_R FILLER_364_173 ();
 DECAPx2_ASAP7_75t_R FILLER_364_195 ();
 FILLER_ASAP7_75t_R FILLER_364_201 ();
 FILLER_ASAP7_75t_R FILLER_364_206 ();
 DECAPx1_ASAP7_75t_R FILLER_364_214 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_218 ();
 DECAPx1_ASAP7_75t_R FILLER_364_231 ();
 DECAPx2_ASAP7_75t_R FILLER_364_250 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_256 ();
 DECAPx10_ASAP7_75t_R FILLER_364_260 ();
 DECAPx4_ASAP7_75t_R FILLER_364_282 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_364_292 ();
 FILLER_ASAP7_75t_R FILLER_364_327 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_335 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_342 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_352 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_428 ();
 FILLER_ASAP7_75t_R FILLER_364_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_524 ();
 DECAPx6_ASAP7_75t_R FILLER_364_559 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_364_573 ();
 DECAPx1_ASAP7_75t_R FILLER_364_583 ();
 FILLERxp5_ASAP7_75t_R FILLER_364_587 ();
 DECAPx10_ASAP7_75t_R FILLER_364_600 ();
 DECAPx10_ASAP7_75t_R FILLER_364_622 ();
 DECAPx2_ASAP7_75t_R FILLER_364_644 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_364_650 ();
 FILLER_ASAP7_75t_R FILLER_364_668 ();
 DECAPx10_ASAP7_75t_R FILLER_364_679 ();
 DECAPx10_ASAP7_75t_R FILLER_364_701 ();
 DECAPx10_ASAP7_75t_R FILLER_364_723 ();
 DECAPx10_ASAP7_75t_R FILLER_364_745 ();
 DECAPx10_ASAP7_75t_R FILLER_364_767 ();
 DECAPx10_ASAP7_75t_R FILLER_364_789 ();
 DECAPx10_ASAP7_75t_R FILLER_364_811 ();
 DECAPx10_ASAP7_75t_R FILLER_364_833 ();
 DECAPx10_ASAP7_75t_R FILLER_364_855 ();
 DECAPx10_ASAP7_75t_R FILLER_364_877 ();
 DECAPx10_ASAP7_75t_R FILLER_364_899 ();
 DECAPx4_ASAP7_75t_R FILLER_364_921 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_364_931 ();
 DECAPx10_ASAP7_75t_R FILLER_365_2 ();
 DECAPx10_ASAP7_75t_R FILLER_365_24 ();
 DECAPx10_ASAP7_75t_R FILLER_365_46 ();
 DECAPx10_ASAP7_75t_R FILLER_365_68 ();
 DECAPx10_ASAP7_75t_R FILLER_365_90 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_365_112 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_365_121 ();
 DECAPx10_ASAP7_75t_R FILLER_365_127 ();
 DECAPx4_ASAP7_75t_R FILLER_365_149 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_365_159 ();
 DECAPx4_ASAP7_75t_R FILLER_365_165 ();
 FILLER_ASAP7_75t_R FILLER_365_175 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_365_203 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_365_258 ();
 DECAPx2_ASAP7_75t_R FILLER_365_287 ();
 FILLER_ASAP7_75t_R FILLER_365_293 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_317 ();
 FILLER_ASAP7_75t_R FILLER_365_349 ();
 FILLER_ASAP7_75t_R FILLER_365_362 ();
 FILLER_ASAP7_75t_R FILLER_365_385 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_393 ();
 FILLER_ASAP7_75t_R FILLER_365_428 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_476 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_518 ();
 DECAPx2_ASAP7_75t_R FILLER_365_536 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_542 ();
 DECAPx2_ASAP7_75t_R FILLER_365_546 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_556 ();
 DECAPx2_ASAP7_75t_R FILLER_365_571 ();
 FILLER_ASAP7_75t_R FILLER_365_577 ();
 DECAPx10_ASAP7_75t_R FILLER_365_599 ();
 DECAPx10_ASAP7_75t_R FILLER_365_621 ();
 DECAPx10_ASAP7_75t_R FILLER_365_643 ();
 FILLER_ASAP7_75t_R FILLER_365_665 ();
 DECAPx10_ASAP7_75t_R FILLER_365_673 ();
 DECAPx10_ASAP7_75t_R FILLER_365_695 ();
 DECAPx10_ASAP7_75t_R FILLER_365_717 ();
 DECAPx10_ASAP7_75t_R FILLER_365_739 ();
 DECAPx10_ASAP7_75t_R FILLER_365_761 ();
 DECAPx10_ASAP7_75t_R FILLER_365_783 ();
 DECAPx10_ASAP7_75t_R FILLER_365_805 ();
 DECAPx10_ASAP7_75t_R FILLER_365_827 ();
 DECAPx10_ASAP7_75t_R FILLER_365_849 ();
 DECAPx10_ASAP7_75t_R FILLER_365_871 ();
 DECAPx10_ASAP7_75t_R FILLER_365_893 ();
 DECAPx4_ASAP7_75t_R FILLER_365_915 ();
 DECAPx2_ASAP7_75t_R FILLER_365_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_365_933 ();
 DECAPx10_ASAP7_75t_R FILLER_366_2 ();
 DECAPx10_ASAP7_75t_R FILLER_366_24 ();
 DECAPx10_ASAP7_75t_R FILLER_366_46 ();
 DECAPx10_ASAP7_75t_R FILLER_366_68 ();
 DECAPx10_ASAP7_75t_R FILLER_366_90 ();
 DECAPx10_ASAP7_75t_R FILLER_366_112 ();
 DECAPx10_ASAP7_75t_R FILLER_366_134 ();
 DECAPx6_ASAP7_75t_R FILLER_366_156 ();
 DECAPx2_ASAP7_75t_R FILLER_366_170 ();
 FILLER_ASAP7_75t_R FILLER_366_220 ();
 DECAPx10_ASAP7_75t_R FILLER_366_225 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_247 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_254 ();
 FILLER_ASAP7_75t_R FILLER_366_261 ();
 DECAPx1_ASAP7_75t_R FILLER_366_275 ();
 FILLER_ASAP7_75t_R FILLER_366_305 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_373 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_400 ();
 FILLER_ASAP7_75t_R FILLER_366_460 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_464 ();
 DECAPx10_ASAP7_75t_R FILLER_366_541 ();
 DECAPx10_ASAP7_75t_R FILLER_366_563 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_366_585 ();
 DECAPx4_ASAP7_75t_R FILLER_366_602 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_366_612 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_627 ();
 DECAPx10_ASAP7_75t_R FILLER_366_643 ();
 DECAPx10_ASAP7_75t_R FILLER_366_665 ();
 DECAPx10_ASAP7_75t_R FILLER_366_687 ();
 DECAPx10_ASAP7_75t_R FILLER_366_709 ();
 DECAPx10_ASAP7_75t_R FILLER_366_731 ();
 DECAPx10_ASAP7_75t_R FILLER_366_753 ();
 DECAPx10_ASAP7_75t_R FILLER_366_775 ();
 DECAPx10_ASAP7_75t_R FILLER_366_797 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_819 ();
 DECAPx10_ASAP7_75t_R FILLER_366_825 ();
 DECAPx10_ASAP7_75t_R FILLER_366_847 ();
 DECAPx10_ASAP7_75t_R FILLER_366_869 ();
 DECAPx10_ASAP7_75t_R FILLER_366_891 ();
 DECAPx6_ASAP7_75t_R FILLER_366_913 ();
 DECAPx2_ASAP7_75t_R FILLER_366_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_366_933 ();
 DECAPx10_ASAP7_75t_R FILLER_367_2 ();
 DECAPx10_ASAP7_75t_R FILLER_367_24 ();
 DECAPx10_ASAP7_75t_R FILLER_367_46 ();
 DECAPx10_ASAP7_75t_R FILLER_367_68 ();
 DECAPx10_ASAP7_75t_R FILLER_367_90 ();
 DECAPx10_ASAP7_75t_R FILLER_367_112 ();
 DECAPx10_ASAP7_75t_R FILLER_367_134 ();
 DECAPx10_ASAP7_75t_R FILLER_367_156 ();
 DECAPx4_ASAP7_75t_R FILLER_367_178 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_188 ();
 FILLER_ASAP7_75t_R FILLER_367_198 ();
 DECAPx10_ASAP7_75t_R FILLER_367_209 ();
 DECAPx4_ASAP7_75t_R FILLER_367_231 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_367_241 ();
 DECAPx1_ASAP7_75t_R FILLER_367_270 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_274 ();
 FILLER_ASAP7_75t_R FILLER_367_290 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_469 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_493 ();
 FILLER_ASAP7_75t_R FILLER_367_504 ();
 FILLER_ASAP7_75t_R FILLER_367_517 ();
 DECAPx4_ASAP7_75t_R FILLER_367_552 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_565 ();
 DECAPx6_ASAP7_75t_R FILLER_367_575 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_367_589 ();
 FILLER_ASAP7_75t_R FILLER_367_595 ();
 DECAPx2_ASAP7_75t_R FILLER_367_600 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_606 ();
 DECAPx1_ASAP7_75t_R FILLER_367_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_636 ();
 DECAPx2_ASAP7_75t_R FILLER_367_654 ();
 DECAPx10_ASAP7_75t_R FILLER_367_663 ();
 DECAPx10_ASAP7_75t_R FILLER_367_685 ();
 DECAPx10_ASAP7_75t_R FILLER_367_707 ();
 DECAPx10_ASAP7_75t_R FILLER_367_729 ();
 DECAPx10_ASAP7_75t_R FILLER_367_751 ();
 DECAPx10_ASAP7_75t_R FILLER_367_773 ();
 DECAPx10_ASAP7_75t_R FILLER_367_795 ();
 DECAPx10_ASAP7_75t_R FILLER_367_817 ();
 DECAPx10_ASAP7_75t_R FILLER_367_839 ();
 DECAPx10_ASAP7_75t_R FILLER_367_861 ();
 DECAPx10_ASAP7_75t_R FILLER_367_883 ();
 DECAPx6_ASAP7_75t_R FILLER_367_905 ();
 DECAPx2_ASAP7_75t_R FILLER_367_919 ();
 DECAPx2_ASAP7_75t_R FILLER_367_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_367_933 ();
 DECAPx10_ASAP7_75t_R FILLER_368_2 ();
 DECAPx10_ASAP7_75t_R FILLER_368_24 ();
 DECAPx10_ASAP7_75t_R FILLER_368_46 ();
 DECAPx10_ASAP7_75t_R FILLER_368_68 ();
 DECAPx10_ASAP7_75t_R FILLER_368_90 ();
 DECAPx10_ASAP7_75t_R FILLER_368_112 ();
 DECAPx10_ASAP7_75t_R FILLER_368_134 ();
 DECAPx10_ASAP7_75t_R FILLER_368_156 ();
 DECAPx10_ASAP7_75t_R FILLER_368_178 ();
 DECAPx10_ASAP7_75t_R FILLER_368_200 ();
 DECAPx10_ASAP7_75t_R FILLER_368_222 ();
 DECAPx6_ASAP7_75t_R FILLER_368_244 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_258 ();
 DECAPx6_ASAP7_75t_R FILLER_368_262 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_368_276 ();
 FILLER_ASAP7_75t_R FILLER_368_298 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_306 ();
 FILLER_ASAP7_75t_R FILLER_368_328 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_336 ();
 FILLER_ASAP7_75t_R FILLER_368_432 ();
 FILLER_ASAP7_75t_R FILLER_368_451 ();
 FILLER_ASAP7_75t_R FILLER_368_460 ();
 FILLER_ASAP7_75t_R FILLER_368_464 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_497 ();
 FILLER_ASAP7_75t_R FILLER_368_532 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_592 ();
 FILLER_ASAP7_75t_R FILLER_368_598 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_626 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_644 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_660 ();
 DECAPx10_ASAP7_75t_R FILLER_368_673 ();
 DECAPx10_ASAP7_75t_R FILLER_368_695 ();
 DECAPx10_ASAP7_75t_R FILLER_368_717 ();
 DECAPx10_ASAP7_75t_R FILLER_368_739 ();
 DECAPx10_ASAP7_75t_R FILLER_368_761 ();
 DECAPx10_ASAP7_75t_R FILLER_368_783 ();
 DECAPx10_ASAP7_75t_R FILLER_368_805 ();
 DECAPx10_ASAP7_75t_R FILLER_368_827 ();
 DECAPx10_ASAP7_75t_R FILLER_368_849 ();
 DECAPx10_ASAP7_75t_R FILLER_368_871 ();
 DECAPx10_ASAP7_75t_R FILLER_368_893 ();
 DECAPx6_ASAP7_75t_R FILLER_368_915 ();
 DECAPx1_ASAP7_75t_R FILLER_368_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_368_933 ();
 DECAPx10_ASAP7_75t_R FILLER_369_2 ();
 DECAPx10_ASAP7_75t_R FILLER_369_24 ();
 DECAPx10_ASAP7_75t_R FILLER_369_46 ();
 DECAPx10_ASAP7_75t_R FILLER_369_68 ();
 DECAPx10_ASAP7_75t_R FILLER_369_90 ();
 DECAPx10_ASAP7_75t_R FILLER_369_112 ();
 DECAPx10_ASAP7_75t_R FILLER_369_134 ();
 DECAPx10_ASAP7_75t_R FILLER_369_156 ();
 DECAPx10_ASAP7_75t_R FILLER_369_178 ();
 DECAPx10_ASAP7_75t_R FILLER_369_200 ();
 DECAPx10_ASAP7_75t_R FILLER_369_222 ();
 DECAPx10_ASAP7_75t_R FILLER_369_244 ();
 DECAPx2_ASAP7_75t_R FILLER_369_266 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_369_272 ();
 FILLER_ASAP7_75t_R FILLER_369_343 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_467 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_484 ();
 FILLER_ASAP7_75t_R FILLER_369_531 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_550 ();
 FILLER_ASAP7_75t_R FILLER_369_576 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_615 ();
 DECAPx1_ASAP7_75t_R FILLER_369_636 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_640 ();
 FILLER_ASAP7_75t_R FILLER_369_655 ();
 DECAPx10_ASAP7_75t_R FILLER_369_677 ();
 DECAPx10_ASAP7_75t_R FILLER_369_699 ();
 DECAPx10_ASAP7_75t_R FILLER_369_721 ();
 DECAPx10_ASAP7_75t_R FILLER_369_743 ();
 DECAPx10_ASAP7_75t_R FILLER_369_765 ();
 DECAPx10_ASAP7_75t_R FILLER_369_787 ();
 DECAPx2_ASAP7_75t_R FILLER_369_814 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_820 ();
 DECAPx10_ASAP7_75t_R FILLER_369_826 ();
 DECAPx10_ASAP7_75t_R FILLER_369_848 ();
 DECAPx10_ASAP7_75t_R FILLER_369_870 ();
 DECAPx10_ASAP7_75t_R FILLER_369_892 ();
 DECAPx4_ASAP7_75t_R FILLER_369_914 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_924 ();
 DECAPx2_ASAP7_75t_R FILLER_369_927 ();
 FILLERxp5_ASAP7_75t_R FILLER_369_933 ();
 DECAPx10_ASAP7_75t_R FILLER_370_2 ();
 DECAPx10_ASAP7_75t_R FILLER_370_24 ();
 DECAPx10_ASAP7_75t_R FILLER_370_46 ();
 DECAPx10_ASAP7_75t_R FILLER_370_68 ();
 DECAPx10_ASAP7_75t_R FILLER_370_90 ();
 DECAPx10_ASAP7_75t_R FILLER_370_112 ();
 DECAPx10_ASAP7_75t_R FILLER_370_134 ();
 DECAPx10_ASAP7_75t_R FILLER_370_156 ();
 DECAPx10_ASAP7_75t_R FILLER_370_178 ();
 DECAPx10_ASAP7_75t_R FILLER_370_200 ();
 DECAPx10_ASAP7_75t_R FILLER_370_222 ();
 DECAPx10_ASAP7_75t_R FILLER_370_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_370_266 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_456 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_464 ();
 FILLER_ASAP7_75t_R FILLER_370_478 ();
 FILLER_ASAP7_75t_R FILLER_370_485 ();
 FILLER_ASAP7_75t_R FILLER_370_535 ();
 DECAPx2_ASAP7_75t_R FILLER_370_574 ();
 DECAPx6_ASAP7_75t_R FILLER_370_586 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_600 ();
 FILLER_ASAP7_75t_R FILLER_370_617 ();
 DECAPx10_ASAP7_75t_R FILLER_370_624 ();
 DECAPx10_ASAP7_75t_R FILLER_370_652 ();
 DECAPx10_ASAP7_75t_R FILLER_370_674 ();
 DECAPx10_ASAP7_75t_R FILLER_370_696 ();
 DECAPx10_ASAP7_75t_R FILLER_370_718 ();
 DECAPx10_ASAP7_75t_R FILLER_370_740 ();
 DECAPx10_ASAP7_75t_R FILLER_370_762 ();
 DECAPx6_ASAP7_75t_R FILLER_370_784 ();
 DECAPx2_ASAP7_75t_R FILLER_370_798 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_804 ();
 DECAPx2_ASAP7_75t_R FILLER_370_820 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_826 ();
 DECAPx10_ASAP7_75t_R FILLER_370_849 ();
 DECAPx10_ASAP7_75t_R FILLER_370_871 ();
 DECAPx10_ASAP7_75t_R FILLER_370_893 ();
 DECAPx6_ASAP7_75t_R FILLER_370_915 ();
 DECAPx1_ASAP7_75t_R FILLER_370_929 ();
 FILLERxp5_ASAP7_75t_R FILLER_370_933 ();
 DECAPx10_ASAP7_75t_R FILLER_371_2 ();
 DECAPx10_ASAP7_75t_R FILLER_371_24 ();
 DECAPx10_ASAP7_75t_R FILLER_371_46 ();
 DECAPx10_ASAP7_75t_R FILLER_371_68 ();
 DECAPx10_ASAP7_75t_R FILLER_371_90 ();
 DECAPx10_ASAP7_75t_R FILLER_371_112 ();
 DECAPx10_ASAP7_75t_R FILLER_371_134 ();
 DECAPx10_ASAP7_75t_R FILLER_371_156 ();
 DECAPx10_ASAP7_75t_R FILLER_371_178 ();
 DECAPx10_ASAP7_75t_R FILLER_371_200 ();
 DECAPx10_ASAP7_75t_R FILLER_371_222 ();
 DECAPx4_ASAP7_75t_R FILLER_371_244 ();
 TAPCELL_WITH_FILLER_ASAP7_75t_R FILLER_371_254 ();
 FILLER_ASAP7_75t_R FILLER_371_464 ();
 DECAPx10_ASAP7_75t_R FILLER_371_586 ();
 DECAPx10_ASAP7_75t_R FILLER_371_608 ();
 DECAPx10_ASAP7_75t_R FILLER_371_630 ();
 DECAPx10_ASAP7_75t_R FILLER_371_652 ();
 DECAPx10_ASAP7_75t_R FILLER_371_674 ();
 DECAPx10_ASAP7_75t_R FILLER_371_696 ();
 DECAPx10_ASAP7_75t_R FILLER_371_718 ();
 DECAPx10_ASAP7_75t_R FILLER_371_740 ();
 DECAPx10_ASAP7_75t_R FILLER_371_762 ();
 DECAPx4_ASAP7_75t_R FILLER_371_784 ();
 FILLERxp5_ASAP7_75t_R FILLER_371_794 ();
 DECAPx10_ASAP7_75t_R FILLER_371_832 ();
 DECAPx10_ASAP7_75t_R FILLER_371_854 ();
 DECAPx10_ASAP7_75t_R FILLER_371_876 ();
 DECAPx10_ASAP7_75t_R FILLER_371_898 ();
 DECAPx1_ASAP7_75t_R FILLER_371_920 ();
 DECAPx2_ASAP7_75t_R FILLER_371_926 ();
 FILLER_ASAP7_75t_R FILLER_371_932 ();
 assign alert_major_o = net461;
endmodule
